* NGSPICE file created from user_project_wrapper.ext - technology: sky130B

* Black-box entry subcircuit for core abstract view
.subckt core dbg_in[0] dbg_in[1] dbg_in[2] dbg_in[3] dbg_out[0] dbg_out[10] dbg_out[11]
+ dbg_out[12] dbg_out[13] dbg_out[14] dbg_out[15] dbg_out[16] dbg_out[17] dbg_out[18]
+ dbg_out[19] dbg_out[1] dbg_out[20] dbg_out[21] dbg_out[22] dbg_out[23] dbg_out[24]
+ dbg_out[25] dbg_out[26] dbg_out[27] dbg_out[28] dbg_out[29] dbg_out[2] dbg_out[30]
+ dbg_out[31] dbg_out[32] dbg_out[33] dbg_out[34] dbg_out[35] dbg_out[3] dbg_out[4]
+ dbg_out[5] dbg_out[6] dbg_out[7] dbg_out[8] dbg_out[9] dbg_pc[0] dbg_pc[10] dbg_pc[11]
+ dbg_pc[12] dbg_pc[13] dbg_pc[14] dbg_pc[15] dbg_pc[1] dbg_pc[2] dbg_pc[3] dbg_pc[4]
+ dbg_pc[5] dbg_pc[6] dbg_pc[7] dbg_pc[8] dbg_pc[9] dbg_r0[0] dbg_r0[10] dbg_r0[11]
+ dbg_r0[12] dbg_r0[13] dbg_r0[14] dbg_r0[15] dbg_r0[1] dbg_r0[2] dbg_r0[3] dbg_r0[4]
+ dbg_r0[5] dbg_r0[6] dbg_r0[7] dbg_r0[8] dbg_r0[9] i_clk i_irq i_mem_ack i_mem_data[0]
+ i_mem_data[10] i_mem_data[11] i_mem_data[12] i_mem_data[13] i_mem_data[14] i_mem_data[15]
+ i_mem_data[1] i_mem_data[2] i_mem_data[3] i_mem_data[4] i_mem_data[5] i_mem_data[6]
+ i_mem_data[7] i_mem_data[8] i_mem_data[9] i_mem_exception i_req_data[0] i_req_data[10]
+ i_req_data[11] i_req_data[12] i_req_data[13] i_req_data[14] i_req_data[15] i_req_data[16]
+ i_req_data[17] i_req_data[18] i_req_data[19] i_req_data[1] i_req_data[20] i_req_data[21]
+ i_req_data[22] i_req_data[23] i_req_data[24] i_req_data[25] i_req_data[26] i_req_data[27]
+ i_req_data[28] i_req_data[29] i_req_data[2] i_req_data[30] i_req_data[31] i_req_data[3]
+ i_req_data[4] i_req_data[5] i_req_data[6] i_req_data[7] i_req_data[8] i_req_data[9]
+ i_req_data_valid i_rst o_c_data_page o_c_instr_page o_icache_flush o_mem_addr[0]
+ o_mem_addr[10] o_mem_addr[11] o_mem_addr[12] o_mem_addr[13] o_mem_addr[14] o_mem_addr[15]
+ o_mem_addr[1] o_mem_addr[2] o_mem_addr[3] o_mem_addr[4] o_mem_addr[5] o_mem_addr[6]
+ o_mem_addr[7] o_mem_addr[8] o_mem_addr[9] o_mem_data[0] o_mem_data[10] o_mem_data[11]
+ o_mem_data[12] o_mem_data[13] o_mem_data[14] o_mem_data[15] o_mem_data[1] o_mem_data[2]
+ o_mem_data[3] o_mem_data[4] o_mem_data[5] o_mem_data[6] o_mem_data[7] o_mem_data[8]
+ o_mem_data[9] o_mem_req o_mem_sel[0] o_mem_sel[1] o_mem_we o_req_active o_req_addr[0]
+ o_req_addr[10] o_req_addr[11] o_req_addr[12] o_req_addr[13] o_req_addr[14] o_req_addr[15]
+ o_req_addr[1] o_req_addr[2] o_req_addr[3] o_req_addr[4] o_req_addr[5] o_req_addr[6]
+ o_req_addr[7] o_req_addr[8] o_req_addr[9] o_req_ppl_submit sr_bus_addr[0] sr_bus_addr[10]
+ sr_bus_addr[11] sr_bus_addr[12] sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15]
+ sr_bus_addr[1] sr_bus_addr[2] sr_bus_addr[3] sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6]
+ sr_bus_addr[7] sr_bus_addr[8] sr_bus_addr[9] sr_bus_data_o[0] sr_bus_data_o[10]
+ sr_bus_data_o[11] sr_bus_data_o[12] sr_bus_data_o[13] sr_bus_data_o[14] sr_bus_data_o[15]
+ sr_bus_data_o[1] sr_bus_data_o[2] sr_bus_data_o[3] sr_bus_data_o[4] sr_bus_data_o[5]
+ sr_bus_data_o[6] sr_bus_data_o[7] sr_bus_data_o[8] sr_bus_data_o[9] sr_bus_we vccd1
+ vssd1
.ends

* Black-box entry subcircuit for wb_cross_clk abstract view
.subckt wb_cross_clk clk_m clk_s m_rst m_wb_4_burst m_wb_8_burst m_wb_ack m_wb_adr[0]
+ m_wb_adr[10] m_wb_adr[11] m_wb_adr[12] m_wb_adr[13] m_wb_adr[14] m_wb_adr[15] m_wb_adr[16]
+ m_wb_adr[17] m_wb_adr[18] m_wb_adr[19] m_wb_adr[1] m_wb_adr[20] m_wb_adr[21] m_wb_adr[22]
+ m_wb_adr[23] m_wb_adr[2] m_wb_adr[3] m_wb_adr[4] m_wb_adr[5] m_wb_adr[6] m_wb_adr[7]
+ m_wb_adr[8] m_wb_adr[9] m_wb_cyc m_wb_err m_wb_i_dat[0] m_wb_i_dat[10] m_wb_i_dat[11]
+ m_wb_i_dat[12] m_wb_i_dat[13] m_wb_i_dat[14] m_wb_i_dat[15] m_wb_i_dat[1] m_wb_i_dat[2]
+ m_wb_i_dat[3] m_wb_i_dat[4] m_wb_i_dat[5] m_wb_i_dat[6] m_wb_i_dat[7] m_wb_i_dat[8]
+ m_wb_i_dat[9] m_wb_o_dat[0] m_wb_o_dat[10] m_wb_o_dat[11] m_wb_o_dat[12] m_wb_o_dat[13]
+ m_wb_o_dat[14] m_wb_o_dat[15] m_wb_o_dat[1] m_wb_o_dat[2] m_wb_o_dat[3] m_wb_o_dat[4]
+ m_wb_o_dat[5] m_wb_o_dat[6] m_wb_o_dat[7] m_wb_o_dat[8] m_wb_o_dat[9] m_wb_sel[0]
+ m_wb_sel[1] m_wb_stb m_wb_we s_rst s_wb_4_burst s_wb_8_burst s_wb_ack s_wb_adr[0]
+ s_wb_adr[10] s_wb_adr[11] s_wb_adr[12] s_wb_adr[13] s_wb_adr[14] s_wb_adr[15] s_wb_adr[16]
+ s_wb_adr[17] s_wb_adr[18] s_wb_adr[19] s_wb_adr[1] s_wb_adr[20] s_wb_adr[21] s_wb_adr[22]
+ s_wb_adr[23] s_wb_adr[2] s_wb_adr[3] s_wb_adr[4] s_wb_adr[5] s_wb_adr[6] s_wb_adr[7]
+ s_wb_adr[8] s_wb_adr[9] s_wb_cyc s_wb_err s_wb_i_dat[0] s_wb_i_dat[10] s_wb_i_dat[11]
+ s_wb_i_dat[12] s_wb_i_dat[13] s_wb_i_dat[14] s_wb_i_dat[15] s_wb_i_dat[1] s_wb_i_dat[2]
+ s_wb_i_dat[3] s_wb_i_dat[4] s_wb_i_dat[5] s_wb_i_dat[6] s_wb_i_dat[7] s_wb_i_dat[8]
+ s_wb_i_dat[9] s_wb_o_dat[0] s_wb_o_dat[10] s_wb_o_dat[11] s_wb_o_dat[12] s_wb_o_dat[13]
+ s_wb_o_dat[14] s_wb_o_dat[15] s_wb_o_dat[1] s_wb_o_dat[2] s_wb_o_dat[3] s_wb_o_dat[4]
+ s_wb_o_dat[5] s_wb_o_dat[6] s_wb_o_dat[7] s_wb_o_dat[8] s_wb_o_dat[9] s_wb_sel[0]
+ s_wb_sel[1] s_wb_stb s_wb_we vccd1 vssd1
.ends

* Black-box entry subcircuit for wb_compressor abstract view
.subckt wb_compressor cw_ack cw_dir cw_err cw_io_i[0] cw_io_i[10] cw_io_i[11] cw_io_i[12]
+ cw_io_i[13] cw_io_i[14] cw_io_i[15] cw_io_i[1] cw_io_i[2] cw_io_i[3] cw_io_i[4]
+ cw_io_i[5] cw_io_i[6] cw_io_i[7] cw_io_i[8] cw_io_i[9] cw_io_o[0] cw_io_o[10] cw_io_o[11]
+ cw_io_o[12] cw_io_o[13] cw_io_o[14] cw_io_o[15] cw_io_o[1] cw_io_o[2] cw_io_o[3]
+ cw_io_o[4] cw_io_o[5] cw_io_o[6] cw_io_o[7] cw_io_o[8] cw_io_o[9] cw_req i_clk i_rst
+ vccd1 vssd1 wb_4_burst wb_8_burst wb_ack wb_adr[0] wb_adr[10] wb_adr[11] wb_adr[12]
+ wb_adr[13] wb_adr[14] wb_adr[15] wb_adr[16] wb_adr[17] wb_adr[18] wb_adr[19] wb_adr[1]
+ wb_adr[20] wb_adr[21] wb_adr[22] wb_adr[23] wb_adr[2] wb_adr[3] wb_adr[4] wb_adr[5]
+ wb_adr[6] wb_adr[7] wb_adr[8] wb_adr[9] wb_cyc wb_err wb_i_dat[0] wb_i_dat[10] wb_i_dat[11]
+ wb_i_dat[12] wb_i_dat[13] wb_i_dat[14] wb_i_dat[15] wb_i_dat[1] wb_i_dat[2] wb_i_dat[3]
+ wb_i_dat[4] wb_i_dat[5] wb_i_dat[6] wb_i_dat[7] wb_i_dat[8] wb_i_dat[9] wb_o_dat[0]
+ wb_o_dat[10] wb_o_dat[11] wb_o_dat[12] wb_o_dat[13] wb_o_dat[14] wb_o_dat[15] wb_o_dat[1]
+ wb_o_dat[2] wb_o_dat[3] wb_o_dat[4] wb_o_dat[5] wb_o_dat[6] wb_o_dat[7] wb_o_dat[8]
+ wb_o_dat[9] wb_sel[0] wb_sel[1] wb_stb wb_we
.ends

* Black-box entry subcircuit for dcache abstract view
.subckt dcache i_clk i_rst mem_ack mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12]
+ mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[16] mem_addr[17] mem_addr[18] mem_addr[19]
+ mem_addr[1] mem_addr[20] mem_addr[21] mem_addr[22] mem_addr[23] mem_addr[2] mem_addr[3]
+ mem_addr[4] mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_cache_enable
+ mem_exception mem_i_data[0] mem_i_data[10] mem_i_data[11] mem_i_data[12] mem_i_data[13]
+ mem_i_data[14] mem_i_data[15] mem_i_data[1] mem_i_data[2] mem_i_data[3] mem_i_data[4]
+ mem_i_data[5] mem_i_data[6] mem_i_data[7] mem_i_data[8] mem_i_data[9] mem_o_data[0]
+ mem_o_data[10] mem_o_data[11] mem_o_data[12] mem_o_data[13] mem_o_data[14] mem_o_data[15]
+ mem_o_data[1] mem_o_data[2] mem_o_data[3] mem_o_data[4] mem_o_data[5] mem_o_data[6]
+ mem_o_data[7] mem_o_data[8] mem_o_data[9] mem_req mem_sel[0] mem_sel[1] mem_we vccd1
+ vssd1 wb_4_burst wb_ack wb_adr[0] wb_adr[10] wb_adr[11] wb_adr[12] wb_adr[13] wb_adr[14]
+ wb_adr[15] wb_adr[16] wb_adr[17] wb_adr[18] wb_adr[19] wb_adr[1] wb_adr[20] wb_adr[21]
+ wb_adr[22] wb_adr[23] wb_adr[2] wb_adr[3] wb_adr[4] wb_adr[5] wb_adr[6] wb_adr[7]
+ wb_adr[8] wb_adr[9] wb_cyc wb_err wb_i_dat[0] wb_i_dat[10] wb_i_dat[11] wb_i_dat[12]
+ wb_i_dat[13] wb_i_dat[14] wb_i_dat[15] wb_i_dat[1] wb_i_dat[2] wb_i_dat[3] wb_i_dat[4]
+ wb_i_dat[5] wb_i_dat[6] wb_i_dat[7] wb_i_dat[8] wb_i_dat[9] wb_o_dat[0] wb_o_dat[10]
+ wb_o_dat[11] wb_o_dat[12] wb_o_dat[13] wb_o_dat[14] wb_o_dat[15] wb_o_dat[1] wb_o_dat[2]
+ wb_o_dat[3] wb_o_dat[4] wb_o_dat[5] wb_o_dat[6] wb_o_dat[7] wb_o_dat[8] wb_o_dat[9]
+ wb_sel[0] wb_sel[1] wb_stb wb_we
.ends

* Black-box entry subcircuit for clk_div abstract view
.subckt clk_div clock_sel div[0] div[1] div[2] div[3] div_we i_clk i_rst o_clk vccd1
+ vssd1
.ends

* Black-box entry subcircuit for upper_core_logic abstract view
.subckt upper_core_logic cc_data_page cc_instr_page data_cacheable data_mem_addr[0]
+ data_mem_addr[10] data_mem_addr[11] data_mem_addr[12] data_mem_addr[13] data_mem_addr[14]
+ data_mem_addr[15] data_mem_addr[1] data_mem_addr[2] data_mem_addr[3] data_mem_addr[4]
+ data_mem_addr[5] data_mem_addr[6] data_mem_addr[7] data_mem_addr[8] data_mem_addr[9]
+ data_mem_addr_paged[0] data_mem_addr_paged[10] data_mem_addr_paged[11] data_mem_addr_paged[12]
+ data_mem_addr_paged[13] data_mem_addr_paged[14] data_mem_addr_paged[15] data_mem_addr_paged[16]
+ data_mem_addr_paged[17] data_mem_addr_paged[18] data_mem_addr_paged[19] data_mem_addr_paged[1]
+ data_mem_addr_paged[20] data_mem_addr_paged[21] data_mem_addr_paged[22] data_mem_addr_paged[23]
+ data_mem_addr_paged[2] data_mem_addr_paged[3] data_mem_addr_paged[4] data_mem_addr_paged[5]
+ data_mem_addr_paged[6] data_mem_addr_paged[7] data_mem_addr_paged[8] data_mem_addr_paged[9]
+ fetch_wb_adr[0] fetch_wb_adr[10] fetch_wb_adr[11] fetch_wb_adr[12] fetch_wb_adr[13]
+ fetch_wb_adr[14] fetch_wb_adr[15] fetch_wb_adr[1] fetch_wb_adr[2] fetch_wb_adr[3]
+ fetch_wb_adr[4] fetch_wb_adr[5] fetch_wb_adr[6] fetch_wb_adr[7] fetch_wb_adr[8]
+ fetch_wb_adr[9] fetch_wb_adr_paged[0] fetch_wb_adr_paged[10] fetch_wb_adr_paged[11]
+ fetch_wb_adr_paged[12] fetch_wb_adr_paged[13] fetch_wb_adr_paged[14] fetch_wb_adr_paged[15]
+ fetch_wb_adr_paged[16] fetch_wb_adr_paged[17] fetch_wb_adr_paged[18] fetch_wb_adr_paged[19]
+ fetch_wb_adr_paged[1] fetch_wb_adr_paged[20] fetch_wb_adr_paged[21] fetch_wb_adr_paged[22]
+ fetch_wb_adr_paged[23] fetch_wb_adr_paged[2] fetch_wb_adr_paged[3] fetch_wb_adr_paged[4]
+ fetch_wb_adr_paged[5] fetch_wb_adr_paged[6] fetch_wb_adr_paged[7] fetch_wb_adr_paged[8]
+ fetch_wb_adr_paged[9] fetch_wb_o_dat[0] fetch_wb_o_dat[10] fetch_wb_o_dat[11] fetch_wb_o_dat[12]
+ fetch_wb_o_dat[13] fetch_wb_o_dat[14] fetch_wb_o_dat[15] fetch_wb_o_dat[1] fetch_wb_o_dat[2]
+ fetch_wb_o_dat[3] fetch_wb_o_dat[4] fetch_wb_o_dat[5] fetch_wb_o_dat[6] fetch_wb_o_dat[7]
+ fetch_wb_o_dat[8] fetch_wb_o_dat[9] i_clk i_rst sr_bus_addr[0] sr_bus_addr[10] sr_bus_addr[11]
+ sr_bus_addr[12] sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15] sr_bus_addr[1] sr_bus_addr[2]
+ sr_bus_addr[3] sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6] sr_bus_addr[7] sr_bus_addr[8]
+ sr_bus_addr[9] sr_bus_data_o[0] sr_bus_data_o[10] sr_bus_data_o[11] sr_bus_data_o[12]
+ sr_bus_data_o[13] sr_bus_data_o[14] sr_bus_data_o[15] sr_bus_data_o[1] sr_bus_data_o[2]
+ sr_bus_data_o[3] sr_bus_data_o[4] sr_bus_data_o[5] sr_bus_data_o[6] sr_bus_data_o[7]
+ sr_bus_data_o[8] sr_bus_data_o[9] sr_bus_we vccd1 vssd1 wb0_8_burst wb1_4_burst
+ wb1_8_burst
.ends

* Black-box entry subcircuit for uprj_w_const abstract view
.subckt uprj_w_const b0_drv[0] b0_drv[10] b0_drv[11] b0_drv[12] b0_drv[13] b0_drv[14]
+ b0_drv[15] b0_drv[16] b0_drv[17] b0_drv[18] b0_drv[19] b0_drv[1] b0_drv[20] b0_drv[21]
+ b0_drv[22] b0_drv[23] b0_drv[24] b0_drv[25] b0_drv[26] b0_drv[27] b0_drv[28] b0_drv[29]
+ b0_drv[2] b0_drv[30] b0_drv[31] b0_drv[32] b0_drv[33] b0_drv[34] b0_drv[35] b0_drv[36]
+ b0_drv[37] b0_drv[38] b0_drv[39] b0_drv[3] b0_drv[40] b0_drv[41] b0_drv[42] b0_drv[43]
+ b0_drv[44] b0_drv[45] b0_drv[46] b0_drv[47] b0_drv[48] b0_drv[49] b0_drv[4] b0_drv[50]
+ b0_drv[51] b0_drv[52] b0_drv[53] b0_drv[54] b0_drv[55] b0_drv[56] b0_drv[57] b0_drv[58]
+ b0_drv[59] b0_drv[5] b0_drv[60] b0_drv[61] b0_drv[62] b0_drv[63] b0_drv[64] b0_drv[65]
+ b0_drv[66] b0_drv[67] b0_drv[68] b0_drv[69] b0_drv[6] b0_drv[70] b0_drv[71] b0_drv[72]
+ b0_drv[73] b0_drv[74] b0_drv[75] b0_drv[76] b0_drv[77] b0_drv[78] b0_drv[79] b0_drv[7]
+ b0_drv[80] b0_drv[81] b0_drv[82] b0_drv[8] b0_drv[9] cw_clk_i cw_clk_o cw_dir cw_dir_b_o
+ cw_dir_b_oo cw_dir_o cw_req_i cw_req_o cw_rst_i cw_rst_o i_pin_rst i_wb_rst io_oeb_15_0[0]
+ io_oeb_15_0[10] io_oeb_15_0[11] io_oeb_15_0[12] io_oeb_15_0[13] io_oeb_15_0[14]
+ io_oeb_15_0[15] io_oeb_15_0[1] io_oeb_15_0[2] io_oeb_15_0[3] io_oeb_15_0[4] io_oeb_15_0[5]
+ io_oeb_15_0[6] io_oeb_15_0[7] io_oeb_15_0[8] io_oeb_15_0[9] io_oeb_18_16[0] io_oeb_18_16[1]
+ io_oeb_18_16[2] io_oeb_20_19[0] io_oeb_20_19[1] io_oeb_21 io_oeb_22 io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[1] io_out[2] io_out[3] io_out[4]
+ io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] io_out_20_19[0] io_out_20_19[1]
+ io_out_22 la_data_out_16_17[0] la_data_out_16_17[1] la_data_out_21 la_data_out_37_36[0]
+ la_data_out_37_36[1] la_data_out_77_62[0] la_data_out_77_62[10] la_data_out_77_62[11]
+ la_data_out_77_62[12] la_data_out_77_62[13] la_data_out_77_62[14] la_data_out_77_62[15]
+ la_data_out_77_62[1] la_data_out_77_62[2] la_data_out_77_62[3] la_data_out_77_62[4]
+ la_data_out_77_62[5] la_data_out_77_62[6] la_data_out_77_62[7] la_data_out_77_62[8]
+ la_data_out_77_62[9] la_data_out_97_95[0] la_data_out_97_95[1] la_data_out_97_95[2]
+ la_datb_i[0] la_datb_i[1] la_datb_i[2] la_datb_o[0] la_datb_o[1] la_datb_o[2] o_s_rst
+ oeb_out[0] oeb_out[10] oeb_out[11] oeb_out[12] oeb_out[13] oeb_out[14] oeb_out[1]
+ oeb_out[2] oeb_out[3] oeb_out[4] oeb_out[5] oeb_out[6] oeb_out[7] oeb_out[8] oeb_out[9]
+ soft_rst vccd1 vssd1
.ends

* Black-box entry subcircuit for top_cw_logic abstract view
.subckt top_cw_logic c_wb_4_burst c_wb_8_burst c_wb_ack_cmp c_wb_adr[0] c_wb_adr[10]
+ c_wb_adr[11] c_wb_adr[12] c_wb_adr[13] c_wb_adr[14] c_wb_adr[15] c_wb_adr[16] c_wb_adr[17]
+ c_wb_adr[18] c_wb_adr[19] c_wb_adr[1] c_wb_adr[20] c_wb_adr[21] c_wb_adr[22] c_wb_adr[23]
+ c_wb_adr[2] c_wb_adr[3] c_wb_adr[4] c_wb_adr[5] c_wb_adr[6] c_wb_adr[7] c_wb_adr[8]
+ c_wb_adr[9] c_wb_cyc c_wb_err_cmp c_wb_i_dat_cmp[0] c_wb_i_dat_cmp[10] c_wb_i_dat_cmp[11]
+ c_wb_i_dat_cmp[12] c_wb_i_dat_cmp[13] c_wb_i_dat_cmp[14] c_wb_i_dat_cmp[15] c_wb_i_dat_cmp[1]
+ c_wb_i_dat_cmp[2] c_wb_i_dat_cmp[3] c_wb_i_dat_cmp[4] c_wb_i_dat_cmp[5] c_wb_i_dat_cmp[6]
+ c_wb_i_dat_cmp[7] c_wb_i_dat_cmp[8] c_wb_i_dat_cmp[9] c_wb_o_dat[0] c_wb_o_dat[10]
+ c_wb_o_dat[11] c_wb_o_dat[12] c_wb_o_dat[13] c_wb_o_dat[14] c_wb_o_dat[15] c_wb_o_dat[1]
+ c_wb_o_dat[2] c_wb_o_dat[3] c_wb_o_dat[4] c_wb_o_dat[5] c_wb_o_dat[6] c_wb_o_dat[7]
+ c_wb_o_dat[8] c_wb_o_dat[9] c_wb_sel[0] c_wb_sel[1] c_wb_stb c_wb_we cc_wb_4_burst
+ cc_wb_8_burst cc_wb_adr[0] cc_wb_adr[10] cc_wb_adr[11] cc_wb_adr[12] cc_wb_adr[13]
+ cc_wb_adr[14] cc_wb_adr[15] cc_wb_adr[16] cc_wb_adr[17] cc_wb_adr[18] cc_wb_adr[19]
+ cc_wb_adr[1] cc_wb_adr[20] cc_wb_adr[21] cc_wb_adr[22] cc_wb_adr[23] cc_wb_adr[2]
+ cc_wb_adr[3] cc_wb_adr[4] cc_wb_adr[5] cc_wb_adr[6] cc_wb_adr[7] cc_wb_adr[8] cc_wb_adr[9]
+ cc_wb_cyc cc_wb_o_dat[0] cc_wb_o_dat[10] cc_wb_o_dat[11] cc_wb_o_dat[12] cc_wb_o_dat[13]
+ cc_wb_o_dat[14] cc_wb_o_dat[15] cc_wb_o_dat[1] cc_wb_o_dat[2] cc_wb_o_dat[3] cc_wb_o_dat[4]
+ cc_wb_o_dat[5] cc_wb_o_dat[6] cc_wb_o_dat[7] cc_wb_o_dat[8] cc_wb_o_dat[9] cc_wb_sel[0]
+ cc_wb_sel[1] cc_wb_stb cc_wb_we cw_ack cw_clk cw_err cw_io_i[0] cw_io_i[10] cw_io_i[11]
+ cw_io_i[12] cw_io_i[13] cw_io_i[14] cw_io_i[15] cw_io_i[1] cw_io_i[2] cw_io_i[3]
+ cw_io_i[4] cw_io_i[5] cw_io_i[6] cw_io_i[7] cw_io_i[8] cw_io_i[9] cw_rst cw_rst_z
+ i_clk i_irq i_rst ic_split_clock irq_s la_cw_ack la_cw_io_i[0] la_cw_io_i[10] la_cw_io_i[11]
+ la_cw_io_i[12] la_cw_io_i[13] la_cw_io_i[14] la_cw_io_i[15] la_cw_io_i[1] la_cw_io_i[2]
+ la_cw_io_i[3] la_cw_io_i[4] la_cw_io_i[5] la_cw_io_i[6] la_cw_io_i[7] la_cw_io_i[8]
+ la_cw_io_i[9] la_cw_ovr m_cw_ack m_cw_err m_cw_io_i[0] m_cw_io_i[10] m_cw_io_i[11]
+ m_cw_io_i[12] m_cw_io_i[13] m_cw_io_i[14] m_cw_io_i[15] m_cw_io_i[1] m_cw_io_i[2]
+ m_cw_io_i[3] m_cw_io_i[4] m_cw_io_i[5] m_cw_io_i[6] m_cw_io_i[7] m_cw_io_i[8] m_cw_io_i[9]
+ s_rst u_wb_4_burst u_wb_8_burst u_wb_ack u_wb_ack_cc u_wb_ack_clk u_wb_ack_mxed
+ u_wb_adr[0] u_wb_adr[10] u_wb_adr[11] u_wb_adr[12] u_wb_adr[13] u_wb_adr[14] u_wb_adr[15]
+ u_wb_adr[16] u_wb_adr[17] u_wb_adr[18] u_wb_adr[19] u_wb_adr[1] u_wb_adr[20] u_wb_adr[21]
+ u_wb_adr[22] u_wb_adr[23] u_wb_adr[2] u_wb_adr[3] u_wb_adr[4] u_wb_adr[5] u_wb_adr[6]
+ u_wb_adr[7] u_wb_adr[8] u_wb_adr[9] u_wb_cyc u_wb_err u_wb_err_cc u_wb_i_dat[0]
+ u_wb_i_dat[10] u_wb_i_dat[11] u_wb_i_dat[12] u_wb_i_dat[13] u_wb_i_dat[14] u_wb_i_dat[15]
+ u_wb_i_dat[1] u_wb_i_dat[2] u_wb_i_dat[3] u_wb_i_dat[4] u_wb_i_dat[5] u_wb_i_dat[6]
+ u_wb_i_dat[7] u_wb_i_dat[8] u_wb_i_dat[9] u_wb_i_dat_cc[0] u_wb_i_dat_cc[10] u_wb_i_dat_cc[11]
+ u_wb_i_dat_cc[12] u_wb_i_dat_cc[13] u_wb_i_dat_cc[14] u_wb_i_dat_cc[15] u_wb_i_dat_cc[1]
+ u_wb_i_dat_cc[2] u_wb_i_dat_cc[3] u_wb_i_dat_cc[4] u_wb_i_dat_cc[5] u_wb_i_dat_cc[6]
+ u_wb_i_dat_cc[7] u_wb_i_dat_cc[8] u_wb_i_dat_cc[9] u_wb_o_dat[0] u_wb_o_dat[10]
+ u_wb_o_dat[11] u_wb_o_dat[12] u_wb_o_dat[13] u_wb_o_dat[14] u_wb_o_dat[15] u_wb_o_dat[1]
+ u_wb_o_dat[2] u_wb_o_dat[3] u_wb_o_dat[4] u_wb_o_dat[5] u_wb_o_dat[6] u_wb_o_dat[7]
+ u_wb_o_dat[8] u_wb_o_dat[9] u_wb_sel[0] u_wb_sel[1] u_wb_stb u_wb_we vccd1 vssd1
.ends

* Black-box entry subcircuit for wishbone_arbiter abstract view
.subckt wishbone_arbiter i_clk i_rst i_wb0_cyc i_wb1_cyc o_sel_sig o_wb_cyc owb_4_burst
+ owb_8_burst owb_ack owb_adr[0] owb_adr[10] owb_adr[11] owb_adr[12] owb_adr[13] owb_adr[14]
+ owb_adr[15] owb_adr[16] owb_adr[17] owb_adr[18] owb_adr[19] owb_adr[1] owb_adr[20]
+ owb_adr[21] owb_adr[22] owb_adr[23] owb_adr[2] owb_adr[3] owb_adr[4] owb_adr[5]
+ owb_adr[6] owb_adr[7] owb_adr[8] owb_adr[9] owb_err owb_o_dat[0] owb_o_dat[10] owb_o_dat[11]
+ owb_o_dat[12] owb_o_dat[13] owb_o_dat[14] owb_o_dat[15] owb_o_dat[1] owb_o_dat[2]
+ owb_o_dat[3] owb_o_dat[4] owb_o_dat[5] owb_o_dat[6] owb_o_dat[7] owb_o_dat[8] owb_o_dat[9]
+ owb_sel[0] owb_sel[1] owb_stb owb_we vccd1 vssd1 wb0_4_burst wb0_8_burst wb0_ack
+ wb0_adr[0] wb0_adr[10] wb0_adr[11] wb0_adr[12] wb0_adr[13] wb0_adr[14] wb0_adr[15]
+ wb0_adr[16] wb0_adr[17] wb0_adr[18] wb0_adr[19] wb0_adr[1] wb0_adr[20] wb0_adr[21]
+ wb0_adr[22] wb0_adr[23] wb0_adr[2] wb0_adr[3] wb0_adr[4] wb0_adr[5] wb0_adr[6] wb0_adr[7]
+ wb0_adr[8] wb0_adr[9] wb0_err wb0_o_dat[0] wb0_o_dat[10] wb0_o_dat[11] wb0_o_dat[12]
+ wb0_o_dat[13] wb0_o_dat[14] wb0_o_dat[15] wb0_o_dat[1] wb0_o_dat[2] wb0_o_dat[3]
+ wb0_o_dat[4] wb0_o_dat[5] wb0_o_dat[6] wb0_o_dat[7] wb0_o_dat[8] wb0_o_dat[9] wb0_sel[0]
+ wb0_sel[1] wb0_stb wb0_we wb1_4_burst wb1_8_burst wb1_ack wb1_adr[0] wb1_adr[10]
+ wb1_adr[11] wb1_adr[12] wb1_adr[13] wb1_adr[14] wb1_adr[15] wb1_adr[16] wb1_adr[17]
+ wb1_adr[18] wb1_adr[19] wb1_adr[1] wb1_adr[20] wb1_adr[21] wb1_adr[22] wb1_adr[23]
+ wb1_adr[2] wb1_adr[3] wb1_adr[4] wb1_adr[5] wb1_adr[6] wb1_adr[7] wb1_adr[8] wb1_adr[9]
+ wb1_err wb1_o_dat[0] wb1_o_dat[10] wb1_o_dat[11] wb1_o_dat[12] wb1_o_dat[13] wb1_o_dat[14]
+ wb1_o_dat[15] wb1_o_dat[1] wb1_o_dat[2] wb1_o_dat[3] wb1_o_dat[4] wb1_o_dat[5] wb1_o_dat[6]
+ wb1_o_dat[7] wb1_o_dat[8] wb1_o_dat[9] wb1_sel[0] wb1_sel[1] wb1_stb wb1_we
.ends

* Black-box entry subcircuit for icache abstract view
.subckt icache i_clk i_rst mem_ack mem_addr[0] mem_addr[10] mem_addr[11] mem_addr[12]
+ mem_addr[13] mem_addr[14] mem_addr[15] mem_addr[1] mem_addr[2] mem_addr[3] mem_addr[4]
+ mem_addr[5] mem_addr[6] mem_addr[7] mem_addr[8] mem_addr[9] mem_cache_flush mem_data[0]
+ mem_data[10] mem_data[11] mem_data[12] mem_data[13] mem_data[14] mem_data[15] mem_data[16]
+ mem_data[17] mem_data[18] mem_data[19] mem_data[1] mem_data[20] mem_data[21] mem_data[22]
+ mem_data[23] mem_data[24] mem_data[25] mem_data[26] mem_data[27] mem_data[28] mem_data[29]
+ mem_data[2] mem_data[30] mem_data[31] mem_data[3] mem_data[4] mem_data[5] mem_data[6]
+ mem_data[7] mem_data[8] mem_data[9] mem_ppl_submit mem_req vccd1 vssd1 wb_ack wb_adr[0]
+ wb_adr[10] wb_adr[11] wb_adr[12] wb_adr[13] wb_adr[14] wb_adr[15] wb_adr[1] wb_adr[2]
+ wb_adr[3] wb_adr[4] wb_adr[5] wb_adr[6] wb_adr[7] wb_adr[8] wb_adr[9] wb_cyc wb_err
+ wb_i_dat[0] wb_i_dat[10] wb_i_dat[11] wb_i_dat[12] wb_i_dat[13] wb_i_dat[14] wb_i_dat[15]
+ wb_i_dat[1] wb_i_dat[2] wb_i_dat[3] wb_i_dat[4] wb_i_dat[5] wb_i_dat[6] wb_i_dat[7]
+ wb_i_dat[8] wb_i_dat[9] wb_sel[0] wb_sel[1] wb_stb wb_we
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xtop_cw.upc.core la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_out[0]
+ la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] uprj_w_const/la_datb_i[2] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] top_cw.upc.core/dbg_pc[0] top_cw.upc.core/dbg_pc[10]
+ top_cw.upc.core/dbg_pc[11] top_cw.upc.core/dbg_pc[12] top_cw.upc.core/dbg_pc[13]
+ top_cw.upc.core/dbg_pc[14] top_cw.upc.core/dbg_pc[15] top_cw.upc.core/dbg_pc[1]
+ top_cw.upc.core/dbg_pc[2] top_cw.upc.core/dbg_pc[3] top_cw.upc.core/dbg_pc[4] top_cw.upc.core/dbg_pc[5]
+ top_cw.upc.core/dbg_pc[6] top_cw.upc.core/dbg_pc[7] top_cw.upc.core/dbg_pc[8] top_cw.upc.core/dbg_pc[9]
+ top_cw.upc.core/dbg_r0[0] top_cw.upc.core/dbg_r0[10] top_cw.upc.core/dbg_r0[11]
+ top_cw.upc.core/dbg_r0[12] top_cw.upc.core/dbg_r0[13] top_cw.upc.core/dbg_r0[14]
+ top_cw.upc.core/dbg_r0[15] top_cw.upc.core/dbg_r0[1] top_cw.upc.core/dbg_r0[2] top_cw.upc.core/dbg_r0[3]
+ top_cw.upc.core/dbg_r0[4] top_cw.upc.core/dbg_r0[5] top_cw.upc.core/dbg_r0[6] top_cw.upc.core/dbg_r0[7]
+ top_cw.upc.core/dbg_r0[8] top_cw.upc.core/dbg_r0[9] user_clock2 top_cw.upc.core/i_irq
+ top_cw.upc.dcache/mem_ack top_cw.upc.core/i_mem_data[0] top_cw.upc.core/i_mem_data[10]
+ top_cw.upc.core/i_mem_data[11] top_cw.upc.core/i_mem_data[12] top_cw.upc.core/i_mem_data[13]
+ top_cw.upc.core/i_mem_data[14] top_cw.upc.core/i_mem_data[15] top_cw.upc.core/i_mem_data[1]
+ top_cw.upc.core/i_mem_data[2] top_cw.upc.core/i_mem_data[3] top_cw.upc.core/i_mem_data[4]
+ top_cw.upc.core/i_mem_data[5] top_cw.upc.core/i_mem_data[6] top_cw.upc.core/i_mem_data[7]
+ top_cw.upc.core/i_mem_data[8] top_cw.upc.core/i_mem_data[9] top_cw.upc.dcache/mem_exception
+ top_cw.upc.icache/mem_data[0] top_cw.upc.icache/mem_data[10] top_cw.upc.icache/mem_data[11]
+ top_cw.upc.icache/mem_data[12] top_cw.upc.icache/mem_data[13] top_cw.upc.icache/mem_data[14]
+ top_cw.upc.icache/mem_data[15] top_cw.upc.icache/mem_data[16] top_cw.upc.icache/mem_data[17]
+ top_cw.upc.icache/mem_data[18] top_cw.upc.icache/mem_data[19] top_cw.upc.icache/mem_data[1]
+ top_cw.upc.icache/mem_data[20] top_cw.upc.icache/mem_data[21] top_cw.upc.icache/mem_data[22]
+ top_cw.upc.icache/mem_data[23] top_cw.upc.icache/mem_data[24] top_cw.upc.icache/mem_data[25]
+ top_cw.upc.icache/mem_data[26] top_cw.upc.icache/mem_data[27] top_cw.upc.icache/mem_data[28]
+ top_cw.upc.icache/mem_data[29] top_cw.upc.icache/mem_data[2] top_cw.upc.icache/mem_data[30]
+ top_cw.upc.icache/mem_data[31] top_cw.upc.icache/mem_data[3] top_cw.upc.icache/mem_data[4]
+ top_cw.upc.icache/mem_data[5] top_cw.upc.icache/mem_data[6] top_cw.upc.icache/mem_data[7]
+ top_cw.upc.icache/mem_data[8] top_cw.upc.icache/mem_data[9] top_cw.upc.icache/mem_ack
+ top_cw.clk_div/i_rst top_cw.upc.core/o_c_data_page top_cw.upc.core/o_c_instr_page
+ top_cw.upc.core/o_icache_flush top_cw.upc.core/o_mem_addr[0] top_cw.upc.core/o_mem_addr[10]
+ top_cw.upc.core/o_mem_addr[11] top_cw.upc.core/o_mem_addr[12] top_cw.upc.core/o_mem_addr[13]
+ top_cw.upc.core/o_mem_addr[14] top_cw.upc.core/o_mem_addr[15] top_cw.upc.core/o_mem_addr[1]
+ top_cw.upc.core/o_mem_addr[2] top_cw.upc.core/o_mem_addr[3] top_cw.upc.core/o_mem_addr[4]
+ top_cw.upc.core/o_mem_addr[5] top_cw.upc.core/o_mem_addr[6] top_cw.upc.core/o_mem_addr[7]
+ top_cw.upc.core/o_mem_addr[8] top_cw.upc.core/o_mem_addr[9] top_cw.upc.core/o_mem_data[0]
+ top_cw.upc.core/o_mem_data[10] top_cw.upc.core/o_mem_data[11] top_cw.upc.core/o_mem_data[12]
+ top_cw.upc.core/o_mem_data[13] top_cw.upc.core/o_mem_data[14] top_cw.upc.core/o_mem_data[15]
+ top_cw.upc.core/o_mem_data[1] top_cw.upc.core/o_mem_data[2] top_cw.upc.core/o_mem_data[3]
+ top_cw.upc.core/o_mem_data[4] top_cw.upc.core/o_mem_data[5] top_cw.upc.core/o_mem_data[6]
+ top_cw.upc.core/o_mem_data[7] top_cw.upc.core/o_mem_data[8] top_cw.upc.core/o_mem_data[9]
+ top_cw.upc.dcache/mem_req top_cw.upc.dcache/mem_sel[0] top_cw.upc.dcache/mem_sel[1]
+ top_cw.upc.dcache/mem_we top_cw.upc.icache/mem_req top_cw.upc.icache/mem_addr[0]
+ top_cw.upc.icache/mem_addr[10] top_cw.upc.icache/mem_addr[11] top_cw.upc.icache/mem_addr[12]
+ top_cw.upc.icache/mem_addr[13] top_cw.upc.icache/mem_addr[14] top_cw.upc.icache/mem_addr[15]
+ top_cw.upc.icache/mem_addr[1] top_cw.upc.icache/mem_addr[2] top_cw.upc.icache/mem_addr[3]
+ top_cw.upc.icache/mem_addr[4] top_cw.upc.icache/mem_addr[5] top_cw.upc.icache/mem_addr[6]
+ top_cw.upc.icache/mem_addr[7] top_cw.upc.icache/mem_addr[8] top_cw.upc.icache/mem_addr[9]
+ top_cw.upc.icache/mem_ppl_submit top_cw.upc.core/sr_bus_addr[0] top_cw.upc.core/sr_bus_addr[10]
+ top_cw.upc.core/sr_bus_addr[11] top_cw.upc.core/sr_bus_addr[12] top_cw.upc.core/sr_bus_addr[13]
+ top_cw.upc.core/sr_bus_addr[14] top_cw.upc.core/sr_bus_addr[15] top_cw.upc.core/sr_bus_addr[1]
+ top_cw.upc.core/sr_bus_addr[2] top_cw.upc.core/sr_bus_addr[3] top_cw.upc.core/sr_bus_addr[4]
+ top_cw.upc.core/sr_bus_addr[5] top_cw.upc.core/sr_bus_addr[6] top_cw.upc.core/sr_bus_addr[7]
+ top_cw.upc.core/sr_bus_addr[8] top_cw.upc.core/sr_bus_addr[9] top_cw.upc.core/sr_bus_data_o[0]
+ top_cw.upc.core/sr_bus_data_o[10] top_cw.upc.core/sr_bus_data_o[11] top_cw.upc.core/sr_bus_data_o[12]
+ top_cw.upc.core/sr_bus_data_o[13] top_cw.upc.core/sr_bus_data_o[14] top_cw.upc.core/sr_bus_data_o[15]
+ top_cw.upc.core/sr_bus_data_o[1] top_cw.upc.core/sr_bus_data_o[2] top_cw.upc.core/sr_bus_data_o[3]
+ top_cw.upc.core/sr_bus_data_o[4] top_cw.upc.core/sr_bus_data_o[5] top_cw.upc.core/sr_bus_data_o[6]
+ top_cw.upc.core/sr_bus_data_o[7] top_cw.upc.core/sr_bus_data_o[8] top_cw.upc.core/sr_bus_data_o[9]
+ top_cw.upc.core/sr_bus_we vccd1 vssd1 core
Xtop_cw.wb_cross_clk user_clock2 top_cw.clk_div/o_clk top_cw.clk_div/i_rst top_cw.wb_cross_clk/m_wb_4_burst
+ top_cw.wb_cross_clk/m_wb_8_burst top_cw.wb_cross_clk/m_wb_ack la_data_out[38] la_data_out[48]
+ la_data_out[49] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[39]
+ la_data_out[58] la_data_out[59] la_data_out[60] la_data_out[61] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] top_cw.wb_cross_clk/m_wb_cyc top_cw.wb_cross_clk/m_wb_err
+ top_cw.wb_cross_clk/m_wb_i_dat[0] top_cw.wb_cross_clk/m_wb_i_dat[10] top_cw.wb_cross_clk/m_wb_i_dat[11]
+ top_cw.wb_cross_clk/m_wb_i_dat[12] top_cw.wb_cross_clk/m_wb_i_dat[13] top_cw.wb_cross_clk/m_wb_i_dat[14]
+ top_cw.wb_cross_clk/m_wb_i_dat[15] top_cw.wb_cross_clk/m_wb_i_dat[1] top_cw.wb_cross_clk/m_wb_i_dat[2]
+ top_cw.wb_cross_clk/m_wb_i_dat[3] top_cw.wb_cross_clk/m_wb_i_dat[4] top_cw.wb_cross_clk/m_wb_i_dat[5]
+ top_cw.wb_cross_clk/m_wb_i_dat[6] top_cw.wb_cross_clk/m_wb_i_dat[7] top_cw.wb_cross_clk/m_wb_i_dat[8]
+ top_cw.wb_cross_clk/m_wb_i_dat[9] top_cw.clk_div/div[0] top_cw.wb_cross_clk/m_wb_o_dat[10]
+ top_cw.wb_cross_clk/m_wb_o_dat[11] top_cw.wb_cross_clk/m_wb_o_dat[12] top_cw.wb_cross_clk/m_wb_o_dat[13]
+ top_cw.wb_cross_clk/m_wb_o_dat[14] top_cw.wb_cross_clk/m_wb_o_dat[15] top_cw.clk_div/div[1]
+ top_cw.clk_div/div[2] top_cw.clk_div/div[3] top_cw.wb_cross_clk/m_wb_o_dat[4] top_cw.wb_cross_clk/m_wb_o_dat[5]
+ top_cw.wb_cross_clk/m_wb_o_dat[6] top_cw.wb_cross_clk/m_wb_o_dat[7] top_cw.wb_cross_clk/m_wb_o_dat[8]
+ top_cw.wb_cross_clk/m_wb_o_dat[9] top_cw.wb_cross_clk/m_wb_sel[0] top_cw.wb_cross_clk/m_wb_sel[1]
+ uprj_w_const/la_datb_i[0] uprj_w_const/la_datb_i[1] uprj_w_const/cw_rst_i top_cw.wb_cross_clk/s_wb_4_burst
+ top_cw.wb_cross_clk/s_wb_8_burst top_cw.wb_compressor/wb_ack top_cw.wb_cross_clk/s_wb_adr[0]
+ top_cw.wb_cross_clk/s_wb_adr[10] top_cw.wb_cross_clk/s_wb_adr[11] top_cw.wb_cross_clk/s_wb_adr[12]
+ top_cw.wb_cross_clk/s_wb_adr[13] top_cw.wb_cross_clk/s_wb_adr[14] top_cw.wb_cross_clk/s_wb_adr[15]
+ top_cw.wb_cross_clk/s_wb_adr[16] top_cw.wb_cross_clk/s_wb_adr[17] top_cw.wb_cross_clk/s_wb_adr[18]
+ top_cw.wb_cross_clk/s_wb_adr[19] top_cw.wb_cross_clk/s_wb_adr[1] top_cw.wb_cross_clk/s_wb_adr[20]
+ top_cw.wb_cross_clk/s_wb_adr[21] top_cw.wb_cross_clk/s_wb_adr[22] top_cw.wb_cross_clk/s_wb_adr[23]
+ top_cw.wb_cross_clk/s_wb_adr[2] top_cw.wb_cross_clk/s_wb_adr[3] top_cw.wb_cross_clk/s_wb_adr[4]
+ top_cw.wb_cross_clk/s_wb_adr[5] top_cw.wb_cross_clk/s_wb_adr[6] top_cw.wb_cross_clk/s_wb_adr[7]
+ top_cw.wb_cross_clk/s_wb_adr[8] top_cw.wb_cross_clk/s_wb_adr[9] top_cw.wb_cross_clk/s_wb_cyc
+ top_cw.wb_compressor/wb_err top_cw.wb_compressor/wb_i_dat[0] top_cw.wb_compressor/wb_i_dat[10]
+ top_cw.wb_compressor/wb_i_dat[11] top_cw.wb_compressor/wb_i_dat[12] top_cw.wb_compressor/wb_i_dat[13]
+ top_cw.wb_compressor/wb_i_dat[14] top_cw.wb_compressor/wb_i_dat[15] top_cw.wb_compressor/wb_i_dat[1]
+ top_cw.wb_compressor/wb_i_dat[2] top_cw.wb_compressor/wb_i_dat[3] top_cw.wb_compressor/wb_i_dat[4]
+ top_cw.wb_compressor/wb_i_dat[5] top_cw.wb_compressor/wb_i_dat[6] top_cw.wb_compressor/wb_i_dat[7]
+ top_cw.wb_compressor/wb_i_dat[8] top_cw.wb_compressor/wb_i_dat[9] top_cw.wb_cross_clk/s_wb_o_dat[0]
+ top_cw.wb_cross_clk/s_wb_o_dat[10] top_cw.wb_cross_clk/s_wb_o_dat[11] top_cw.wb_cross_clk/s_wb_o_dat[12]
+ top_cw.wb_cross_clk/s_wb_o_dat[13] top_cw.wb_cross_clk/s_wb_o_dat[14] top_cw.wb_cross_clk/s_wb_o_dat[15]
+ top_cw.wb_cross_clk/s_wb_o_dat[1] top_cw.wb_cross_clk/s_wb_o_dat[2] top_cw.wb_cross_clk/s_wb_o_dat[3]
+ top_cw.wb_cross_clk/s_wb_o_dat[4] top_cw.wb_cross_clk/s_wb_o_dat[5] top_cw.wb_cross_clk/s_wb_o_dat[6]
+ top_cw.wb_cross_clk/s_wb_o_dat[7] top_cw.wb_cross_clk/s_wb_o_dat[8] top_cw.wb_cross_clk/s_wb_o_dat[9]
+ top_cw.wb_cross_clk/s_wb_sel[0] top_cw.wb_cross_clk/s_wb_sel[1] top_cw.wb_cross_clk/s_wb_stb
+ top_cw.wb_cross_clk/s_wb_we vccd1 vssd1 wb_cross_clk
Xtop_cw.wb_compressor top_cw.wb_compressor/cw_ack uprj_w_const/cw_dir top_cw.wb_compressor/cw_err
+ top_cw.wb_compressor/cw_io_i[0] top_cw.wb_compressor/cw_io_i[10] top_cw.wb_compressor/cw_io_i[11]
+ top_cw.wb_compressor/cw_io_i[12] top_cw.wb_compressor/cw_io_i[13] top_cw.wb_compressor/cw_io_i[14]
+ top_cw.wb_compressor/cw_io_i[15] top_cw.wb_compressor/cw_io_i[1] top_cw.wb_compressor/cw_io_i[2]
+ top_cw.wb_compressor/cw_io_i[3] top_cw.wb_compressor/cw_io_i[4] top_cw.wb_compressor/cw_io_i[5]
+ top_cw.wb_compressor/cw_io_i[6] top_cw.wb_compressor/cw_io_i[7] top_cw.wb_compressor/cw_io_i[8]
+ top_cw.wb_compressor/cw_io_i[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] uprj_w_const/cw_req_i top_cw.clk_div/o_clk uprj_w_const/cw_rst_i
+ vccd1 vssd1 top_cw.wb_compressor/wb_4_burst top_cw.wb_compressor/wb_8_burst top_cw.wb_compressor/wb_ack
+ top_cw.wb_compressor/wb_adr[0] top_cw.wb_compressor/wb_adr[10] top_cw.wb_compressor/wb_adr[11]
+ top_cw.wb_compressor/wb_adr[12] top_cw.wb_compressor/wb_adr[13] top_cw.wb_compressor/wb_adr[14]
+ top_cw.wb_compressor/wb_adr[15] top_cw.wb_compressor/wb_adr[16] top_cw.wb_compressor/wb_adr[17]
+ top_cw.wb_compressor/wb_adr[18] top_cw.wb_compressor/wb_adr[19] top_cw.wb_compressor/wb_adr[1]
+ top_cw.wb_compressor/wb_adr[20] top_cw.wb_compressor/wb_adr[21] top_cw.wb_compressor/wb_adr[22]
+ top_cw.wb_compressor/wb_adr[23] top_cw.wb_compressor/wb_adr[2] top_cw.wb_compressor/wb_adr[3]
+ top_cw.wb_compressor/wb_adr[4] top_cw.wb_compressor/wb_adr[5] top_cw.wb_compressor/wb_adr[6]
+ top_cw.wb_compressor/wb_adr[7] top_cw.wb_compressor/wb_adr[8] top_cw.wb_compressor/wb_adr[9]
+ top_cw.wb_compressor/wb_cyc top_cw.wb_compressor/wb_err top_cw.wb_compressor/wb_i_dat[0]
+ top_cw.wb_compressor/wb_i_dat[10] top_cw.wb_compressor/wb_i_dat[11] top_cw.wb_compressor/wb_i_dat[12]
+ top_cw.wb_compressor/wb_i_dat[13] top_cw.wb_compressor/wb_i_dat[14] top_cw.wb_compressor/wb_i_dat[15]
+ top_cw.wb_compressor/wb_i_dat[1] top_cw.wb_compressor/wb_i_dat[2] top_cw.wb_compressor/wb_i_dat[3]
+ top_cw.wb_compressor/wb_i_dat[4] top_cw.wb_compressor/wb_i_dat[5] top_cw.wb_compressor/wb_i_dat[6]
+ top_cw.wb_compressor/wb_i_dat[7] top_cw.wb_compressor/wb_i_dat[8] top_cw.wb_compressor/wb_i_dat[9]
+ top_cw.wb_compressor/wb_o_dat[0] top_cw.wb_compressor/wb_o_dat[10] top_cw.wb_compressor/wb_o_dat[11]
+ top_cw.wb_compressor/wb_o_dat[12] top_cw.wb_compressor/wb_o_dat[13] top_cw.wb_compressor/wb_o_dat[14]
+ top_cw.wb_compressor/wb_o_dat[15] top_cw.wb_compressor/wb_o_dat[1] top_cw.wb_compressor/wb_o_dat[2]
+ top_cw.wb_compressor/wb_o_dat[3] top_cw.wb_compressor/wb_o_dat[4] top_cw.wb_compressor/wb_o_dat[5]
+ top_cw.wb_compressor/wb_o_dat[6] top_cw.wb_compressor/wb_o_dat[7] top_cw.wb_compressor/wb_o_dat[8]
+ top_cw.wb_compressor/wb_o_dat[9] top_cw.wb_compressor/wb_sel[0] top_cw.wb_compressor/wb_sel[1]
+ top_cw.wb_compressor/wb_stb top_cw.wb_compressor/wb_we wb_compressor
Xtop_cw.upc.dcache user_clock2 top_cw.clk_div/i_rst top_cw.upc.dcache/mem_ack top_cw.upc.dcache/mem_addr[0]
+ top_cw.upc.dcache/mem_addr[10] top_cw.upc.dcache/mem_addr[11] top_cw.upc.dcache/mem_addr[12]
+ top_cw.upc.dcache/mem_addr[13] top_cw.upc.dcache/mem_addr[14] top_cw.upc.dcache/mem_addr[15]
+ top_cw.upc.dcache/mem_addr[16] top_cw.upc.dcache/mem_addr[17] top_cw.upc.dcache/mem_addr[18]
+ top_cw.upc.dcache/mem_addr[19] top_cw.upc.dcache/mem_addr[1] top_cw.upc.dcache/mem_addr[20]
+ top_cw.upc.dcache/mem_addr[21] top_cw.upc.dcache/mem_addr[22] top_cw.upc.dcache/mem_addr[23]
+ top_cw.upc.dcache/mem_addr[2] top_cw.upc.dcache/mem_addr[3] top_cw.upc.dcache/mem_addr[4]
+ top_cw.upc.dcache/mem_addr[5] top_cw.upc.dcache/mem_addr[6] top_cw.upc.dcache/mem_addr[7]
+ top_cw.upc.dcache/mem_addr[8] top_cw.upc.dcache/mem_addr[9] top_cw.upc.dcache/mem_cache_enable
+ top_cw.upc.dcache/mem_exception top_cw.upc.core/o_mem_data[0] top_cw.upc.core/o_mem_data[10]
+ top_cw.upc.core/o_mem_data[11] top_cw.upc.core/o_mem_data[12] top_cw.upc.core/o_mem_data[13]
+ top_cw.upc.core/o_mem_data[14] top_cw.upc.core/o_mem_data[15] top_cw.upc.core/o_mem_data[1]
+ top_cw.upc.core/o_mem_data[2] top_cw.upc.core/o_mem_data[3] top_cw.upc.core/o_mem_data[4]
+ top_cw.upc.core/o_mem_data[5] top_cw.upc.core/o_mem_data[6] top_cw.upc.core/o_mem_data[7]
+ top_cw.upc.core/o_mem_data[8] top_cw.upc.core/o_mem_data[9] top_cw.upc.core/i_mem_data[0]
+ top_cw.upc.core/i_mem_data[10] top_cw.upc.core/i_mem_data[11] top_cw.upc.core/i_mem_data[12]
+ top_cw.upc.core/i_mem_data[13] top_cw.upc.core/i_mem_data[14] top_cw.upc.core/i_mem_data[15]
+ top_cw.upc.core/i_mem_data[1] top_cw.upc.core/i_mem_data[2] top_cw.upc.core/i_mem_data[3]
+ top_cw.upc.core/i_mem_data[4] top_cw.upc.core/i_mem_data[5] top_cw.upc.core/i_mem_data[6]
+ top_cw.upc.core/i_mem_data[7] top_cw.upc.core/i_mem_data[8] top_cw.upc.core/i_mem_data[9]
+ top_cw.upc.dcache/mem_req top_cw.upc.dcache/mem_sel[0] top_cw.upc.dcache/mem_sel[1]
+ top_cw.upc.dcache/mem_we vccd1 vssd1 top_cw.upc.dcache/wb_4_burst top_cw.upc.dcache/wb_ack
+ top_cw.upc.dcache/wb_adr[0] top_cw.upc.dcache/wb_adr[10] top_cw.upc.dcache/wb_adr[11]
+ top_cw.upc.dcache/wb_adr[12] top_cw.upc.dcache/wb_adr[13] top_cw.upc.dcache/wb_adr[14]
+ top_cw.upc.dcache/wb_adr[15] top_cw.upc.dcache/wb_adr[16] top_cw.upc.dcache/wb_adr[17]
+ top_cw.upc.dcache/wb_adr[18] top_cw.upc.dcache/wb_adr[19] top_cw.upc.dcache/wb_adr[1]
+ top_cw.upc.dcache/wb_adr[20] top_cw.upc.dcache/wb_adr[21] top_cw.upc.dcache/wb_adr[22]
+ top_cw.upc.dcache/wb_adr[23] top_cw.upc.dcache/wb_adr[2] top_cw.upc.dcache/wb_adr[3]
+ top_cw.upc.dcache/wb_adr[4] top_cw.upc.dcache/wb_adr[5] top_cw.upc.dcache/wb_adr[6]
+ top_cw.upc.dcache/wb_adr[7] top_cw.upc.dcache/wb_adr[8] top_cw.upc.dcache/wb_adr[9]
+ top_cw.upc.dcache/wb_cyc top_cw.upc.dcache/wb_err top_cw.upc.icache/wb_i_dat[0]
+ top_cw.upc.icache/wb_i_dat[10] top_cw.upc.icache/wb_i_dat[11] top_cw.upc.icache/wb_i_dat[12]
+ top_cw.upc.icache/wb_i_dat[13] top_cw.upc.icache/wb_i_dat[14] top_cw.upc.icache/wb_i_dat[15]
+ top_cw.upc.icache/wb_i_dat[1] top_cw.upc.icache/wb_i_dat[2] top_cw.upc.icache/wb_i_dat[3]
+ top_cw.upc.icache/wb_i_dat[4] top_cw.upc.icache/wb_i_dat[5] top_cw.upc.icache/wb_i_dat[6]
+ top_cw.upc.icache/wb_i_dat[7] top_cw.upc.icache/wb_i_dat[8] top_cw.upc.icache/wb_i_dat[9]
+ top_cw.upc.dcache/wb_o_dat[0] top_cw.upc.dcache/wb_o_dat[10] top_cw.upc.dcache/wb_o_dat[11]
+ top_cw.upc.dcache/wb_o_dat[12] top_cw.upc.dcache/wb_o_dat[13] top_cw.upc.dcache/wb_o_dat[14]
+ top_cw.upc.dcache/wb_o_dat[15] top_cw.upc.dcache/wb_o_dat[1] top_cw.upc.dcache/wb_o_dat[2]
+ top_cw.upc.dcache/wb_o_dat[3] top_cw.upc.dcache/wb_o_dat[4] top_cw.upc.dcache/wb_o_dat[5]
+ top_cw.upc.dcache/wb_o_dat[6] top_cw.upc.dcache/wb_o_dat[7] top_cw.upc.dcache/wb_o_dat[8]
+ top_cw.upc.dcache/wb_o_dat[9] top_cw.upc.dcache/wb_sel[0] top_cw.upc.dcache/wb_sel[1]
+ top_cw.upc.dcache/wb_stb top_cw.upc.dcache/wb_we dcache
Xtop_cw.clk_div la_data_in[104] top_cw.clk_div/div[0] top_cw.clk_div/div[1] top_cw.clk_div/div[2]
+ top_cw.clk_div/div[3] top_cw.clk_div/div_we user_clock2 top_cw.clk_div/i_rst top_cw.clk_div/o_clk
+ vccd1 vssd1 clk_div
Xtop_cw.upc.upper_core_logic top_cw.upc.core/o_c_data_page top_cw.upc.core/o_c_instr_page
+ top_cw.upc.dcache/mem_cache_enable top_cw.upc.core/o_mem_addr[0] top_cw.upc.core/o_mem_addr[10]
+ top_cw.upc.core/o_mem_addr[11] top_cw.upc.core/o_mem_addr[12] top_cw.upc.core/o_mem_addr[13]
+ top_cw.upc.core/o_mem_addr[14] top_cw.upc.core/o_mem_addr[15] top_cw.upc.core/o_mem_addr[1]
+ top_cw.upc.core/o_mem_addr[2] top_cw.upc.core/o_mem_addr[3] top_cw.upc.core/o_mem_addr[4]
+ top_cw.upc.core/o_mem_addr[5] top_cw.upc.core/o_mem_addr[6] top_cw.upc.core/o_mem_addr[7]
+ top_cw.upc.core/o_mem_addr[8] top_cw.upc.core/o_mem_addr[9] top_cw.upc.dcache/mem_addr[0]
+ top_cw.upc.dcache/mem_addr[10] top_cw.upc.dcache/mem_addr[11] top_cw.upc.dcache/mem_addr[12]
+ top_cw.upc.dcache/mem_addr[13] top_cw.upc.dcache/mem_addr[14] top_cw.upc.dcache/mem_addr[15]
+ top_cw.upc.dcache/mem_addr[16] top_cw.upc.dcache/mem_addr[17] top_cw.upc.dcache/mem_addr[18]
+ top_cw.upc.dcache/mem_addr[19] top_cw.upc.dcache/mem_addr[1] top_cw.upc.dcache/mem_addr[20]
+ top_cw.upc.dcache/mem_addr[21] top_cw.upc.dcache/mem_addr[22] top_cw.upc.dcache/mem_addr[23]
+ top_cw.upc.dcache/mem_addr[2] top_cw.upc.dcache/mem_addr[3] top_cw.upc.dcache/mem_addr[4]
+ top_cw.upc.dcache/mem_addr[5] top_cw.upc.dcache/mem_addr[6] top_cw.upc.dcache/mem_addr[7]
+ top_cw.upc.dcache/mem_addr[8] top_cw.upc.dcache/mem_addr[9] top_cw.upc.icache/wb_adr[0]
+ top_cw.upc.icache/wb_adr[10] top_cw.upc.icache/wb_adr[11] top_cw.upc.icache/wb_adr[12]
+ top_cw.upc.icache/wb_adr[13] top_cw.upc.icache/wb_adr[14] top_cw.upc.icache/wb_adr[15]
+ top_cw.upc.icache/wb_adr[1] top_cw.upc.icache/wb_adr[2] top_cw.upc.icache/wb_adr[3]
+ top_cw.upc.icache/wb_adr[4] top_cw.upc.icache/wb_adr[5] top_cw.upc.icache/wb_adr[6]
+ top_cw.upc.icache/wb_adr[7] top_cw.upc.icache/wb_adr[8] top_cw.upc.icache/wb_adr[9]
+ top_cw.upc.wb_arbiter/wb1_adr[0] top_cw.upc.wb_arbiter/wb1_adr[10] top_cw.upc.wb_arbiter/wb1_adr[11]
+ top_cw.upc.wb_arbiter/wb1_adr[12] top_cw.upc.wb_arbiter/wb1_adr[13] top_cw.upc.wb_arbiter/wb1_adr[14]
+ top_cw.upc.wb_arbiter/wb1_adr[15] top_cw.upc.wb_arbiter/wb1_adr[16] top_cw.upc.wb_arbiter/wb1_adr[17]
+ top_cw.upc.wb_arbiter/wb1_adr[18] top_cw.upc.wb_arbiter/wb1_adr[19] top_cw.upc.wb_arbiter/wb1_adr[1]
+ top_cw.upc.wb_arbiter/wb1_adr[20] top_cw.upc.wb_arbiter/wb1_adr[21] top_cw.upc.wb_arbiter/wb1_adr[22]
+ top_cw.upc.wb_arbiter/wb1_adr[23] top_cw.upc.wb_arbiter/wb1_adr[2] top_cw.upc.wb_arbiter/wb1_adr[3]
+ top_cw.upc.wb_arbiter/wb1_adr[4] top_cw.upc.wb_arbiter/wb1_adr[5] top_cw.upc.wb_arbiter/wb1_adr[6]
+ top_cw.upc.wb_arbiter/wb1_adr[7] top_cw.upc.wb_arbiter/wb1_adr[8] top_cw.upc.wb_arbiter/wb1_adr[9]
+ top_cw.upc.wb_arbiter/wb1_o_dat[0] top_cw.upc.wb_arbiter/wb1_o_dat[10] top_cw.upc.wb_arbiter/wb1_o_dat[11]
+ top_cw.upc.wb_arbiter/wb1_o_dat[12] top_cw.upc.wb_arbiter/wb1_o_dat[13] top_cw.upc.wb_arbiter/wb1_o_dat[14]
+ top_cw.upc.wb_arbiter/wb1_o_dat[15] top_cw.upc.wb_arbiter/wb1_o_dat[1] top_cw.upc.wb_arbiter/wb1_o_dat[2]
+ top_cw.upc.wb_arbiter/wb1_o_dat[3] top_cw.upc.wb_arbiter/wb1_o_dat[4] top_cw.upc.wb_arbiter/wb1_o_dat[5]
+ top_cw.upc.wb_arbiter/wb1_o_dat[6] top_cw.upc.wb_arbiter/wb1_o_dat[7] top_cw.upc.wb_arbiter/wb1_o_dat[8]
+ top_cw.upc.wb_arbiter/wb1_o_dat[9] user_clock2 top_cw.clk_div/i_rst top_cw.upc.core/sr_bus_addr[0]
+ top_cw.upc.core/sr_bus_addr[10] top_cw.upc.core/sr_bus_addr[11] top_cw.upc.core/sr_bus_addr[12]
+ top_cw.upc.core/sr_bus_addr[13] top_cw.upc.core/sr_bus_addr[14] top_cw.upc.core/sr_bus_addr[15]
+ top_cw.upc.core/sr_bus_addr[1] top_cw.upc.core/sr_bus_addr[2] top_cw.upc.core/sr_bus_addr[3]
+ top_cw.upc.core/sr_bus_addr[4] top_cw.upc.core/sr_bus_addr[5] top_cw.upc.core/sr_bus_addr[6]
+ top_cw.upc.core/sr_bus_addr[7] top_cw.upc.core/sr_bus_addr[8] top_cw.upc.core/sr_bus_addr[9]
+ top_cw.upc.core/sr_bus_data_o[0] top_cw.upc.core/sr_bus_data_o[10] top_cw.upc.core/sr_bus_data_o[11]
+ top_cw.upc.core/sr_bus_data_o[12] top_cw.upc.core/sr_bus_data_o[13] top_cw.upc.core/sr_bus_data_o[14]
+ top_cw.upc.core/sr_bus_data_o[15] top_cw.upc.core/sr_bus_data_o[1] top_cw.upc.core/sr_bus_data_o[2]
+ top_cw.upc.core/sr_bus_data_o[3] top_cw.upc.core/sr_bus_data_o[4] top_cw.upc.core/sr_bus_data_o[5]
+ top_cw.upc.core/sr_bus_data_o[6] top_cw.upc.core/sr_bus_data_o[7] top_cw.upc.core/sr_bus_data_o[8]
+ top_cw.upc.core/sr_bus_data_o[9] top_cw.upc.core/sr_bus_we vccd1 vssd1 top_cw.upc.wb_arbiter/wb0_8_burst
+ top_cw.upc.wb_arbiter/wb1_4_burst top_cw.upc.wb_arbiter/wb1_8_burst upper_core_logic
Xuprj_w_const la_data_out[98] la_data_out[108] la_data_out[109] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[99] la_data_out[118] la_data_out[119] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[100] la_data_out[78] la_data_out[79]
+ la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[101] la_data_out[88]
+ la_data_out[89] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] user_irq[0] user_irq[1] user_irq[2] la_data_out[102] wbs_ack_o wbs_dat_o[0]
+ wbs_dat_o[1] wbs_dat_o[2] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7]
+ wbs_dat_o[8] la_data_out[103] wbs_dat_o[9] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12]
+ wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18]
+ la_data_out[104] wbs_dat_o[19] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23]
+ wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] la_data_out[105]
+ wbs_dat_o[29] wbs_dat_o[30] wbs_dat_o[31] la_data_out[106] la_data_out[107] top_cw.clk_div/o_clk
+ io_out[16] uprj_w_const/cw_dir uprj_w_const/cw_dir_o io_out[18] uprj_w_const/cw_dir_o
+ uprj_w_const/cw_req_i io_out[17] uprj_w_const/cw_rst_i io_out[21] io_in[23] wb_rst_i
+ io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[1]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[20] io_oeb[21] io_oeb[22] io_out[23]
+ io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[24] io_out[25] io_out[26]
+ io_out[27] io_out[28] io_out[29] io_out[30] io_out[31] io_out[32] io_out[19] io_out[20]
+ io_out[22] la_data_out[16] la_data_out[17] la_data_out[21] la_data_out[36] la_data_out[37]
+ la_data_out[62] la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75]
+ la_data_out[76] la_data_out[77] la_data_out[63] la_data_out[64] la_data_out[65]
+ la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[70]
+ la_data_out[71] la_data_out[95] la_data_out[96] la_data_out[97] uprj_w_const/la_datb_i[0]
+ uprj_w_const/la_datb_i[1] uprj_w_const/la_datb_i[2] la_data_out[36] la_data_out[37]
+ la_data_out[21] uprj_w_const/o_s_rst io_oeb[23] io_oeb[33] io_oeb[34] io_oeb[35]
+ io_oeb[36] io_oeb[37] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[30] io_oeb[31] io_oeb[32] la_data_in[105] vccd1 vssd1 uprj_w_const
Xtop_cw.top_cw_logic top_cw.wb_compressor/wb_4_burst top_cw.wb_compressor/wb_8_burst
+ top_cw.wb_compressor/wb_ack top_cw.wb_compressor/wb_adr[0] top_cw.wb_compressor/wb_adr[10]
+ top_cw.wb_compressor/wb_adr[11] top_cw.wb_compressor/wb_adr[12] top_cw.wb_compressor/wb_adr[13]
+ top_cw.wb_compressor/wb_adr[14] top_cw.wb_compressor/wb_adr[15] top_cw.wb_compressor/wb_adr[16]
+ top_cw.wb_compressor/wb_adr[17] top_cw.wb_compressor/wb_adr[18] top_cw.wb_compressor/wb_adr[19]
+ top_cw.wb_compressor/wb_adr[1] top_cw.wb_compressor/wb_adr[20] top_cw.wb_compressor/wb_adr[21]
+ top_cw.wb_compressor/wb_adr[22] top_cw.wb_compressor/wb_adr[23] top_cw.wb_compressor/wb_adr[2]
+ top_cw.wb_compressor/wb_adr[3] top_cw.wb_compressor/wb_adr[4] top_cw.wb_compressor/wb_adr[5]
+ top_cw.wb_compressor/wb_adr[6] top_cw.wb_compressor/wb_adr[7] top_cw.wb_compressor/wb_adr[8]
+ top_cw.wb_compressor/wb_adr[9] top_cw.wb_compressor/wb_cyc top_cw.wb_compressor/wb_err
+ top_cw.wb_compressor/wb_i_dat[0] top_cw.wb_compressor/wb_i_dat[10] top_cw.wb_compressor/wb_i_dat[11]
+ top_cw.wb_compressor/wb_i_dat[12] top_cw.wb_compressor/wb_i_dat[13] top_cw.wb_compressor/wb_i_dat[14]
+ top_cw.wb_compressor/wb_i_dat[15] top_cw.wb_compressor/wb_i_dat[1] top_cw.wb_compressor/wb_i_dat[2]
+ top_cw.wb_compressor/wb_i_dat[3] top_cw.wb_compressor/wb_i_dat[4] top_cw.wb_compressor/wb_i_dat[5]
+ top_cw.wb_compressor/wb_i_dat[6] top_cw.wb_compressor/wb_i_dat[7] top_cw.wb_compressor/wb_i_dat[8]
+ top_cw.wb_compressor/wb_i_dat[9] top_cw.wb_compressor/wb_o_dat[0] top_cw.wb_compressor/wb_o_dat[10]
+ top_cw.wb_compressor/wb_o_dat[11] top_cw.wb_compressor/wb_o_dat[12] top_cw.wb_compressor/wb_o_dat[13]
+ top_cw.wb_compressor/wb_o_dat[14] top_cw.wb_compressor/wb_o_dat[15] top_cw.wb_compressor/wb_o_dat[1]
+ top_cw.wb_compressor/wb_o_dat[2] top_cw.wb_compressor/wb_o_dat[3] top_cw.wb_compressor/wb_o_dat[4]
+ top_cw.wb_compressor/wb_o_dat[5] top_cw.wb_compressor/wb_o_dat[6] top_cw.wb_compressor/wb_o_dat[7]
+ top_cw.wb_compressor/wb_o_dat[8] top_cw.wb_compressor/wb_o_dat[9] top_cw.wb_compressor/wb_sel[0]
+ top_cw.wb_compressor/wb_sel[1] top_cw.wb_compressor/wb_stb top_cw.wb_compressor/wb_we
+ top_cw.wb_cross_clk/s_wb_4_burst top_cw.wb_cross_clk/s_wb_8_burst top_cw.wb_cross_clk/s_wb_adr[0]
+ top_cw.wb_cross_clk/s_wb_adr[10] top_cw.wb_cross_clk/s_wb_adr[11] top_cw.wb_cross_clk/s_wb_adr[12]
+ top_cw.wb_cross_clk/s_wb_adr[13] top_cw.wb_cross_clk/s_wb_adr[14] top_cw.wb_cross_clk/s_wb_adr[15]
+ top_cw.wb_cross_clk/s_wb_adr[16] top_cw.wb_cross_clk/s_wb_adr[17] top_cw.wb_cross_clk/s_wb_adr[18]
+ top_cw.wb_cross_clk/s_wb_adr[19] top_cw.wb_cross_clk/s_wb_adr[1] top_cw.wb_cross_clk/s_wb_adr[20]
+ top_cw.wb_cross_clk/s_wb_adr[21] top_cw.wb_cross_clk/s_wb_adr[22] top_cw.wb_cross_clk/s_wb_adr[23]
+ top_cw.wb_cross_clk/s_wb_adr[2] top_cw.wb_cross_clk/s_wb_adr[3] top_cw.wb_cross_clk/s_wb_adr[4]
+ top_cw.wb_cross_clk/s_wb_adr[5] top_cw.wb_cross_clk/s_wb_adr[6] top_cw.wb_cross_clk/s_wb_adr[7]
+ top_cw.wb_cross_clk/s_wb_adr[8] top_cw.wb_cross_clk/s_wb_adr[9] top_cw.wb_cross_clk/s_wb_cyc
+ top_cw.wb_cross_clk/s_wb_o_dat[0] top_cw.wb_cross_clk/s_wb_o_dat[10] top_cw.wb_cross_clk/s_wb_o_dat[11]
+ top_cw.wb_cross_clk/s_wb_o_dat[12] top_cw.wb_cross_clk/s_wb_o_dat[13] top_cw.wb_cross_clk/s_wb_o_dat[14]
+ top_cw.wb_cross_clk/s_wb_o_dat[15] top_cw.wb_cross_clk/s_wb_o_dat[1] top_cw.wb_cross_clk/s_wb_o_dat[2]
+ top_cw.wb_cross_clk/s_wb_o_dat[3] top_cw.wb_cross_clk/s_wb_o_dat[4] top_cw.wb_cross_clk/s_wb_o_dat[5]
+ top_cw.wb_cross_clk/s_wb_o_dat[6] top_cw.wb_cross_clk/s_wb_o_dat[7] top_cw.wb_cross_clk/s_wb_o_dat[8]
+ top_cw.wb_cross_clk/s_wb_o_dat[9] top_cw.wb_cross_clk/s_wb_sel[0] top_cw.wb_cross_clk/s_wb_sel[1]
+ top_cw.wb_cross_clk/s_wb_stb top_cw.wb_cross_clk/s_wb_we io_in[19] top_cw.clk_div/o_clk
+ io_in[20] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[1]
+ io_in[2] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] uprj_w_const/cw_rst_i
+ top_cw.top_cw_logic/cw_rst_z user_clock2 io_in[22] uprj_w_const/o_s_rst la_data_in[104]
+ top_cw.upc.core/i_irq la_data_in[94] la_data_in[78] la_data_in[88] la_data_in[89]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[79] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[98] top_cw.wb_compressor/cw_ack top_cw.wb_compressor/cw_err
+ top_cw.wb_compressor/cw_io_i[0] top_cw.wb_compressor/cw_io_i[10] top_cw.wb_compressor/cw_io_i[11]
+ top_cw.wb_compressor/cw_io_i[12] top_cw.wb_compressor/cw_io_i[13] top_cw.wb_compressor/cw_io_i[14]
+ top_cw.wb_compressor/cw_io_i[15] top_cw.wb_compressor/cw_io_i[1] top_cw.wb_compressor/cw_io_i[2]
+ top_cw.wb_compressor/cw_io_i[3] top_cw.wb_compressor/cw_io_i[4] top_cw.wb_compressor/cw_io_i[5]
+ top_cw.wb_compressor/cw_io_i[6] top_cw.wb_compressor/cw_io_i[7] top_cw.wb_compressor/cw_io_i[8]
+ top_cw.wb_compressor/cw_io_i[9] top_cw.clk_div/i_rst top_cw.wb_cross_clk/m_wb_4_burst
+ top_cw.wb_cross_clk/m_wb_8_burst top_cw.top_cw_logic/u_wb_ack top_cw.wb_cross_clk/m_wb_ack
+ top_cw.clk_div/div_we top_cw.top_cw_logic/u_wb_ack_mxed la_data_out[38] la_data_out[48]
+ la_data_out[49] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[39]
+ la_data_out[58] la_data_out[59] la_data_out[60] la_data_out[61] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] top_cw.wb_cross_clk/m_wb_cyc top_cw.top_cw_logic/u_wb_err
+ top_cw.wb_cross_clk/m_wb_err top_cw.upc.icache/wb_i_dat[0] top_cw.upc.icache/wb_i_dat[10]
+ top_cw.upc.icache/wb_i_dat[11] top_cw.upc.icache/wb_i_dat[12] top_cw.upc.icache/wb_i_dat[13]
+ top_cw.upc.icache/wb_i_dat[14] top_cw.upc.icache/wb_i_dat[15] top_cw.upc.icache/wb_i_dat[1]
+ top_cw.upc.icache/wb_i_dat[2] top_cw.upc.icache/wb_i_dat[3] top_cw.upc.icache/wb_i_dat[4]
+ top_cw.upc.icache/wb_i_dat[5] top_cw.upc.icache/wb_i_dat[6] top_cw.upc.icache/wb_i_dat[7]
+ top_cw.upc.icache/wb_i_dat[8] top_cw.upc.icache/wb_i_dat[9] top_cw.wb_cross_clk/m_wb_i_dat[0]
+ top_cw.wb_cross_clk/m_wb_i_dat[10] top_cw.wb_cross_clk/m_wb_i_dat[11] top_cw.wb_cross_clk/m_wb_i_dat[12]
+ top_cw.wb_cross_clk/m_wb_i_dat[13] top_cw.wb_cross_clk/m_wb_i_dat[14] top_cw.wb_cross_clk/m_wb_i_dat[15]
+ top_cw.wb_cross_clk/m_wb_i_dat[1] top_cw.wb_cross_clk/m_wb_i_dat[2] top_cw.wb_cross_clk/m_wb_i_dat[3]
+ top_cw.wb_cross_clk/m_wb_i_dat[4] top_cw.wb_cross_clk/m_wb_i_dat[5] top_cw.wb_cross_clk/m_wb_i_dat[6]
+ top_cw.wb_cross_clk/m_wb_i_dat[7] top_cw.wb_cross_clk/m_wb_i_dat[8] top_cw.wb_cross_clk/m_wb_i_dat[9]
+ top_cw.clk_div/div[0] top_cw.wb_cross_clk/m_wb_o_dat[10] top_cw.wb_cross_clk/m_wb_o_dat[11]
+ top_cw.wb_cross_clk/m_wb_o_dat[12] top_cw.wb_cross_clk/m_wb_o_dat[13] top_cw.wb_cross_clk/m_wb_o_dat[14]
+ top_cw.wb_cross_clk/m_wb_o_dat[15] top_cw.clk_div/div[1] top_cw.clk_div/div[2] top_cw.clk_div/div[3]
+ top_cw.wb_cross_clk/m_wb_o_dat[4] top_cw.wb_cross_clk/m_wb_o_dat[5] top_cw.wb_cross_clk/m_wb_o_dat[6]
+ top_cw.wb_cross_clk/m_wb_o_dat[7] top_cw.wb_cross_clk/m_wb_o_dat[8] top_cw.wb_cross_clk/m_wb_o_dat[9]
+ top_cw.wb_cross_clk/m_wb_sel[0] top_cw.wb_cross_clk/m_wb_sel[1] uprj_w_const/la_datb_i[0]
+ uprj_w_const/la_datb_i[1] vccd1 vssd1 top_cw_logic
Xtop_cw.upc.wb_arbiter user_clock2 top_cw.clk_div/i_rst top_cw.upc.dcache/wb_cyc top_cw.upc.icache/wb_cyc
+ top_cw.upc.wb_arbiter/o_sel_sig top_cw.wb_cross_clk/m_wb_cyc top_cw.wb_cross_clk/m_wb_4_burst
+ top_cw.wb_cross_clk/m_wb_8_burst top_cw.top_cw_logic/u_wb_ack la_data_out[38] la_data_out[48]
+ la_data_out[49] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[39]
+ la_data_out[58] la_data_out[59] la_data_out[60] la_data_out[61] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] top_cw.top_cw_logic/u_wb_err top_cw.clk_div/div[0]
+ top_cw.wb_cross_clk/m_wb_o_dat[10] top_cw.wb_cross_clk/m_wb_o_dat[11] top_cw.wb_cross_clk/m_wb_o_dat[12]
+ top_cw.wb_cross_clk/m_wb_o_dat[13] top_cw.wb_cross_clk/m_wb_o_dat[14] top_cw.wb_cross_clk/m_wb_o_dat[15]
+ top_cw.clk_div/div[1] top_cw.clk_div/div[2] top_cw.clk_div/div[3] top_cw.wb_cross_clk/m_wb_o_dat[4]
+ top_cw.wb_cross_clk/m_wb_o_dat[5] top_cw.wb_cross_clk/m_wb_o_dat[6] top_cw.wb_cross_clk/m_wb_o_dat[7]
+ top_cw.wb_cross_clk/m_wb_o_dat[8] top_cw.wb_cross_clk/m_wb_o_dat[9] top_cw.wb_cross_clk/m_wb_sel[0]
+ top_cw.wb_cross_clk/m_wb_sel[1] uprj_w_const/la_datb_i[0] uprj_w_const/la_datb_i[1]
+ vccd1 vssd1 top_cw.upc.dcache/wb_4_burst top_cw.upc.wb_arbiter/wb0_8_burst top_cw.upc.dcache/wb_ack
+ top_cw.upc.dcache/wb_adr[0] top_cw.upc.dcache/wb_adr[10] top_cw.upc.dcache/wb_adr[11]
+ top_cw.upc.dcache/wb_adr[12] top_cw.upc.dcache/wb_adr[13] top_cw.upc.dcache/wb_adr[14]
+ top_cw.upc.dcache/wb_adr[15] top_cw.upc.dcache/wb_adr[16] top_cw.upc.dcache/wb_adr[17]
+ top_cw.upc.dcache/wb_adr[18] top_cw.upc.dcache/wb_adr[19] top_cw.upc.dcache/wb_adr[1]
+ top_cw.upc.dcache/wb_adr[20] top_cw.upc.dcache/wb_adr[21] top_cw.upc.dcache/wb_adr[22]
+ top_cw.upc.dcache/wb_adr[23] top_cw.upc.dcache/wb_adr[2] top_cw.upc.dcache/wb_adr[3]
+ top_cw.upc.dcache/wb_adr[4] top_cw.upc.dcache/wb_adr[5] top_cw.upc.dcache/wb_adr[6]
+ top_cw.upc.dcache/wb_adr[7] top_cw.upc.dcache/wb_adr[8] top_cw.upc.dcache/wb_adr[9]
+ top_cw.upc.dcache/wb_err top_cw.upc.dcache/wb_o_dat[0] top_cw.upc.dcache/wb_o_dat[10]
+ top_cw.upc.dcache/wb_o_dat[11] top_cw.upc.dcache/wb_o_dat[12] top_cw.upc.dcache/wb_o_dat[13]
+ top_cw.upc.dcache/wb_o_dat[14] top_cw.upc.dcache/wb_o_dat[15] top_cw.upc.dcache/wb_o_dat[1]
+ top_cw.upc.dcache/wb_o_dat[2] top_cw.upc.dcache/wb_o_dat[3] top_cw.upc.dcache/wb_o_dat[4]
+ top_cw.upc.dcache/wb_o_dat[5] top_cw.upc.dcache/wb_o_dat[6] top_cw.upc.dcache/wb_o_dat[7]
+ top_cw.upc.dcache/wb_o_dat[8] top_cw.upc.dcache/wb_o_dat[9] top_cw.upc.dcache/wb_sel[0]
+ top_cw.upc.dcache/wb_sel[1] top_cw.upc.dcache/wb_stb top_cw.upc.dcache/wb_we top_cw.upc.wb_arbiter/wb1_4_burst
+ top_cw.upc.wb_arbiter/wb1_8_burst top_cw.upc.icache/wb_ack top_cw.upc.wb_arbiter/wb1_adr[0]
+ top_cw.upc.wb_arbiter/wb1_adr[10] top_cw.upc.wb_arbiter/wb1_adr[11] top_cw.upc.wb_arbiter/wb1_adr[12]
+ top_cw.upc.wb_arbiter/wb1_adr[13] top_cw.upc.wb_arbiter/wb1_adr[14] top_cw.upc.wb_arbiter/wb1_adr[15]
+ top_cw.upc.wb_arbiter/wb1_adr[16] top_cw.upc.wb_arbiter/wb1_adr[17] top_cw.upc.wb_arbiter/wb1_adr[18]
+ top_cw.upc.wb_arbiter/wb1_adr[19] top_cw.upc.wb_arbiter/wb1_adr[1] top_cw.upc.wb_arbiter/wb1_adr[20]
+ top_cw.upc.wb_arbiter/wb1_adr[21] top_cw.upc.wb_arbiter/wb1_adr[22] top_cw.upc.wb_arbiter/wb1_adr[23]
+ top_cw.upc.wb_arbiter/wb1_adr[2] top_cw.upc.wb_arbiter/wb1_adr[3] top_cw.upc.wb_arbiter/wb1_adr[4]
+ top_cw.upc.wb_arbiter/wb1_adr[5] top_cw.upc.wb_arbiter/wb1_adr[6] top_cw.upc.wb_arbiter/wb1_adr[7]
+ top_cw.upc.wb_arbiter/wb1_adr[8] top_cw.upc.wb_arbiter/wb1_adr[9] top_cw.upc.icache/wb_err
+ top_cw.upc.wb_arbiter/wb1_o_dat[0] top_cw.upc.wb_arbiter/wb1_o_dat[10] top_cw.upc.wb_arbiter/wb1_o_dat[11]
+ top_cw.upc.wb_arbiter/wb1_o_dat[12] top_cw.upc.wb_arbiter/wb1_o_dat[13] top_cw.upc.wb_arbiter/wb1_o_dat[14]
+ top_cw.upc.wb_arbiter/wb1_o_dat[15] top_cw.upc.wb_arbiter/wb1_o_dat[1] top_cw.upc.wb_arbiter/wb1_o_dat[2]
+ top_cw.upc.wb_arbiter/wb1_o_dat[3] top_cw.upc.wb_arbiter/wb1_o_dat[4] top_cw.upc.wb_arbiter/wb1_o_dat[5]
+ top_cw.upc.wb_arbiter/wb1_o_dat[6] top_cw.upc.wb_arbiter/wb1_o_dat[7] top_cw.upc.wb_arbiter/wb1_o_dat[8]
+ top_cw.upc.wb_arbiter/wb1_o_dat[9] top_cw.upc.icache/wb_sel[0] top_cw.upc.icache/wb_sel[1]
+ top_cw.upc.icache/wb_stb top_cw.upc.icache/wb_we wishbone_arbiter
Xtop_cw.upc.icache user_clock2 top_cw.clk_div/i_rst top_cw.upc.icache/mem_ack top_cw.upc.icache/mem_addr[0]
+ top_cw.upc.icache/mem_addr[10] top_cw.upc.icache/mem_addr[11] top_cw.upc.icache/mem_addr[12]
+ top_cw.upc.icache/mem_addr[13] top_cw.upc.icache/mem_addr[14] top_cw.upc.icache/mem_addr[15]
+ top_cw.upc.icache/mem_addr[1] top_cw.upc.icache/mem_addr[2] top_cw.upc.icache/mem_addr[3]
+ top_cw.upc.icache/mem_addr[4] top_cw.upc.icache/mem_addr[5] top_cw.upc.icache/mem_addr[6]
+ top_cw.upc.icache/mem_addr[7] top_cw.upc.icache/mem_addr[8] top_cw.upc.icache/mem_addr[9]
+ top_cw.upc.core/o_icache_flush top_cw.upc.icache/mem_data[0] top_cw.upc.icache/mem_data[10]
+ top_cw.upc.icache/mem_data[11] top_cw.upc.icache/mem_data[12] top_cw.upc.icache/mem_data[13]
+ top_cw.upc.icache/mem_data[14] top_cw.upc.icache/mem_data[15] top_cw.upc.icache/mem_data[16]
+ top_cw.upc.icache/mem_data[17] top_cw.upc.icache/mem_data[18] top_cw.upc.icache/mem_data[19]
+ top_cw.upc.icache/mem_data[1] top_cw.upc.icache/mem_data[20] top_cw.upc.icache/mem_data[21]
+ top_cw.upc.icache/mem_data[22] top_cw.upc.icache/mem_data[23] top_cw.upc.icache/mem_data[24]
+ top_cw.upc.icache/mem_data[25] top_cw.upc.icache/mem_data[26] top_cw.upc.icache/mem_data[27]
+ top_cw.upc.icache/mem_data[28] top_cw.upc.icache/mem_data[29] top_cw.upc.icache/mem_data[2]
+ top_cw.upc.icache/mem_data[30] top_cw.upc.icache/mem_data[31] top_cw.upc.icache/mem_data[3]
+ top_cw.upc.icache/mem_data[4] top_cw.upc.icache/mem_data[5] top_cw.upc.icache/mem_data[6]
+ top_cw.upc.icache/mem_data[7] top_cw.upc.icache/mem_data[8] top_cw.upc.icache/mem_data[9]
+ top_cw.upc.icache/mem_ppl_submit top_cw.upc.icache/mem_req vccd1 vssd1 top_cw.upc.icache/wb_ack
+ top_cw.upc.icache/wb_adr[0] top_cw.upc.icache/wb_adr[10] top_cw.upc.icache/wb_adr[11]
+ top_cw.upc.icache/wb_adr[12] top_cw.upc.icache/wb_adr[13] top_cw.upc.icache/wb_adr[14]
+ top_cw.upc.icache/wb_adr[15] top_cw.upc.icache/wb_adr[1] top_cw.upc.icache/wb_adr[2]
+ top_cw.upc.icache/wb_adr[3] top_cw.upc.icache/wb_adr[4] top_cw.upc.icache/wb_adr[5]
+ top_cw.upc.icache/wb_adr[6] top_cw.upc.icache/wb_adr[7] top_cw.upc.icache/wb_adr[8]
+ top_cw.upc.icache/wb_adr[9] top_cw.upc.icache/wb_cyc top_cw.upc.icache/wb_err top_cw.upc.icache/wb_i_dat[0]
+ top_cw.upc.icache/wb_i_dat[10] top_cw.upc.icache/wb_i_dat[11] top_cw.upc.icache/wb_i_dat[12]
+ top_cw.upc.icache/wb_i_dat[13] top_cw.upc.icache/wb_i_dat[14] top_cw.upc.icache/wb_i_dat[15]
+ top_cw.upc.icache/wb_i_dat[1] top_cw.upc.icache/wb_i_dat[2] top_cw.upc.icache/wb_i_dat[3]
+ top_cw.upc.icache/wb_i_dat[4] top_cw.upc.icache/wb_i_dat[5] top_cw.upc.icache/wb_i_dat[6]
+ top_cw.upc.icache/wb_i_dat[7] top_cw.upc.icache/wb_i_dat[8] top_cw.upc.icache/wb_i_dat[9]
+ top_cw.upc.icache/wb_sel[0] top_cw.upc.icache/wb_sel[1] top_cw.upc.icache/wb_stb
+ top_cw.upc.icache/wb_we icache
.ends

