magic
tech sky130B
magscale 1 2
timestamp 1662741341
<< nwell >>
rect 1066 161285 161498 161851
rect 1066 160197 161498 160763
rect 1066 159109 161498 159675
rect 1066 158021 161498 158587
rect 1066 156933 161498 157499
rect 1066 155845 161498 156411
rect 1066 154757 161498 155323
rect 1066 153669 161498 154235
rect 1066 152581 161498 153147
rect 1066 151493 161498 152059
rect 1066 150405 161498 150971
rect 1066 149317 161498 149883
rect 1066 148229 161498 148795
rect 1066 147141 161498 147707
rect 1066 146053 161498 146619
rect 1066 144965 161498 145531
rect 1066 143877 161498 144443
rect 1066 142789 161498 143355
rect 1066 141701 161498 142267
rect 1066 140613 161498 141179
rect 1066 139525 161498 140091
rect 1066 138437 161498 139003
rect 1066 137349 161498 137915
rect 1066 136261 161498 136827
rect 1066 135173 161498 135739
rect 1066 134085 161498 134651
rect 1066 132997 161498 133563
rect 1066 131909 161498 132475
rect 1066 130821 161498 131387
rect 1066 129733 161498 130299
rect 1066 128645 161498 129211
rect 1066 127557 161498 128123
rect 1066 126469 161498 127035
rect 1066 125381 161498 125947
rect 1066 124293 161498 124859
rect 1066 123205 161498 123771
rect 1066 122117 161498 122683
rect 1066 121029 161498 121595
rect 1066 119941 161498 120507
rect 1066 118853 161498 119419
rect 1066 117765 161498 118331
rect 1066 116677 161498 117243
rect 1066 115589 161498 116155
rect 1066 114501 161498 115067
rect 1066 113413 161498 113979
rect 1066 112325 161498 112891
rect 1066 111237 161498 111803
rect 1066 110149 161498 110715
rect 1066 109061 161498 109627
rect 1066 107973 161498 108539
rect 1066 106885 161498 107451
rect 1066 105797 161498 106363
rect 1066 104709 161498 105275
rect 1066 103621 161498 104187
rect 1066 102533 161498 103099
rect 1066 101445 161498 102011
rect 1066 100357 161498 100923
rect 1066 99269 161498 99835
rect 1066 98181 161498 98747
rect 1066 97093 161498 97659
rect 1066 96005 161498 96571
rect 1066 94917 161498 95483
rect 1066 93829 161498 94395
rect 1066 92741 161498 93307
rect 1066 91653 161498 92219
rect 1066 90565 161498 91131
rect 1066 89477 161498 90043
rect 1066 88389 161498 88955
rect 1066 87301 161498 87867
rect 1066 86213 161498 86779
rect 1066 85125 161498 85691
rect 1066 84037 161498 84603
rect 1066 82949 161498 83515
rect 1066 81861 161498 82427
rect 1066 80773 161498 81339
rect 1066 79685 161498 80251
rect 1066 78597 161498 79163
rect 1066 77509 161498 78075
rect 1066 76421 161498 76987
rect 1066 75333 161498 75899
rect 1066 74245 161498 74811
rect 1066 73157 161498 73723
rect 1066 72069 161498 72635
rect 1066 70981 161498 71547
rect 1066 69893 161498 70459
rect 1066 68805 161498 69371
rect 1066 67717 161498 68283
rect 1066 66629 161498 67195
rect 1066 65541 161498 66107
rect 1066 64453 161498 65019
rect 1066 63365 161498 63931
rect 1066 62277 161498 62843
rect 1066 61189 161498 61755
rect 1066 60101 161498 60667
rect 1066 59013 161498 59579
rect 1066 57925 161498 58491
rect 1066 56837 161498 57403
rect 1066 55749 161498 56315
rect 1066 54661 161498 55227
rect 1066 53573 161498 54139
rect 1066 52485 161498 53051
rect 1066 51397 161498 51963
rect 1066 50309 161498 50875
rect 1066 49221 161498 49787
rect 1066 48133 161498 48699
rect 1066 47045 161498 47611
rect 1066 45957 161498 46523
rect 1066 44869 161498 45435
rect 1066 43781 161498 44347
rect 1066 42693 161498 43259
rect 1066 41605 161498 42171
rect 1066 40517 161498 41083
rect 1066 39429 161498 39995
rect 1066 38341 161498 38907
rect 1066 37253 161498 37819
rect 1066 36165 161498 36731
rect 1066 35077 161498 35643
rect 1066 33989 161498 34555
rect 1066 32901 161498 33467
rect 1066 31813 161498 32379
rect 1066 30725 161498 31291
rect 1066 29637 161498 30203
rect 1066 28549 161498 29115
rect 1066 27461 161498 28027
rect 1066 26373 161498 26939
rect 1066 25285 161498 25851
rect 1066 24197 161498 24763
rect 1066 23109 161498 23675
rect 1066 22021 161498 22587
rect 1066 20933 161498 21499
rect 1066 19845 161498 20411
rect 1066 18757 161498 19323
rect 1066 17669 161498 18235
rect 1066 16581 161498 17147
rect 1066 15493 161498 16059
rect 1066 14405 161498 14971
rect 1066 13317 161498 13883
rect 1066 12229 161498 12795
rect 1066 11141 161498 11707
rect 1066 10053 161498 10619
rect 1066 8965 161498 9531
rect 1066 7877 161498 8443
rect 1066 6789 161498 7355
rect 1066 5701 161498 6267
rect 1066 4613 161498 5179
rect 1066 3525 161498 4091
rect 1066 2437 161498 3003
<< obsli1 >>
rect 1104 2159 161460 162129
<< obsm1 >>
rect 1104 1844 161460 162444
<< metal2 >>
rect 2042 163952 2098 164752
rect 3974 163952 4030 164752
rect 5906 163952 5962 164752
rect 7838 163952 7894 164752
rect 9770 163952 9826 164752
rect 11702 163952 11758 164752
rect 13634 163952 13690 164752
rect 15566 163952 15622 164752
rect 17498 163952 17554 164752
rect 19430 163952 19486 164752
rect 21362 163952 21418 164752
rect 23294 163952 23350 164752
rect 25226 163952 25282 164752
rect 27158 163952 27214 164752
rect 29090 163952 29146 164752
rect 31022 163952 31078 164752
rect 32954 163952 33010 164752
rect 34886 163952 34942 164752
rect 36818 163952 36874 164752
rect 38750 163952 38806 164752
rect 40682 163952 40738 164752
rect 42614 163952 42670 164752
rect 44546 163952 44602 164752
rect 46478 163952 46534 164752
rect 48410 163952 48466 164752
rect 50342 163952 50398 164752
rect 52274 163952 52330 164752
rect 54206 163952 54262 164752
rect 56138 163952 56194 164752
rect 58070 163952 58126 164752
rect 60002 163952 60058 164752
rect 61934 163952 61990 164752
rect 63866 163952 63922 164752
rect 65798 163952 65854 164752
rect 67730 163952 67786 164752
rect 69662 163952 69718 164752
rect 71594 163952 71650 164752
rect 73526 163952 73582 164752
rect 75458 163952 75514 164752
rect 77390 163952 77446 164752
rect 79322 163952 79378 164752
rect 81254 163952 81310 164752
rect 83186 163952 83242 164752
rect 85118 163952 85174 164752
rect 87050 163952 87106 164752
rect 88982 163952 89038 164752
rect 90914 163952 90970 164752
rect 92846 163952 92902 164752
rect 94778 163952 94834 164752
rect 96710 163952 96766 164752
rect 98642 163952 98698 164752
rect 100574 163952 100630 164752
rect 102506 163952 102562 164752
rect 104438 163952 104494 164752
rect 106370 163952 106426 164752
rect 108302 163952 108358 164752
rect 110234 163952 110290 164752
rect 112166 163952 112222 164752
rect 114098 163952 114154 164752
rect 116030 163952 116086 164752
rect 117962 163952 118018 164752
rect 119894 163952 119950 164752
rect 121826 163952 121882 164752
rect 123758 163952 123814 164752
rect 125690 163952 125746 164752
rect 127622 163952 127678 164752
rect 129554 163952 129610 164752
rect 131486 163952 131542 164752
rect 133418 163952 133474 164752
rect 135350 163952 135406 164752
rect 137282 163952 137338 164752
rect 139214 163952 139270 164752
rect 141146 163952 141202 164752
rect 143078 163952 143134 164752
rect 145010 163952 145066 164752
rect 146942 163952 146998 164752
rect 148874 163952 148930 164752
rect 150806 163952 150862 164752
rect 152738 163952 152794 164752
rect 154670 163952 154726 164752
rect 156602 163952 156658 164752
rect 158534 163952 158590 164752
rect 160466 163952 160522 164752
rect 1214 0 1270 800
rect 3054 0 3110 800
rect 4894 0 4950 800
rect 6734 0 6790 800
rect 8574 0 8630 800
rect 10414 0 10470 800
rect 12254 0 12310 800
rect 14094 0 14150 800
rect 15934 0 15990 800
rect 17774 0 17830 800
rect 19614 0 19670 800
rect 21454 0 21510 800
rect 23294 0 23350 800
rect 25134 0 25190 800
rect 26974 0 27030 800
rect 28814 0 28870 800
rect 30654 0 30710 800
rect 32494 0 32550 800
rect 34334 0 34390 800
rect 36174 0 36230 800
rect 38014 0 38070 800
rect 39854 0 39910 800
rect 41694 0 41750 800
rect 43534 0 43590 800
rect 45374 0 45430 800
rect 47214 0 47270 800
rect 49054 0 49110 800
rect 50894 0 50950 800
rect 52734 0 52790 800
rect 54574 0 54630 800
rect 56414 0 56470 800
rect 58254 0 58310 800
rect 60094 0 60150 800
rect 61934 0 61990 800
rect 63774 0 63830 800
rect 65614 0 65670 800
rect 67454 0 67510 800
rect 69294 0 69350 800
rect 71134 0 71190 800
rect 72974 0 73030 800
rect 74814 0 74870 800
rect 76654 0 76710 800
rect 78494 0 78550 800
rect 80334 0 80390 800
rect 82174 0 82230 800
rect 84014 0 84070 800
rect 85854 0 85910 800
rect 87694 0 87750 800
rect 89534 0 89590 800
rect 91374 0 91430 800
rect 93214 0 93270 800
rect 95054 0 95110 800
rect 96894 0 96950 800
rect 98734 0 98790 800
rect 100574 0 100630 800
rect 102414 0 102470 800
rect 104254 0 104310 800
rect 106094 0 106150 800
rect 107934 0 107990 800
rect 109774 0 109830 800
rect 111614 0 111670 800
rect 113454 0 113510 800
rect 115294 0 115350 800
rect 117134 0 117190 800
rect 118974 0 119030 800
rect 120814 0 120870 800
rect 122654 0 122710 800
rect 124494 0 124550 800
rect 126334 0 126390 800
rect 128174 0 128230 800
rect 130014 0 130070 800
rect 131854 0 131910 800
rect 133694 0 133750 800
rect 135534 0 135590 800
rect 137374 0 137430 800
rect 139214 0 139270 800
rect 141054 0 141110 800
rect 142894 0 142950 800
rect 144734 0 144790 800
rect 146574 0 146630 800
rect 148414 0 148470 800
rect 150254 0 150310 800
rect 152094 0 152150 800
rect 153934 0 153990 800
rect 155774 0 155830 800
rect 157614 0 157670 800
rect 159454 0 159510 800
rect 161294 0 161350 800
<< obsm2 >>
rect 1228 163896 1986 164098
rect 2154 163896 3918 164098
rect 4086 163896 5850 164098
rect 6018 163896 7782 164098
rect 7950 163896 9714 164098
rect 9882 163896 11646 164098
rect 11814 163896 13578 164098
rect 13746 163896 15510 164098
rect 15678 163896 17442 164098
rect 17610 163896 19374 164098
rect 19542 163896 21306 164098
rect 21474 163896 23238 164098
rect 23406 163896 25170 164098
rect 25338 163896 27102 164098
rect 27270 163896 29034 164098
rect 29202 163896 30966 164098
rect 31134 163896 32898 164098
rect 33066 163896 34830 164098
rect 34998 163896 36762 164098
rect 36930 163896 38694 164098
rect 38862 163896 40626 164098
rect 40794 163896 42558 164098
rect 42726 163896 44490 164098
rect 44658 163896 46422 164098
rect 46590 163896 48354 164098
rect 48522 163896 50286 164098
rect 50454 163896 52218 164098
rect 52386 163896 54150 164098
rect 54318 163896 56082 164098
rect 56250 163896 58014 164098
rect 58182 163896 59946 164098
rect 60114 163896 61878 164098
rect 62046 163896 63810 164098
rect 63978 163896 65742 164098
rect 65910 163896 67674 164098
rect 67842 163896 69606 164098
rect 69774 163896 71538 164098
rect 71706 163896 73470 164098
rect 73638 163896 75402 164098
rect 75570 163896 77334 164098
rect 77502 163896 79266 164098
rect 79434 163896 81198 164098
rect 81366 163896 83130 164098
rect 83298 163896 85062 164098
rect 85230 163896 86994 164098
rect 87162 163896 88926 164098
rect 89094 163896 90858 164098
rect 91026 163896 92790 164098
rect 92958 163896 94722 164098
rect 94890 163896 96654 164098
rect 96822 163896 98586 164098
rect 98754 163896 100518 164098
rect 100686 163896 102450 164098
rect 102618 163896 104382 164098
rect 104550 163896 106314 164098
rect 106482 163896 108246 164098
rect 108414 163896 110178 164098
rect 110346 163896 112110 164098
rect 112278 163896 114042 164098
rect 114210 163896 115974 164098
rect 116142 163896 117906 164098
rect 118074 163896 119838 164098
rect 120006 163896 121770 164098
rect 121938 163896 123702 164098
rect 123870 163896 125634 164098
rect 125802 163896 127566 164098
rect 127734 163896 129498 164098
rect 129666 163896 131430 164098
rect 131598 163896 133362 164098
rect 133530 163896 135294 164098
rect 135462 163896 137226 164098
rect 137394 163896 139158 164098
rect 139326 163896 141090 164098
rect 141258 163896 143022 164098
rect 143190 163896 144954 164098
rect 145122 163896 146886 164098
rect 147054 163896 148818 164098
rect 148986 163896 150750 164098
rect 150918 163896 152682 164098
rect 152850 163896 154614 164098
rect 154782 163896 156546 164098
rect 156714 163896 158478 164098
rect 158646 163896 160410 164098
rect 160578 163896 161348 164098
rect 1228 856 161348 163896
rect 1326 734 2998 856
rect 3166 734 4838 856
rect 5006 734 6678 856
rect 6846 734 8518 856
rect 8686 734 10358 856
rect 10526 734 12198 856
rect 12366 734 14038 856
rect 14206 734 15878 856
rect 16046 734 17718 856
rect 17886 734 19558 856
rect 19726 734 21398 856
rect 21566 734 23238 856
rect 23406 734 25078 856
rect 25246 734 26918 856
rect 27086 734 28758 856
rect 28926 734 30598 856
rect 30766 734 32438 856
rect 32606 734 34278 856
rect 34446 734 36118 856
rect 36286 734 37958 856
rect 38126 734 39798 856
rect 39966 734 41638 856
rect 41806 734 43478 856
rect 43646 734 45318 856
rect 45486 734 47158 856
rect 47326 734 48998 856
rect 49166 734 50838 856
rect 51006 734 52678 856
rect 52846 734 54518 856
rect 54686 734 56358 856
rect 56526 734 58198 856
rect 58366 734 60038 856
rect 60206 734 61878 856
rect 62046 734 63718 856
rect 63886 734 65558 856
rect 65726 734 67398 856
rect 67566 734 69238 856
rect 69406 734 71078 856
rect 71246 734 72918 856
rect 73086 734 74758 856
rect 74926 734 76598 856
rect 76766 734 78438 856
rect 78606 734 80278 856
rect 80446 734 82118 856
rect 82286 734 83958 856
rect 84126 734 85798 856
rect 85966 734 87638 856
rect 87806 734 89478 856
rect 89646 734 91318 856
rect 91486 734 93158 856
rect 93326 734 94998 856
rect 95166 734 96838 856
rect 97006 734 98678 856
rect 98846 734 100518 856
rect 100686 734 102358 856
rect 102526 734 104198 856
rect 104366 734 106038 856
rect 106206 734 107878 856
rect 108046 734 109718 856
rect 109886 734 111558 856
rect 111726 734 113398 856
rect 113566 734 115238 856
rect 115406 734 117078 856
rect 117246 734 118918 856
rect 119086 734 120758 856
rect 120926 734 122598 856
rect 122766 734 124438 856
rect 124606 734 126278 856
rect 126446 734 128118 856
rect 128286 734 129958 856
rect 130126 734 131798 856
rect 131966 734 133638 856
rect 133806 734 135478 856
rect 135646 734 137318 856
rect 137486 734 139158 856
rect 139326 734 140998 856
rect 141166 734 142838 856
rect 143006 734 144678 856
rect 144846 734 146518 856
rect 146686 734 148358 856
rect 148526 734 150198 856
rect 150366 734 152038 856
rect 152206 734 153878 856
rect 154046 734 155718 856
rect 155886 734 157558 856
rect 157726 734 159398 856
rect 159566 734 161238 856
<< metal3 >>
rect 161808 123360 162608 123480
rect 161808 41080 162608 41200
<< obsm3 >>
rect 2221 123560 161808 162621
rect 2221 123280 161728 123560
rect 2221 41280 161808 123280
rect 2221 41000 161728 41280
rect 2221 1667 161808 41000
<< metal4 >>
rect 4208 2128 4528 162160
rect 19568 2128 19888 162160
rect 34928 2128 35248 162160
rect 50288 2128 50608 162160
rect 65648 2128 65968 162160
rect 81008 2128 81328 162160
rect 96368 2128 96688 162160
rect 111728 2128 112048 162160
rect 127088 2128 127408 162160
rect 142448 2128 142768 162160
rect 157808 2128 158128 162160
<< obsm4 >>
rect 10731 162240 157261 162621
rect 10731 2048 19488 162240
rect 19968 2048 34848 162240
rect 35328 2048 50208 162240
rect 50688 2048 65568 162240
rect 66048 2048 80928 162240
rect 81408 2048 96288 162240
rect 96768 2048 111648 162240
rect 112128 2048 127008 162240
rect 127488 2048 142368 162240
rect 142848 2048 157261 162240
rect 10731 1667 157261 2048
<< labels >>
rlabel metal2 s 1214 0 1270 800 6 i_addr[0]
port 1 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 i_addr[1]
port 2 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 i_addr[2]
port 3 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 i_addr[3]
port 4 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 i_addr[4]
port 5 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 i_addr[5]
port 6 nsew signal input
rlabel metal3 s 161808 41080 162608 41200 6 i_clk
port 7 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 i_data[0]
port 8 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 i_data[10]
port 9 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 i_data[11]
port 10 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 i_data[12]
port 11 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 i_data[13]
port 12 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 i_data[14]
port 13 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 i_data[15]
port 14 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 i_data[16]
port 15 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 i_data[17]
port 16 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 i_data[18]
port 17 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 i_data[19]
port 18 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 i_data[1]
port 19 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 i_data[20]
port 20 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 i_data[21]
port 21 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 i_data[22]
port 22 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 i_data[23]
port 23 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 i_data[24]
port 24 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 i_data[25]
port 25 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 i_data[26]
port 26 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 i_data[27]
port 27 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 i_data[28]
port 28 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 i_data[29]
port 29 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 i_data[2]
port 30 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 i_data[30]
port 31 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 i_data[31]
port 32 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 i_data[32]
port 33 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 i_data[33]
port 34 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 i_data[34]
port 35 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 i_data[35]
port 36 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 i_data[36]
port 37 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 i_data[37]
port 38 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 i_data[38]
port 39 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 i_data[39]
port 40 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 i_data[3]
port 41 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 i_data[40]
port 42 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 i_data[41]
port 43 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 i_data[42]
port 44 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 i_data[43]
port 45 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 i_data[44]
port 46 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 i_data[45]
port 47 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 i_data[46]
port 48 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 i_data[47]
port 49 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 i_data[48]
port 50 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 i_data[49]
port 51 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 i_data[4]
port 52 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 i_data[50]
port 53 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 i_data[51]
port 54 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 i_data[52]
port 55 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 i_data[53]
port 56 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 i_data[54]
port 57 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 i_data[55]
port 58 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 i_data[56]
port 59 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 i_data[57]
port 60 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 i_data[58]
port 61 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 i_data[59]
port 62 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 i_data[5]
port 63 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 i_data[60]
port 64 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 i_data[61]
port 65 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 i_data[62]
port 66 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 i_data[63]
port 67 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 i_data[64]
port 68 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 i_data[65]
port 69 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 i_data[66]
port 70 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 i_data[67]
port 71 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 i_data[68]
port 72 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 i_data[69]
port 73 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 i_data[6]
port 74 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 i_data[70]
port 75 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 i_data[71]
port 76 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 i_data[72]
port 77 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 i_data[73]
port 78 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 i_data[74]
port 79 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 i_data[75]
port 80 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 i_data[76]
port 81 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 i_data[77]
port 82 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 i_data[78]
port 83 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 i_data[79]
port 84 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 i_data[7]
port 85 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 i_data[80]
port 86 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 i_data[81]
port 87 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 i_data[8]
port 88 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 i_data[9]
port 89 nsew signal input
rlabel metal3 s 161808 123360 162608 123480 6 i_rst
port 90 nsew signal input
rlabel metal2 s 160466 163952 160522 164752 6 i_we
port 91 nsew signal input
rlabel metal2 s 2042 163952 2098 164752 6 o_data[0]
port 92 nsew signal output
rlabel metal2 s 21362 163952 21418 164752 6 o_data[10]
port 93 nsew signal output
rlabel metal2 s 23294 163952 23350 164752 6 o_data[11]
port 94 nsew signal output
rlabel metal2 s 25226 163952 25282 164752 6 o_data[12]
port 95 nsew signal output
rlabel metal2 s 27158 163952 27214 164752 6 o_data[13]
port 96 nsew signal output
rlabel metal2 s 29090 163952 29146 164752 6 o_data[14]
port 97 nsew signal output
rlabel metal2 s 31022 163952 31078 164752 6 o_data[15]
port 98 nsew signal output
rlabel metal2 s 32954 163952 33010 164752 6 o_data[16]
port 99 nsew signal output
rlabel metal2 s 34886 163952 34942 164752 6 o_data[17]
port 100 nsew signal output
rlabel metal2 s 36818 163952 36874 164752 6 o_data[18]
port 101 nsew signal output
rlabel metal2 s 38750 163952 38806 164752 6 o_data[19]
port 102 nsew signal output
rlabel metal2 s 3974 163952 4030 164752 6 o_data[1]
port 103 nsew signal output
rlabel metal2 s 40682 163952 40738 164752 6 o_data[20]
port 104 nsew signal output
rlabel metal2 s 42614 163952 42670 164752 6 o_data[21]
port 105 nsew signal output
rlabel metal2 s 44546 163952 44602 164752 6 o_data[22]
port 106 nsew signal output
rlabel metal2 s 46478 163952 46534 164752 6 o_data[23]
port 107 nsew signal output
rlabel metal2 s 48410 163952 48466 164752 6 o_data[24]
port 108 nsew signal output
rlabel metal2 s 50342 163952 50398 164752 6 o_data[25]
port 109 nsew signal output
rlabel metal2 s 52274 163952 52330 164752 6 o_data[26]
port 110 nsew signal output
rlabel metal2 s 54206 163952 54262 164752 6 o_data[27]
port 111 nsew signal output
rlabel metal2 s 56138 163952 56194 164752 6 o_data[28]
port 112 nsew signal output
rlabel metal2 s 58070 163952 58126 164752 6 o_data[29]
port 113 nsew signal output
rlabel metal2 s 5906 163952 5962 164752 6 o_data[2]
port 114 nsew signal output
rlabel metal2 s 60002 163952 60058 164752 6 o_data[30]
port 115 nsew signal output
rlabel metal2 s 61934 163952 61990 164752 6 o_data[31]
port 116 nsew signal output
rlabel metal2 s 63866 163952 63922 164752 6 o_data[32]
port 117 nsew signal output
rlabel metal2 s 65798 163952 65854 164752 6 o_data[33]
port 118 nsew signal output
rlabel metal2 s 67730 163952 67786 164752 6 o_data[34]
port 119 nsew signal output
rlabel metal2 s 69662 163952 69718 164752 6 o_data[35]
port 120 nsew signal output
rlabel metal2 s 71594 163952 71650 164752 6 o_data[36]
port 121 nsew signal output
rlabel metal2 s 73526 163952 73582 164752 6 o_data[37]
port 122 nsew signal output
rlabel metal2 s 75458 163952 75514 164752 6 o_data[38]
port 123 nsew signal output
rlabel metal2 s 77390 163952 77446 164752 6 o_data[39]
port 124 nsew signal output
rlabel metal2 s 7838 163952 7894 164752 6 o_data[3]
port 125 nsew signal output
rlabel metal2 s 79322 163952 79378 164752 6 o_data[40]
port 126 nsew signal output
rlabel metal2 s 81254 163952 81310 164752 6 o_data[41]
port 127 nsew signal output
rlabel metal2 s 83186 163952 83242 164752 6 o_data[42]
port 128 nsew signal output
rlabel metal2 s 85118 163952 85174 164752 6 o_data[43]
port 129 nsew signal output
rlabel metal2 s 87050 163952 87106 164752 6 o_data[44]
port 130 nsew signal output
rlabel metal2 s 88982 163952 89038 164752 6 o_data[45]
port 131 nsew signal output
rlabel metal2 s 90914 163952 90970 164752 6 o_data[46]
port 132 nsew signal output
rlabel metal2 s 92846 163952 92902 164752 6 o_data[47]
port 133 nsew signal output
rlabel metal2 s 94778 163952 94834 164752 6 o_data[48]
port 134 nsew signal output
rlabel metal2 s 96710 163952 96766 164752 6 o_data[49]
port 135 nsew signal output
rlabel metal2 s 9770 163952 9826 164752 6 o_data[4]
port 136 nsew signal output
rlabel metal2 s 98642 163952 98698 164752 6 o_data[50]
port 137 nsew signal output
rlabel metal2 s 100574 163952 100630 164752 6 o_data[51]
port 138 nsew signal output
rlabel metal2 s 102506 163952 102562 164752 6 o_data[52]
port 139 nsew signal output
rlabel metal2 s 104438 163952 104494 164752 6 o_data[53]
port 140 nsew signal output
rlabel metal2 s 106370 163952 106426 164752 6 o_data[54]
port 141 nsew signal output
rlabel metal2 s 108302 163952 108358 164752 6 o_data[55]
port 142 nsew signal output
rlabel metal2 s 110234 163952 110290 164752 6 o_data[56]
port 143 nsew signal output
rlabel metal2 s 112166 163952 112222 164752 6 o_data[57]
port 144 nsew signal output
rlabel metal2 s 114098 163952 114154 164752 6 o_data[58]
port 145 nsew signal output
rlabel metal2 s 116030 163952 116086 164752 6 o_data[59]
port 146 nsew signal output
rlabel metal2 s 11702 163952 11758 164752 6 o_data[5]
port 147 nsew signal output
rlabel metal2 s 117962 163952 118018 164752 6 o_data[60]
port 148 nsew signal output
rlabel metal2 s 119894 163952 119950 164752 6 o_data[61]
port 149 nsew signal output
rlabel metal2 s 121826 163952 121882 164752 6 o_data[62]
port 150 nsew signal output
rlabel metal2 s 123758 163952 123814 164752 6 o_data[63]
port 151 nsew signal output
rlabel metal2 s 125690 163952 125746 164752 6 o_data[64]
port 152 nsew signal output
rlabel metal2 s 127622 163952 127678 164752 6 o_data[65]
port 153 nsew signal output
rlabel metal2 s 129554 163952 129610 164752 6 o_data[66]
port 154 nsew signal output
rlabel metal2 s 131486 163952 131542 164752 6 o_data[67]
port 155 nsew signal output
rlabel metal2 s 133418 163952 133474 164752 6 o_data[68]
port 156 nsew signal output
rlabel metal2 s 135350 163952 135406 164752 6 o_data[69]
port 157 nsew signal output
rlabel metal2 s 13634 163952 13690 164752 6 o_data[6]
port 158 nsew signal output
rlabel metal2 s 137282 163952 137338 164752 6 o_data[70]
port 159 nsew signal output
rlabel metal2 s 139214 163952 139270 164752 6 o_data[71]
port 160 nsew signal output
rlabel metal2 s 141146 163952 141202 164752 6 o_data[72]
port 161 nsew signal output
rlabel metal2 s 143078 163952 143134 164752 6 o_data[73]
port 162 nsew signal output
rlabel metal2 s 145010 163952 145066 164752 6 o_data[74]
port 163 nsew signal output
rlabel metal2 s 146942 163952 146998 164752 6 o_data[75]
port 164 nsew signal output
rlabel metal2 s 148874 163952 148930 164752 6 o_data[76]
port 165 nsew signal output
rlabel metal2 s 150806 163952 150862 164752 6 o_data[77]
port 166 nsew signal output
rlabel metal2 s 152738 163952 152794 164752 6 o_data[78]
port 167 nsew signal output
rlabel metal2 s 154670 163952 154726 164752 6 o_data[79]
port 168 nsew signal output
rlabel metal2 s 15566 163952 15622 164752 6 o_data[7]
port 169 nsew signal output
rlabel metal2 s 156602 163952 156658 164752 6 o_data[80]
port 170 nsew signal output
rlabel metal2 s 158534 163952 158590 164752 6 o_data[81]
port 171 nsew signal output
rlabel metal2 s 17498 163952 17554 164752 6 o_data[8]
port 172 nsew signal output
rlabel metal2 s 19430 163952 19486 164752 6 o_data[9]
port 173 nsew signal output
rlabel metal4 s 4208 2128 4528 162160 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 162160 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 162160 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 162160 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 162160 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 162160 6 vccd1
port 174 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 162160 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 162160 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 162160 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 162160 6 vssd1
port 175 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 162160 6 vssd1
port 175 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 162608 164752
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 68129924
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/dcache_ram/runs/22_09_09_18_21/results/signoff/dcache_ram.magic.gds
string GDS_START 339778
<< end >>

