VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 800.000 ;
  PIN dbg_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END dbg_in[0]
  PIN dbg_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END dbg_in[1]
  PIN dbg_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END dbg_in[2]
  PIN dbg_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END dbg_in[3]
  PIN dbg_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END dbg_out[0]
  PIN dbg_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END dbg_out[10]
  PIN dbg_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END dbg_out[11]
  PIN dbg_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END dbg_out[12]
  PIN dbg_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END dbg_out[13]
  PIN dbg_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END dbg_out[14]
  PIN dbg_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END dbg_out[15]
  PIN dbg_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END dbg_out[16]
  PIN dbg_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END dbg_out[17]
  PIN dbg_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END dbg_out[18]
  PIN dbg_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END dbg_out[19]
  PIN dbg_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END dbg_out[1]
  PIN dbg_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END dbg_out[20]
  PIN dbg_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END dbg_out[21]
  PIN dbg_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END dbg_out[22]
  PIN dbg_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END dbg_out[23]
  PIN dbg_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END dbg_out[24]
  PIN dbg_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END dbg_out[25]
  PIN dbg_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END dbg_out[26]
  PIN dbg_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END dbg_out[27]
  PIN dbg_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END dbg_out[28]
  PIN dbg_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END dbg_out[29]
  PIN dbg_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END dbg_out[2]
  PIN dbg_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END dbg_out[30]
  PIN dbg_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END dbg_out[31]
  PIN dbg_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END dbg_out[32]
  PIN dbg_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END dbg_out[33]
  PIN dbg_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END dbg_out[34]
  PIN dbg_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END dbg_out[35]
  PIN dbg_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END dbg_out[3]
  PIN dbg_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END dbg_out[4]
  PIN dbg_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END dbg_out[5]
  PIN dbg_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END dbg_out[6]
  PIN dbg_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END dbg_out[7]
  PIN dbg_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END dbg_out[8]
  PIN dbg_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END dbg_out[9]
  PIN dbg_pc[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END dbg_pc[0]
  PIN dbg_pc[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END dbg_pc[10]
  PIN dbg_pc[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END dbg_pc[11]
  PIN dbg_pc[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END dbg_pc[12]
  PIN dbg_pc[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END dbg_pc[13]
  PIN dbg_pc[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END dbg_pc[14]
  PIN dbg_pc[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END dbg_pc[15]
  PIN dbg_pc[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END dbg_pc[1]
  PIN dbg_pc[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END dbg_pc[2]
  PIN dbg_pc[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END dbg_pc[3]
  PIN dbg_pc[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END dbg_pc[4]
  PIN dbg_pc[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END dbg_pc[5]
  PIN dbg_pc[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END dbg_pc[6]
  PIN dbg_pc[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END dbg_pc[7]
  PIN dbg_pc[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END dbg_pc[8]
  PIN dbg_pc[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END dbg_pc[9]
  PIN dbg_r0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END dbg_r0[0]
  PIN dbg_r0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END dbg_r0[10]
  PIN dbg_r0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END dbg_r0[11]
  PIN dbg_r0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END dbg_r0[12]
  PIN dbg_r0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END dbg_r0[13]
  PIN dbg_r0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END dbg_r0[14]
  PIN dbg_r0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END dbg_r0[15]
  PIN dbg_r0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END dbg_r0[1]
  PIN dbg_r0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END dbg_r0[2]
  PIN dbg_r0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END dbg_r0[3]
  PIN dbg_r0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END dbg_r0[4]
  PIN dbg_r0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END dbg_r0[5]
  PIN dbg_r0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END dbg_r0[6]
  PIN dbg_r0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END dbg_r0[7]
  PIN dbg_r0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END dbg_r0[8]
  PIN dbg_r0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END dbg_r0[9]
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.040 400.000 34.640 ;
    END
  END i_clk
  PIN i_core_int_sreg[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 703.160 400.000 703.760 ;
    END
  END i_core_int_sreg[0]
  PIN i_core_int_sreg[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 743.960 400.000 744.560 ;
    END
  END i_core_int_sreg[10]
  PIN i_core_int_sreg[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 748.040 400.000 748.640 ;
    END
  END i_core_int_sreg[11]
  PIN i_core_int_sreg[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 752.120 400.000 752.720 ;
    END
  END i_core_int_sreg[12]
  PIN i_core_int_sreg[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 756.200 400.000 756.800 ;
    END
  END i_core_int_sreg[13]
  PIN i_core_int_sreg[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 760.280 400.000 760.880 ;
    END
  END i_core_int_sreg[14]
  PIN i_core_int_sreg[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 764.360 400.000 764.960 ;
    END
  END i_core_int_sreg[15]
  PIN i_core_int_sreg[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 707.240 400.000 707.840 ;
    END
  END i_core_int_sreg[1]
  PIN i_core_int_sreg[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 711.320 400.000 711.920 ;
    END
  END i_core_int_sreg[2]
  PIN i_core_int_sreg[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 715.400 400.000 716.000 ;
    END
  END i_core_int_sreg[3]
  PIN i_core_int_sreg[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 719.480 400.000 720.080 ;
    END
  END i_core_int_sreg[4]
  PIN i_core_int_sreg[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 723.560 400.000 724.160 ;
    END
  END i_core_int_sreg[5]
  PIN i_core_int_sreg[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 727.640 400.000 728.240 ;
    END
  END i_core_int_sreg[6]
  PIN i_core_int_sreg[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 731.720 400.000 732.320 ;
    END
  END i_core_int_sreg[7]
  PIN i_core_int_sreg[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 735.800 400.000 736.400 ;
    END
  END i_core_int_sreg[8]
  PIN i_core_int_sreg[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 739.880 400.000 740.480 ;
    END
  END i_core_int_sreg[9]
  PIN i_disable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 695.000 400.000 695.600 ;
    END
  END i_disable
  PIN i_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 544.040 400.000 544.640 ;
    END
  END i_irq
  PIN i_mc_core_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 699.080 400.000 699.680 ;
    END
  END i_mc_core_int
  PIN i_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 287.000 400.000 287.600 ;
    END
  END i_mem_ack
  PIN i_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 140.120 400.000 140.720 ;
    END
  END i_mem_data[0]
  PIN i_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.720 400.000 222.320 ;
    END
  END i_mem_data[10]
  PIN i_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.880 400.000 230.480 ;
    END
  END i_mem_data[11]
  PIN i_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 238.040 400.000 238.640 ;
    END
  END i_mem_data[12]
  PIN i_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.200 400.000 246.800 ;
    END
  END i_mem_data[13]
  PIN i_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 254.360 400.000 254.960 ;
    END
  END i_mem_data[14]
  PIN i_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 262.520 400.000 263.120 ;
    END
  END i_mem_data[15]
  PIN i_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.280 400.000 148.880 ;
    END
  END i_mem_data[1]
  PIN i_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END i_mem_data[2]
  PIN i_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 164.600 400.000 165.200 ;
    END
  END i_mem_data[3]
  PIN i_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.760 400.000 173.360 ;
    END
  END i_mem_data[4]
  PIN i_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.920 400.000 181.520 ;
    END
  END i_mem_data[5]
  PIN i_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.080 400.000 189.680 ;
    END
  END i_mem_data[6]
  PIN i_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END i_mem_data[7]
  PIN i_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 205.400 400.000 206.000 ;
    END
  END i_mem_data[8]
  PIN i_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 213.560 400.000 214.160 ;
    END
  END i_mem_data[9]
  PIN i_mem_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 291.080 400.000 291.680 ;
    END
  END i_mem_exception
  PIN i_req_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 307.400 400.000 308.000 ;
    END
  END i_req_data[0]
  PIN i_req_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 389.000 400.000 389.600 ;
    END
  END i_req_data[10]
  PIN i_req_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.160 400.000 397.760 ;
    END
  END i_req_data[11]
  PIN i_req_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 405.320 400.000 405.920 ;
    END
  END i_req_data[12]
  PIN i_req_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 413.480 400.000 414.080 ;
    END
  END i_req_data[13]
  PIN i_req_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 421.640 400.000 422.240 ;
    END
  END i_req_data[14]
  PIN i_req_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 429.800 400.000 430.400 ;
    END
  END i_req_data[15]
  PIN i_req_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 437.960 400.000 438.560 ;
    END
  END i_req_data[16]
  PIN i_req_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 442.040 400.000 442.640 ;
    END
  END i_req_data[17]
  PIN i_req_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 446.120 400.000 446.720 ;
    END
  END i_req_data[18]
  PIN i_req_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 450.200 400.000 450.800 ;
    END
  END i_req_data[19]
  PIN i_req_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 315.560 400.000 316.160 ;
    END
  END i_req_data[1]
  PIN i_req_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 454.280 400.000 454.880 ;
    END
  END i_req_data[20]
  PIN i_req_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 458.360 400.000 458.960 ;
    END
  END i_req_data[21]
  PIN i_req_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 462.440 400.000 463.040 ;
    END
  END i_req_data[22]
  PIN i_req_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 466.520 400.000 467.120 ;
    END
  END i_req_data[23]
  PIN i_req_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 470.600 400.000 471.200 ;
    END
  END i_req_data[24]
  PIN i_req_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 474.680 400.000 475.280 ;
    END
  END i_req_data[25]
  PIN i_req_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 478.760 400.000 479.360 ;
    END
  END i_req_data[26]
  PIN i_req_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 482.840 400.000 483.440 ;
    END
  END i_req_data[27]
  PIN i_req_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 486.920 400.000 487.520 ;
    END
  END i_req_data[28]
  PIN i_req_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 491.000 400.000 491.600 ;
    END
  END i_req_data[29]
  PIN i_req_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.720 400.000 324.320 ;
    END
  END i_req_data[2]
  PIN i_req_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 495.080 400.000 495.680 ;
    END
  END i_req_data[30]
  PIN i_req_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 499.160 400.000 499.760 ;
    END
  END i_req_data[31]
  PIN i_req_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 331.880 400.000 332.480 ;
    END
  END i_req_data[3]
  PIN i_req_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 340.040 400.000 340.640 ;
    END
  END i_req_data[4]
  PIN i_req_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.200 400.000 348.800 ;
    END
  END i_req_data[5]
  PIN i_req_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 356.360 400.000 356.960 ;
    END
  END i_req_data[6]
  PIN i_req_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 364.520 400.000 365.120 ;
    END
  END i_req_data[7]
  PIN i_req_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.680 400.000 373.280 ;
    END
  END i_req_data[8]
  PIN i_req_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.840 400.000 381.440 ;
    END
  END i_req_data[9]
  PIN i_req_data_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.160 400.000 295.760 ;
    END
  END i_req_data_valid
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 38.120 400.000 38.720 ;
    END
  END i_rst
  PIN o_c_data_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 548.120 400.000 548.720 ;
    END
  END o_c_data_page
  PIN o_c_instr_long
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 503.240 400.000 503.840 ;
    END
  END o_c_instr_long
  PIN o_c_instr_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 552.200 400.000 552.800 ;
    END
  END o_c_instr_page
  PIN o_icache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 690.920 400.000 691.520 ;
    END
  END o_icache_flush
  PIN o_instr_long_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 511.400 400.000 512.000 ;
    END
  END o_instr_long_addr[0]
  PIN o_instr_long_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 515.480 400.000 516.080 ;
    END
  END o_instr_long_addr[1]
  PIN o_instr_long_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 519.560 400.000 520.160 ;
    END
  END o_instr_long_addr[2]
  PIN o_instr_long_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 523.640 400.000 524.240 ;
    END
  END o_instr_long_addr[3]
  PIN o_instr_long_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 527.720 400.000 528.320 ;
    END
  END o_instr_long_addr[4]
  PIN o_instr_long_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 531.800 400.000 532.400 ;
    END
  END o_instr_long_addr[5]
  PIN o_instr_long_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 535.880 400.000 536.480 ;
    END
  END o_instr_long_addr[6]
  PIN o_instr_long_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 539.960 400.000 540.560 ;
    END
  END o_instr_long_addr[7]
  PIN o_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.200 400.000 42.800 ;
    END
  END o_mem_addr[0]
  PIN o_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 115.640 400.000 116.240 ;
    END
  END o_mem_addr[10]
  PIN o_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.720 400.000 120.320 ;
    END
  END o_mem_addr[11]
  PIN o_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.800 400.000 124.400 ;
    END
  END o_mem_addr[12]
  PIN o_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 127.880 400.000 128.480 ;
    END
  END o_mem_addr[13]
  PIN o_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 131.960 400.000 132.560 ;
    END
  END o_mem_addr[14]
  PIN o_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 136.040 400.000 136.640 ;
    END
  END o_mem_addr[15]
  PIN o_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 50.360 400.000 50.960 ;
    END
  END o_mem_addr[1]
  PIN o_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 58.520 400.000 59.120 ;
    END
  END o_mem_addr[2]
  PIN o_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 66.680 400.000 67.280 ;
    END
  END o_mem_addr[3]
  PIN o_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.840 400.000 75.440 ;
    END
  END o_mem_addr[4]
  PIN o_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 83.000 400.000 83.600 ;
    END
  END o_mem_addr[5]
  PIN o_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 91.160 400.000 91.760 ;
    END
  END o_mem_addr[6]
  PIN o_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 99.320 400.000 99.920 ;
    END
  END o_mem_addr[7]
  PIN o_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 107.480 400.000 108.080 ;
    END
  END o_mem_addr[8]
  PIN o_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 111.560 400.000 112.160 ;
    END
  END o_mem_addr[9]
  PIN o_mem_addr_high[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 46.280 400.000 46.880 ;
    END
  END o_mem_addr_high[0]
  PIN o_mem_addr_high[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 54.440 400.000 55.040 ;
    END
  END o_mem_addr_high[1]
  PIN o_mem_addr_high[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 62.600 400.000 63.200 ;
    END
  END o_mem_addr_high[2]
  PIN o_mem_addr_high[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 70.760 400.000 71.360 ;
    END
  END o_mem_addr_high[3]
  PIN o_mem_addr_high[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.920 400.000 79.520 ;
    END
  END o_mem_addr_high[4]
  PIN o_mem_addr_high[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 87.080 400.000 87.680 ;
    END
  END o_mem_addr_high[5]
  PIN o_mem_addr_high[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.240 400.000 95.840 ;
    END
  END o_mem_addr_high[6]
  PIN o_mem_addr_high[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 103.400 400.000 104.000 ;
    END
  END o_mem_addr_high[7]
  PIN o_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 144.200 400.000 144.800 ;
    END
  END o_mem_data[0]
  PIN o_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.800 400.000 226.400 ;
    END
  END o_mem_data[10]
  PIN o_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 233.960 400.000 234.560 ;
    END
  END o_mem_data[11]
  PIN o_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 242.120 400.000 242.720 ;
    END
  END o_mem_data[12]
  PIN o_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.280 400.000 250.880 ;
    END
  END o_mem_data[13]
  PIN o_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 258.440 400.000 259.040 ;
    END
  END o_mem_data[14]
  PIN o_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 266.600 400.000 267.200 ;
    END
  END o_mem_data[15]
  PIN o_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 152.360 400.000 152.960 ;
    END
  END o_mem_data[1]
  PIN o_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 160.520 400.000 161.120 ;
    END
  END o_mem_data[2]
  PIN o_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 168.680 400.000 169.280 ;
    END
  END o_mem_data[3]
  PIN o_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.840 400.000 177.440 ;
    END
  END o_mem_data[4]
  PIN o_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 185.000 400.000 185.600 ;
    END
  END o_mem_data[5]
  PIN o_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.160 400.000 193.760 ;
    END
  END o_mem_data[6]
  PIN o_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 201.320 400.000 201.920 ;
    END
  END o_mem_data[7]
  PIN o_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 209.480 400.000 210.080 ;
    END
  END o_mem_data[8]
  PIN o_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 217.640 400.000 218.240 ;
    END
  END o_mem_data[9]
  PIN o_mem_long
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 507.320 400.000 507.920 ;
    END
  END o_mem_long
  PIN o_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 270.680 400.000 271.280 ;
    END
  END o_mem_req
  PIN o_mem_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.840 400.000 279.440 ;
    END
  END o_mem_sel[0]
  PIN o_mem_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.920 400.000 283.520 ;
    END
  END o_mem_sel[1]
  PIN o_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 274.760 400.000 275.360 ;
    END
  END o_mem_we
  PIN o_req_active
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 299.240 400.000 299.840 ;
    END
  END o_req_active
  PIN o_req_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 311.480 400.000 312.080 ;
    END
  END o_req_addr[0]
  PIN o_req_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.080 400.000 393.680 ;
    END
  END o_req_addr[10]
  PIN o_req_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 401.240 400.000 401.840 ;
    END
  END o_req_addr[11]
  PIN o_req_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 409.400 400.000 410.000 ;
    END
  END o_req_addr[12]
  PIN o_req_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 417.560 400.000 418.160 ;
    END
  END o_req_addr[13]
  PIN o_req_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 425.720 400.000 426.320 ;
    END
  END o_req_addr[14]
  PIN o_req_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 433.880 400.000 434.480 ;
    END
  END o_req_addr[15]
  PIN o_req_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 319.640 400.000 320.240 ;
    END
  END o_req_addr[1]
  PIN o_req_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 327.800 400.000 328.400 ;
    END
  END o_req_addr[2]
  PIN o_req_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 335.960 400.000 336.560 ;
    END
  END o_req_addr[3]
  PIN o_req_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.120 400.000 344.720 ;
    END
  END o_req_addr[4]
  PIN o_req_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.280 400.000 352.880 ;
    END
  END o_req_addr[5]
  PIN o_req_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 360.440 400.000 361.040 ;
    END
  END o_req_addr[6]
  PIN o_req_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 368.600 400.000 369.200 ;
    END
  END o_req_addr[7]
  PIN o_req_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.760 400.000 377.360 ;
    END
  END o_req_addr[8]
  PIN o_req_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 384.920 400.000 385.520 ;
    END
  END o_req_addr[9]
  PIN o_req_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 303.320 400.000 303.920 ;
    END
  END o_req_ppl_submit
  PIN sr_bus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 560.360 400.000 560.960 ;
    END
  END sr_bus_addr[0]
  PIN sr_bus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 641.960 400.000 642.560 ;
    END
  END sr_bus_addr[10]
  PIN sr_bus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 650.120 400.000 650.720 ;
    END
  END sr_bus_addr[11]
  PIN sr_bus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 658.280 400.000 658.880 ;
    END
  END sr_bus_addr[12]
  PIN sr_bus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 666.440 400.000 667.040 ;
    END
  END sr_bus_addr[13]
  PIN sr_bus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 674.600 400.000 675.200 ;
    END
  END sr_bus_addr[14]
  PIN sr_bus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 682.760 400.000 683.360 ;
    END
  END sr_bus_addr[15]
  PIN sr_bus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 568.520 400.000 569.120 ;
    END
  END sr_bus_addr[1]
  PIN sr_bus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 576.680 400.000 577.280 ;
    END
  END sr_bus_addr[2]
  PIN sr_bus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 584.840 400.000 585.440 ;
    END
  END sr_bus_addr[3]
  PIN sr_bus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 593.000 400.000 593.600 ;
    END
  END sr_bus_addr[4]
  PIN sr_bus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 601.160 400.000 601.760 ;
    END
  END sr_bus_addr[5]
  PIN sr_bus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 609.320 400.000 609.920 ;
    END
  END sr_bus_addr[6]
  PIN sr_bus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 617.480 400.000 618.080 ;
    END
  END sr_bus_addr[7]
  PIN sr_bus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 625.640 400.000 626.240 ;
    END
  END sr_bus_addr[8]
  PIN sr_bus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 633.800 400.000 634.400 ;
    END
  END sr_bus_addr[9]
  PIN sr_bus_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 564.440 400.000 565.040 ;
    END
  END sr_bus_data_o[0]
  PIN sr_bus_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 646.040 400.000 646.640 ;
    END
  END sr_bus_data_o[10]
  PIN sr_bus_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 654.200 400.000 654.800 ;
    END
  END sr_bus_data_o[11]
  PIN sr_bus_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 662.360 400.000 662.960 ;
    END
  END sr_bus_data_o[12]
  PIN sr_bus_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 670.520 400.000 671.120 ;
    END
  END sr_bus_data_o[13]
  PIN sr_bus_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 678.680 400.000 679.280 ;
    END
  END sr_bus_data_o[14]
  PIN sr_bus_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 686.840 400.000 687.440 ;
    END
  END sr_bus_data_o[15]
  PIN sr_bus_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 572.600 400.000 573.200 ;
    END
  END sr_bus_data_o[1]
  PIN sr_bus_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 580.760 400.000 581.360 ;
    END
  END sr_bus_data_o[2]
  PIN sr_bus_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 588.920 400.000 589.520 ;
    END
  END sr_bus_data_o[3]
  PIN sr_bus_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 597.080 400.000 597.680 ;
    END
  END sr_bus_data_o[4]
  PIN sr_bus_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 605.240 400.000 605.840 ;
    END
  END sr_bus_data_o[5]
  PIN sr_bus_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 613.400 400.000 614.000 ;
    END
  END sr_bus_data_o[6]
  PIN sr_bus_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 621.560 400.000 622.160 ;
    END
  END sr_bus_data_o[7]
  PIN sr_bus_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 629.720 400.000 630.320 ;
    END
  END sr_bus_data_o[8]
  PIN sr_bus_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 637.880 400.000 638.480 ;
    END
  END sr_bus_data_o[9]
  PIN sr_bus_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 556.280 400.000 556.880 ;
    END
  END sr_bus_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 788.885 ;
      LAYER met1 ;
        RECT 3.750 9.560 398.290 789.040 ;
      LAYER met2 ;
        RECT 3.780 4.280 398.260 788.985 ;
        RECT 4.330 4.000 9.010 4.280 ;
        RECT 9.850 4.000 14.530 4.280 ;
        RECT 15.370 4.000 20.050 4.280 ;
        RECT 20.890 4.000 25.570 4.280 ;
        RECT 26.410 4.000 31.090 4.280 ;
        RECT 31.930 4.000 36.610 4.280 ;
        RECT 37.450 4.000 42.130 4.280 ;
        RECT 42.970 4.000 47.650 4.280 ;
        RECT 48.490 4.000 53.170 4.280 ;
        RECT 54.010 4.000 58.690 4.280 ;
        RECT 59.530 4.000 64.210 4.280 ;
        RECT 65.050 4.000 69.730 4.280 ;
        RECT 70.570 4.000 75.250 4.280 ;
        RECT 76.090 4.000 80.770 4.280 ;
        RECT 81.610 4.000 86.290 4.280 ;
        RECT 87.130 4.000 91.810 4.280 ;
        RECT 92.650 4.000 97.330 4.280 ;
        RECT 98.170 4.000 102.850 4.280 ;
        RECT 103.690 4.000 108.370 4.280 ;
        RECT 109.210 4.000 113.890 4.280 ;
        RECT 114.730 4.000 119.410 4.280 ;
        RECT 120.250 4.000 124.930 4.280 ;
        RECT 125.770 4.000 130.450 4.280 ;
        RECT 131.290 4.000 135.970 4.280 ;
        RECT 136.810 4.000 141.490 4.280 ;
        RECT 142.330 4.000 147.010 4.280 ;
        RECT 147.850 4.000 152.530 4.280 ;
        RECT 153.370 4.000 158.050 4.280 ;
        RECT 158.890 4.000 163.570 4.280 ;
        RECT 164.410 4.000 169.090 4.280 ;
        RECT 169.930 4.000 174.610 4.280 ;
        RECT 175.450 4.000 180.130 4.280 ;
        RECT 180.970 4.000 185.650 4.280 ;
        RECT 186.490 4.000 191.170 4.280 ;
        RECT 192.010 4.000 196.690 4.280 ;
        RECT 197.530 4.000 202.210 4.280 ;
        RECT 203.050 4.000 207.730 4.280 ;
        RECT 208.570 4.000 213.250 4.280 ;
        RECT 214.090 4.000 218.770 4.280 ;
        RECT 219.610 4.000 224.290 4.280 ;
        RECT 225.130 4.000 229.810 4.280 ;
        RECT 230.650 4.000 235.330 4.280 ;
        RECT 236.170 4.000 240.850 4.280 ;
        RECT 241.690 4.000 246.370 4.280 ;
        RECT 247.210 4.000 251.890 4.280 ;
        RECT 252.730 4.000 257.410 4.280 ;
        RECT 258.250 4.000 262.930 4.280 ;
        RECT 263.770 4.000 268.450 4.280 ;
        RECT 269.290 4.000 273.970 4.280 ;
        RECT 274.810 4.000 279.490 4.280 ;
        RECT 280.330 4.000 285.010 4.280 ;
        RECT 285.850 4.000 290.530 4.280 ;
        RECT 291.370 4.000 296.050 4.280 ;
        RECT 296.890 4.000 301.570 4.280 ;
        RECT 302.410 4.000 307.090 4.280 ;
        RECT 307.930 4.000 312.610 4.280 ;
        RECT 313.450 4.000 318.130 4.280 ;
        RECT 318.970 4.000 323.650 4.280 ;
        RECT 324.490 4.000 329.170 4.280 ;
        RECT 330.010 4.000 334.690 4.280 ;
        RECT 335.530 4.000 340.210 4.280 ;
        RECT 341.050 4.000 345.730 4.280 ;
        RECT 346.570 4.000 351.250 4.280 ;
        RECT 352.090 4.000 356.770 4.280 ;
        RECT 357.610 4.000 362.290 4.280 ;
        RECT 363.130 4.000 367.810 4.280 ;
        RECT 368.650 4.000 373.330 4.280 ;
        RECT 374.170 4.000 378.850 4.280 ;
        RECT 379.690 4.000 384.370 4.280 ;
        RECT 385.210 4.000 389.890 4.280 ;
        RECT 390.730 4.000 395.410 4.280 ;
        RECT 396.250 4.000 398.260 4.280 ;
      LAYER met3 ;
        RECT 18.005 765.360 396.000 788.965 ;
        RECT 18.005 763.960 395.600 765.360 ;
        RECT 18.005 761.280 396.000 763.960 ;
        RECT 18.005 759.880 395.600 761.280 ;
        RECT 18.005 757.200 396.000 759.880 ;
        RECT 18.005 755.800 395.600 757.200 ;
        RECT 18.005 753.120 396.000 755.800 ;
        RECT 18.005 751.720 395.600 753.120 ;
        RECT 18.005 749.040 396.000 751.720 ;
        RECT 18.005 747.640 395.600 749.040 ;
        RECT 18.005 744.960 396.000 747.640 ;
        RECT 18.005 743.560 395.600 744.960 ;
        RECT 18.005 740.880 396.000 743.560 ;
        RECT 18.005 739.480 395.600 740.880 ;
        RECT 18.005 736.800 396.000 739.480 ;
        RECT 18.005 735.400 395.600 736.800 ;
        RECT 18.005 732.720 396.000 735.400 ;
        RECT 18.005 731.320 395.600 732.720 ;
        RECT 18.005 728.640 396.000 731.320 ;
        RECT 18.005 727.240 395.600 728.640 ;
        RECT 18.005 724.560 396.000 727.240 ;
        RECT 18.005 723.160 395.600 724.560 ;
        RECT 18.005 720.480 396.000 723.160 ;
        RECT 18.005 719.080 395.600 720.480 ;
        RECT 18.005 716.400 396.000 719.080 ;
        RECT 18.005 715.000 395.600 716.400 ;
        RECT 18.005 712.320 396.000 715.000 ;
        RECT 18.005 710.920 395.600 712.320 ;
        RECT 18.005 708.240 396.000 710.920 ;
        RECT 18.005 706.840 395.600 708.240 ;
        RECT 18.005 704.160 396.000 706.840 ;
        RECT 18.005 702.760 395.600 704.160 ;
        RECT 18.005 700.080 396.000 702.760 ;
        RECT 18.005 698.680 395.600 700.080 ;
        RECT 18.005 696.000 396.000 698.680 ;
        RECT 18.005 694.600 395.600 696.000 ;
        RECT 18.005 691.920 396.000 694.600 ;
        RECT 18.005 690.520 395.600 691.920 ;
        RECT 18.005 687.840 396.000 690.520 ;
        RECT 18.005 686.440 395.600 687.840 ;
        RECT 18.005 683.760 396.000 686.440 ;
        RECT 18.005 682.360 395.600 683.760 ;
        RECT 18.005 679.680 396.000 682.360 ;
        RECT 18.005 678.280 395.600 679.680 ;
        RECT 18.005 675.600 396.000 678.280 ;
        RECT 18.005 674.200 395.600 675.600 ;
        RECT 18.005 671.520 396.000 674.200 ;
        RECT 18.005 670.120 395.600 671.520 ;
        RECT 18.005 667.440 396.000 670.120 ;
        RECT 18.005 666.040 395.600 667.440 ;
        RECT 18.005 663.360 396.000 666.040 ;
        RECT 18.005 661.960 395.600 663.360 ;
        RECT 18.005 659.280 396.000 661.960 ;
        RECT 18.005 657.880 395.600 659.280 ;
        RECT 18.005 655.200 396.000 657.880 ;
        RECT 18.005 653.800 395.600 655.200 ;
        RECT 18.005 651.120 396.000 653.800 ;
        RECT 18.005 649.720 395.600 651.120 ;
        RECT 18.005 647.040 396.000 649.720 ;
        RECT 18.005 645.640 395.600 647.040 ;
        RECT 18.005 642.960 396.000 645.640 ;
        RECT 18.005 641.560 395.600 642.960 ;
        RECT 18.005 638.880 396.000 641.560 ;
        RECT 18.005 637.480 395.600 638.880 ;
        RECT 18.005 634.800 396.000 637.480 ;
        RECT 18.005 633.400 395.600 634.800 ;
        RECT 18.005 630.720 396.000 633.400 ;
        RECT 18.005 629.320 395.600 630.720 ;
        RECT 18.005 626.640 396.000 629.320 ;
        RECT 18.005 625.240 395.600 626.640 ;
        RECT 18.005 622.560 396.000 625.240 ;
        RECT 18.005 621.160 395.600 622.560 ;
        RECT 18.005 618.480 396.000 621.160 ;
        RECT 18.005 617.080 395.600 618.480 ;
        RECT 18.005 614.400 396.000 617.080 ;
        RECT 18.005 613.000 395.600 614.400 ;
        RECT 18.005 610.320 396.000 613.000 ;
        RECT 18.005 608.920 395.600 610.320 ;
        RECT 18.005 606.240 396.000 608.920 ;
        RECT 18.005 604.840 395.600 606.240 ;
        RECT 18.005 602.160 396.000 604.840 ;
        RECT 18.005 600.760 395.600 602.160 ;
        RECT 18.005 598.080 396.000 600.760 ;
        RECT 18.005 596.680 395.600 598.080 ;
        RECT 18.005 594.000 396.000 596.680 ;
        RECT 18.005 592.600 395.600 594.000 ;
        RECT 18.005 589.920 396.000 592.600 ;
        RECT 18.005 588.520 395.600 589.920 ;
        RECT 18.005 585.840 396.000 588.520 ;
        RECT 18.005 584.440 395.600 585.840 ;
        RECT 18.005 581.760 396.000 584.440 ;
        RECT 18.005 580.360 395.600 581.760 ;
        RECT 18.005 577.680 396.000 580.360 ;
        RECT 18.005 576.280 395.600 577.680 ;
        RECT 18.005 573.600 396.000 576.280 ;
        RECT 18.005 572.200 395.600 573.600 ;
        RECT 18.005 569.520 396.000 572.200 ;
        RECT 18.005 568.120 395.600 569.520 ;
        RECT 18.005 565.440 396.000 568.120 ;
        RECT 18.005 564.040 395.600 565.440 ;
        RECT 18.005 561.360 396.000 564.040 ;
        RECT 18.005 559.960 395.600 561.360 ;
        RECT 18.005 557.280 396.000 559.960 ;
        RECT 18.005 555.880 395.600 557.280 ;
        RECT 18.005 553.200 396.000 555.880 ;
        RECT 18.005 551.800 395.600 553.200 ;
        RECT 18.005 549.120 396.000 551.800 ;
        RECT 18.005 547.720 395.600 549.120 ;
        RECT 18.005 545.040 396.000 547.720 ;
        RECT 18.005 543.640 395.600 545.040 ;
        RECT 18.005 540.960 396.000 543.640 ;
        RECT 18.005 539.560 395.600 540.960 ;
        RECT 18.005 536.880 396.000 539.560 ;
        RECT 18.005 535.480 395.600 536.880 ;
        RECT 18.005 532.800 396.000 535.480 ;
        RECT 18.005 531.400 395.600 532.800 ;
        RECT 18.005 528.720 396.000 531.400 ;
        RECT 18.005 527.320 395.600 528.720 ;
        RECT 18.005 524.640 396.000 527.320 ;
        RECT 18.005 523.240 395.600 524.640 ;
        RECT 18.005 520.560 396.000 523.240 ;
        RECT 18.005 519.160 395.600 520.560 ;
        RECT 18.005 516.480 396.000 519.160 ;
        RECT 18.005 515.080 395.600 516.480 ;
        RECT 18.005 512.400 396.000 515.080 ;
        RECT 18.005 511.000 395.600 512.400 ;
        RECT 18.005 508.320 396.000 511.000 ;
        RECT 18.005 506.920 395.600 508.320 ;
        RECT 18.005 504.240 396.000 506.920 ;
        RECT 18.005 502.840 395.600 504.240 ;
        RECT 18.005 500.160 396.000 502.840 ;
        RECT 18.005 498.760 395.600 500.160 ;
        RECT 18.005 496.080 396.000 498.760 ;
        RECT 18.005 494.680 395.600 496.080 ;
        RECT 18.005 492.000 396.000 494.680 ;
        RECT 18.005 490.600 395.600 492.000 ;
        RECT 18.005 487.920 396.000 490.600 ;
        RECT 18.005 486.520 395.600 487.920 ;
        RECT 18.005 483.840 396.000 486.520 ;
        RECT 18.005 482.440 395.600 483.840 ;
        RECT 18.005 479.760 396.000 482.440 ;
        RECT 18.005 478.360 395.600 479.760 ;
        RECT 18.005 475.680 396.000 478.360 ;
        RECT 18.005 474.280 395.600 475.680 ;
        RECT 18.005 471.600 396.000 474.280 ;
        RECT 18.005 470.200 395.600 471.600 ;
        RECT 18.005 467.520 396.000 470.200 ;
        RECT 18.005 466.120 395.600 467.520 ;
        RECT 18.005 463.440 396.000 466.120 ;
        RECT 18.005 462.040 395.600 463.440 ;
        RECT 18.005 459.360 396.000 462.040 ;
        RECT 18.005 457.960 395.600 459.360 ;
        RECT 18.005 455.280 396.000 457.960 ;
        RECT 18.005 453.880 395.600 455.280 ;
        RECT 18.005 451.200 396.000 453.880 ;
        RECT 18.005 449.800 395.600 451.200 ;
        RECT 18.005 447.120 396.000 449.800 ;
        RECT 18.005 445.720 395.600 447.120 ;
        RECT 18.005 443.040 396.000 445.720 ;
        RECT 18.005 441.640 395.600 443.040 ;
        RECT 18.005 438.960 396.000 441.640 ;
        RECT 18.005 437.560 395.600 438.960 ;
        RECT 18.005 434.880 396.000 437.560 ;
        RECT 18.005 433.480 395.600 434.880 ;
        RECT 18.005 430.800 396.000 433.480 ;
        RECT 18.005 429.400 395.600 430.800 ;
        RECT 18.005 426.720 396.000 429.400 ;
        RECT 18.005 425.320 395.600 426.720 ;
        RECT 18.005 422.640 396.000 425.320 ;
        RECT 18.005 421.240 395.600 422.640 ;
        RECT 18.005 418.560 396.000 421.240 ;
        RECT 18.005 417.160 395.600 418.560 ;
        RECT 18.005 414.480 396.000 417.160 ;
        RECT 18.005 413.080 395.600 414.480 ;
        RECT 18.005 410.400 396.000 413.080 ;
        RECT 18.005 409.000 395.600 410.400 ;
        RECT 18.005 406.320 396.000 409.000 ;
        RECT 18.005 404.920 395.600 406.320 ;
        RECT 18.005 402.240 396.000 404.920 ;
        RECT 18.005 400.840 395.600 402.240 ;
        RECT 18.005 398.160 396.000 400.840 ;
        RECT 18.005 396.760 395.600 398.160 ;
        RECT 18.005 394.080 396.000 396.760 ;
        RECT 18.005 392.680 395.600 394.080 ;
        RECT 18.005 390.000 396.000 392.680 ;
        RECT 18.005 388.600 395.600 390.000 ;
        RECT 18.005 385.920 396.000 388.600 ;
        RECT 18.005 384.520 395.600 385.920 ;
        RECT 18.005 381.840 396.000 384.520 ;
        RECT 18.005 380.440 395.600 381.840 ;
        RECT 18.005 377.760 396.000 380.440 ;
        RECT 18.005 376.360 395.600 377.760 ;
        RECT 18.005 373.680 396.000 376.360 ;
        RECT 18.005 372.280 395.600 373.680 ;
        RECT 18.005 369.600 396.000 372.280 ;
        RECT 18.005 368.200 395.600 369.600 ;
        RECT 18.005 365.520 396.000 368.200 ;
        RECT 18.005 364.120 395.600 365.520 ;
        RECT 18.005 361.440 396.000 364.120 ;
        RECT 18.005 360.040 395.600 361.440 ;
        RECT 18.005 357.360 396.000 360.040 ;
        RECT 18.005 355.960 395.600 357.360 ;
        RECT 18.005 353.280 396.000 355.960 ;
        RECT 18.005 351.880 395.600 353.280 ;
        RECT 18.005 349.200 396.000 351.880 ;
        RECT 18.005 347.800 395.600 349.200 ;
        RECT 18.005 345.120 396.000 347.800 ;
        RECT 18.005 343.720 395.600 345.120 ;
        RECT 18.005 341.040 396.000 343.720 ;
        RECT 18.005 339.640 395.600 341.040 ;
        RECT 18.005 336.960 396.000 339.640 ;
        RECT 18.005 335.560 395.600 336.960 ;
        RECT 18.005 332.880 396.000 335.560 ;
        RECT 18.005 331.480 395.600 332.880 ;
        RECT 18.005 328.800 396.000 331.480 ;
        RECT 18.005 327.400 395.600 328.800 ;
        RECT 18.005 324.720 396.000 327.400 ;
        RECT 18.005 323.320 395.600 324.720 ;
        RECT 18.005 320.640 396.000 323.320 ;
        RECT 18.005 319.240 395.600 320.640 ;
        RECT 18.005 316.560 396.000 319.240 ;
        RECT 18.005 315.160 395.600 316.560 ;
        RECT 18.005 312.480 396.000 315.160 ;
        RECT 18.005 311.080 395.600 312.480 ;
        RECT 18.005 308.400 396.000 311.080 ;
        RECT 18.005 307.000 395.600 308.400 ;
        RECT 18.005 304.320 396.000 307.000 ;
        RECT 18.005 302.920 395.600 304.320 ;
        RECT 18.005 300.240 396.000 302.920 ;
        RECT 18.005 298.840 395.600 300.240 ;
        RECT 18.005 296.160 396.000 298.840 ;
        RECT 18.005 294.760 395.600 296.160 ;
        RECT 18.005 292.080 396.000 294.760 ;
        RECT 18.005 290.680 395.600 292.080 ;
        RECT 18.005 288.000 396.000 290.680 ;
        RECT 18.005 286.600 395.600 288.000 ;
        RECT 18.005 283.920 396.000 286.600 ;
        RECT 18.005 282.520 395.600 283.920 ;
        RECT 18.005 279.840 396.000 282.520 ;
        RECT 18.005 278.440 395.600 279.840 ;
        RECT 18.005 275.760 396.000 278.440 ;
        RECT 18.005 274.360 395.600 275.760 ;
        RECT 18.005 271.680 396.000 274.360 ;
        RECT 18.005 270.280 395.600 271.680 ;
        RECT 18.005 267.600 396.000 270.280 ;
        RECT 18.005 266.200 395.600 267.600 ;
        RECT 18.005 263.520 396.000 266.200 ;
        RECT 18.005 262.120 395.600 263.520 ;
        RECT 18.005 259.440 396.000 262.120 ;
        RECT 18.005 258.040 395.600 259.440 ;
        RECT 18.005 255.360 396.000 258.040 ;
        RECT 18.005 253.960 395.600 255.360 ;
        RECT 18.005 251.280 396.000 253.960 ;
        RECT 18.005 249.880 395.600 251.280 ;
        RECT 18.005 247.200 396.000 249.880 ;
        RECT 18.005 245.800 395.600 247.200 ;
        RECT 18.005 243.120 396.000 245.800 ;
        RECT 18.005 241.720 395.600 243.120 ;
        RECT 18.005 239.040 396.000 241.720 ;
        RECT 18.005 237.640 395.600 239.040 ;
        RECT 18.005 234.960 396.000 237.640 ;
        RECT 18.005 233.560 395.600 234.960 ;
        RECT 18.005 230.880 396.000 233.560 ;
        RECT 18.005 229.480 395.600 230.880 ;
        RECT 18.005 226.800 396.000 229.480 ;
        RECT 18.005 225.400 395.600 226.800 ;
        RECT 18.005 222.720 396.000 225.400 ;
        RECT 18.005 221.320 395.600 222.720 ;
        RECT 18.005 218.640 396.000 221.320 ;
        RECT 18.005 217.240 395.600 218.640 ;
        RECT 18.005 214.560 396.000 217.240 ;
        RECT 18.005 213.160 395.600 214.560 ;
        RECT 18.005 210.480 396.000 213.160 ;
        RECT 18.005 209.080 395.600 210.480 ;
        RECT 18.005 206.400 396.000 209.080 ;
        RECT 18.005 205.000 395.600 206.400 ;
        RECT 18.005 202.320 396.000 205.000 ;
        RECT 18.005 200.920 395.600 202.320 ;
        RECT 18.005 198.240 396.000 200.920 ;
        RECT 18.005 196.840 395.600 198.240 ;
        RECT 18.005 194.160 396.000 196.840 ;
        RECT 18.005 192.760 395.600 194.160 ;
        RECT 18.005 190.080 396.000 192.760 ;
        RECT 18.005 188.680 395.600 190.080 ;
        RECT 18.005 186.000 396.000 188.680 ;
        RECT 18.005 184.600 395.600 186.000 ;
        RECT 18.005 181.920 396.000 184.600 ;
        RECT 18.005 180.520 395.600 181.920 ;
        RECT 18.005 177.840 396.000 180.520 ;
        RECT 18.005 176.440 395.600 177.840 ;
        RECT 18.005 173.760 396.000 176.440 ;
        RECT 18.005 172.360 395.600 173.760 ;
        RECT 18.005 169.680 396.000 172.360 ;
        RECT 18.005 168.280 395.600 169.680 ;
        RECT 18.005 165.600 396.000 168.280 ;
        RECT 18.005 164.200 395.600 165.600 ;
        RECT 18.005 161.520 396.000 164.200 ;
        RECT 18.005 160.120 395.600 161.520 ;
        RECT 18.005 157.440 396.000 160.120 ;
        RECT 18.005 156.040 395.600 157.440 ;
        RECT 18.005 153.360 396.000 156.040 ;
        RECT 18.005 151.960 395.600 153.360 ;
        RECT 18.005 149.280 396.000 151.960 ;
        RECT 18.005 147.880 395.600 149.280 ;
        RECT 18.005 145.200 396.000 147.880 ;
        RECT 18.005 143.800 395.600 145.200 ;
        RECT 18.005 141.120 396.000 143.800 ;
        RECT 18.005 139.720 395.600 141.120 ;
        RECT 18.005 137.040 396.000 139.720 ;
        RECT 18.005 135.640 395.600 137.040 ;
        RECT 18.005 132.960 396.000 135.640 ;
        RECT 18.005 131.560 395.600 132.960 ;
        RECT 18.005 128.880 396.000 131.560 ;
        RECT 18.005 127.480 395.600 128.880 ;
        RECT 18.005 124.800 396.000 127.480 ;
        RECT 18.005 123.400 395.600 124.800 ;
        RECT 18.005 120.720 396.000 123.400 ;
        RECT 18.005 119.320 395.600 120.720 ;
        RECT 18.005 116.640 396.000 119.320 ;
        RECT 18.005 115.240 395.600 116.640 ;
        RECT 18.005 112.560 396.000 115.240 ;
        RECT 18.005 111.160 395.600 112.560 ;
        RECT 18.005 108.480 396.000 111.160 ;
        RECT 18.005 107.080 395.600 108.480 ;
        RECT 18.005 104.400 396.000 107.080 ;
        RECT 18.005 103.000 395.600 104.400 ;
        RECT 18.005 100.320 396.000 103.000 ;
        RECT 18.005 98.920 395.600 100.320 ;
        RECT 18.005 96.240 396.000 98.920 ;
        RECT 18.005 94.840 395.600 96.240 ;
        RECT 18.005 92.160 396.000 94.840 ;
        RECT 18.005 90.760 395.600 92.160 ;
        RECT 18.005 88.080 396.000 90.760 ;
        RECT 18.005 86.680 395.600 88.080 ;
        RECT 18.005 84.000 396.000 86.680 ;
        RECT 18.005 82.600 395.600 84.000 ;
        RECT 18.005 79.920 396.000 82.600 ;
        RECT 18.005 78.520 395.600 79.920 ;
        RECT 18.005 75.840 396.000 78.520 ;
        RECT 18.005 74.440 395.600 75.840 ;
        RECT 18.005 71.760 396.000 74.440 ;
        RECT 18.005 70.360 395.600 71.760 ;
        RECT 18.005 67.680 396.000 70.360 ;
        RECT 18.005 66.280 395.600 67.680 ;
        RECT 18.005 63.600 396.000 66.280 ;
        RECT 18.005 62.200 395.600 63.600 ;
        RECT 18.005 59.520 396.000 62.200 ;
        RECT 18.005 58.120 395.600 59.520 ;
        RECT 18.005 55.440 396.000 58.120 ;
        RECT 18.005 54.040 395.600 55.440 ;
        RECT 18.005 51.360 396.000 54.040 ;
        RECT 18.005 49.960 395.600 51.360 ;
        RECT 18.005 47.280 396.000 49.960 ;
        RECT 18.005 45.880 395.600 47.280 ;
        RECT 18.005 43.200 396.000 45.880 ;
        RECT 18.005 41.800 395.600 43.200 ;
        RECT 18.005 39.120 396.000 41.800 ;
        RECT 18.005 37.720 395.600 39.120 ;
        RECT 18.005 35.040 396.000 37.720 ;
        RECT 18.005 33.640 395.600 35.040 ;
        RECT 18.005 10.715 396.000 33.640 ;
      LAYER met4 ;
        RECT 181.535 18.535 251.040 772.985 ;
        RECT 253.440 18.535 327.840 772.985 ;
        RECT 330.240 18.535 386.105 772.985 ;
  END
END core
END LIBRARY

