magic
tech sky130B
magscale 1 2
timestamp 1663072423
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 235166 700612 235172 700664
rect 235224 700652 235230 700664
rect 253198 700652 253204 700664
rect 235224 700624 253204 700652
rect 235224 700612 235230 700624
rect 253198 700612 253204 700624
rect 253256 700612 253262 700664
rect 202782 700544 202788 700596
rect 202840 700584 202846 700596
rect 253290 700584 253296 700596
rect 202840 700556 253296 700584
rect 202840 700544 202846 700556
rect 253290 700544 253296 700556
rect 253348 700544 253354 700596
rect 348786 700544 348792 700596
rect 348844 700584 348850 700596
rect 409230 700584 409236 700596
rect 348844 700556 409236 700584
rect 348844 700544 348850 700556
rect 409230 700544 409236 700556
rect 409288 700544 409294 700596
rect 154114 700476 154120 700528
rect 154172 700516 154178 700528
rect 260098 700516 260104 700528
rect 154172 700488 260104 700516
rect 154172 700476 154178 700488
rect 260098 700476 260104 700488
rect 260156 700476 260162 700528
rect 404998 700476 405004 700528
rect 405056 700516 405062 700528
rect 559650 700516 559656 700528
rect 405056 700488 559656 700516
rect 405056 700476 405062 700488
rect 559650 700476 559656 700488
rect 559708 700476 559714 700528
rect 137830 700408 137836 700460
rect 137888 700448 137894 700460
rect 253382 700448 253388 700460
rect 137888 700420 253388 700448
rect 137888 700408 137894 700420
rect 253382 700408 253388 700420
rect 253440 700408 253446 700460
rect 317414 700408 317420 700460
rect 317472 700448 317478 700460
rect 543458 700448 543464 700460
rect 317472 700420 543464 700448
rect 317472 700408 317478 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 89162 700340 89168 700392
rect 89220 700380 89226 700392
rect 406470 700380 406476 700392
rect 89220 700352 406476 700380
rect 89220 700340 89226 700352
rect 406470 700340 406476 700352
rect 406528 700340 406534 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 472710 700312 472716 700324
rect 24360 700284 472716 700312
rect 24360 700272 24366 700284
rect 472710 700272 472716 700284
rect 472768 700272 472774 700324
rect 526438 699660 526444 699712
rect 526496 699700 526502 699712
rect 527174 699700 527180 699712
rect 526496 699672 527180 699700
rect 526496 699660 526502 699672
rect 527174 699660 527180 699672
rect 527232 699660 527238 699712
rect 397454 698912 397460 698964
rect 397512 698952 397518 698964
rect 458818 698952 458824 698964
rect 397512 698924 458824 698952
rect 397512 698912 397518 698924
rect 458818 698912 458824 698924
rect 458876 698912 458882 698964
rect 105446 697552 105452 697604
rect 105504 697592 105510 697604
rect 337378 697592 337384 697604
rect 105504 697564 337384 697592
rect 105504 697552 105510 697564
rect 337378 697552 337384 697564
rect 337436 697552 337442 697604
rect 525058 696940 525064 696992
rect 525116 696980 525122 696992
rect 580166 696980 580172 696992
rect 525116 696952 580172 696980
rect 525116 696940 525122 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 267642 694764 267648 694816
rect 267700 694804 267706 694816
rect 427078 694804 427084 694816
rect 267700 694776 427084 694804
rect 267700 694764 267706 694776
rect 427078 694764 427084 694776
rect 427136 694764 427142 694816
rect 316126 683136 316132 683188
rect 316184 683176 316190 683188
rect 580166 683176 580172 683188
rect 316184 683148 580172 683176
rect 316184 683136 316190 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 403710 670692 403716 670744
rect 403768 670732 403774 670744
rect 580166 670732 580172 670744
rect 403768 670704 580172 670732
rect 403768 670692 403774 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3234 667156 3240 667208
rect 3292 667196 3298 667208
rect 479518 667196 479524 667208
rect 3292 667168 479524 667196
rect 3292 667156 3298 667168
rect 479518 667156 479524 667168
rect 479576 667156 479582 667208
rect 40034 665796 40040 665848
rect 40092 665836 40098 665848
rect 476942 665836 476948 665848
rect 40092 665808 476948 665836
rect 40092 665796 40098 665808
rect 476942 665796 476948 665808
rect 477000 665796 477006 665848
rect 46566 663756 46572 663808
rect 46624 663796 46630 663808
rect 352834 663796 352840 663808
rect 46624 663768 352840 663796
rect 46624 663756 46630 663768
rect 352834 663756 352840 663768
rect 352892 663756 352898 663808
rect 51994 663144 52000 663196
rect 52052 663184 52058 663196
rect 276658 663184 276664 663196
rect 52052 663156 276664 663184
rect 52052 663144 52058 663156
rect 276658 663144 276664 663156
rect 276716 663144 276722 663196
rect 51902 663076 51908 663128
rect 51960 663116 51966 663128
rect 276750 663116 276756 663128
rect 51960 663088 276756 663116
rect 51960 663076 51966 663088
rect 276750 663076 276756 663088
rect 276808 663076 276814 663128
rect 46658 663008 46664 663060
rect 46716 663048 46722 663060
rect 276842 663048 276848 663060
rect 46716 663020 276848 663048
rect 46716 663008 46722 663020
rect 276842 663008 276848 663020
rect 276900 663008 276906 663060
rect 52178 662940 52184 662992
rect 52236 662980 52242 662992
rect 353018 662980 353024 662992
rect 52236 662952 353024 662980
rect 52236 662940 52242 662952
rect 353018 662940 353024 662952
rect 353076 662940 353082 662992
rect 51166 662872 51172 662924
rect 51224 662912 51230 662924
rect 352650 662912 352656 662924
rect 51224 662884 352656 662912
rect 51224 662872 51230 662884
rect 352650 662872 352656 662884
rect 352708 662872 352714 662924
rect 47854 662804 47860 662856
rect 47912 662844 47918 662856
rect 349798 662844 349804 662856
rect 47912 662816 349804 662844
rect 47912 662804 47918 662816
rect 349798 662804 349804 662816
rect 349856 662804 349862 662856
rect 51074 662736 51080 662788
rect 51132 662776 51138 662788
rect 355410 662776 355416 662788
rect 51132 662748 355416 662776
rect 51132 662736 51138 662748
rect 355410 662736 355416 662748
rect 355468 662736 355474 662788
rect 50982 662668 50988 662720
rect 51040 662708 51046 662720
rect 355318 662708 355324 662720
rect 51040 662680 355324 662708
rect 51040 662668 51046 662680
rect 355318 662668 355324 662680
rect 355376 662668 355382 662720
rect 46474 662600 46480 662652
rect 46532 662640 46538 662652
rect 352742 662640 352748 662652
rect 46532 662612 352748 662640
rect 46532 662600 46538 662612
rect 352742 662600 352748 662612
rect 352800 662600 352806 662652
rect 45462 662532 45468 662584
rect 45520 662572 45526 662584
rect 352558 662572 352564 662584
rect 45520 662544 352564 662572
rect 45520 662532 45526 662544
rect 352558 662532 352564 662544
rect 352616 662532 352622 662584
rect 51810 662464 51816 662516
rect 51868 662504 51874 662516
rect 403250 662504 403256 662516
rect 51868 662476 403256 662504
rect 51868 662464 51874 662476
rect 403250 662464 403256 662476
rect 403308 662464 403314 662516
rect 46382 662396 46388 662448
rect 46440 662436 46446 662448
rect 405274 662436 405280 662448
rect 46440 662408 405280 662436
rect 46440 662396 46446 662408
rect 405274 662396 405280 662408
rect 405332 662396 405338 662448
rect 52086 661784 52092 661836
rect 52144 661824 52150 661836
rect 279510 661824 279516 661836
rect 52144 661796 279516 661824
rect 52144 661784 52150 661796
rect 279510 661784 279516 661796
rect 279568 661784 279574 661836
rect 218054 661716 218060 661768
rect 218112 661756 218118 661768
rect 521838 661756 521844 661768
rect 218112 661728 521844 661756
rect 218112 661716 218118 661728
rect 521838 661716 521844 661728
rect 521896 661716 521902 661768
rect 6914 661648 6920 661700
rect 6972 661688 6978 661700
rect 520734 661688 520740 661700
rect 6972 661660 520740 661688
rect 6972 661648 6978 661660
rect 520734 661648 520740 661660
rect 520792 661648 520798 661700
rect 48866 661580 48872 661632
rect 48924 661620 48930 661632
rect 279602 661620 279608 661632
rect 48924 661592 279608 661620
rect 48924 661580 48930 661592
rect 279602 661580 279608 661592
rect 279660 661580 279666 661632
rect 48498 661512 48504 661564
rect 48556 661552 48562 661564
rect 310514 661552 310520 661564
rect 48556 661524 310520 661552
rect 48556 661512 48562 661524
rect 310514 661512 310520 661524
rect 310572 661512 310578 661564
rect 50890 661444 50896 661496
rect 50948 661484 50954 661496
rect 356698 661484 356704 661496
rect 50948 661456 356704 661484
rect 50948 661444 50954 661456
rect 356698 661444 356704 661456
rect 356756 661444 356762 661496
rect 50798 661376 50804 661428
rect 50856 661416 50862 661428
rect 358814 661416 358820 661428
rect 50856 661388 358820 661416
rect 50856 661376 50862 661388
rect 358814 661376 358820 661388
rect 358872 661376 358878 661428
rect 50614 661308 50620 661360
rect 50672 661348 50678 661360
rect 401594 661348 401600 661360
rect 50672 661320 401600 661348
rect 50672 661308 50678 661320
rect 401594 661308 401600 661320
rect 401652 661308 401658 661360
rect 51718 661240 51724 661292
rect 51776 661280 51782 661292
rect 407114 661280 407120 661292
rect 51776 661252 407120 661280
rect 51776 661240 51782 661252
rect 407114 661240 407120 661252
rect 407172 661240 407178 661292
rect 50338 661172 50344 661224
rect 50396 661212 50402 661224
rect 478322 661212 478328 661224
rect 50396 661184 478328 661212
rect 50396 661172 50402 661184
rect 478322 661172 478328 661184
rect 478380 661172 478386 661224
rect 50522 661104 50528 661156
rect 50580 661144 50586 661156
rect 478414 661144 478420 661156
rect 50580 661116 478420 661144
rect 50580 661104 50586 661116
rect 478414 661104 478420 661116
rect 478472 661104 478478 661156
rect 3510 661036 3516 661088
rect 3568 661076 3574 661088
rect 522022 661076 522028 661088
rect 3568 661048 522028 661076
rect 3568 661036 3574 661048
rect 522022 661036 522028 661048
rect 522080 661036 522086 661088
rect 49602 660560 49608 660612
rect 49660 660600 49666 660612
rect 278130 660600 278136 660612
rect 49660 660572 278136 660600
rect 49660 660560 49666 660572
rect 278130 660560 278136 660572
rect 278188 660560 278194 660612
rect 50706 660492 50712 660544
rect 50764 660532 50770 660544
rect 279694 660532 279700 660544
rect 50764 660504 279700 660532
rect 50764 660492 50770 660504
rect 279694 660492 279700 660504
rect 279752 660492 279758 660544
rect 50430 660424 50436 660476
rect 50488 660464 50494 660476
rect 502334 660464 502340 660476
rect 50488 660436 502340 660464
rect 50488 660424 50494 660436
rect 502334 660424 502340 660436
rect 502392 660424 502398 660476
rect 49418 660356 49424 660408
rect 49476 660396 49482 660408
rect 279142 660396 279148 660408
rect 49476 660368 279148 660396
rect 49476 660356 49482 660368
rect 279142 660356 279148 660368
rect 279200 660356 279206 660408
rect 331214 660356 331220 660408
rect 331272 660396 331278 660408
rect 520458 660396 520464 660408
rect 331272 660368 520464 660396
rect 331272 660356 331278 660368
rect 520458 660356 520464 660368
rect 520516 660356 520522 660408
rect 49878 660288 49884 660340
rect 49936 660328 49942 660340
rect 507854 660328 507860 660340
rect 49936 660300 507860 660328
rect 49936 660288 49942 660300
rect 507854 660288 507860 660300
rect 507912 660288 507918 660340
rect 49510 660220 49516 660272
rect 49568 660260 49574 660272
rect 280062 660260 280068 660272
rect 49568 660232 280068 660260
rect 49568 660220 49574 660232
rect 280062 660220 280068 660232
rect 280120 660220 280126 660272
rect 48130 660152 48136 660204
rect 48188 660192 48194 660204
rect 279326 660192 279332 660204
rect 48188 660164 279332 660192
rect 48188 660152 48194 660164
rect 279326 660152 279332 660164
rect 279384 660152 279390 660204
rect 48038 660084 48044 660136
rect 48096 660124 48102 660136
rect 279234 660124 279240 660136
rect 48096 660096 279240 660124
rect 48096 660084 48102 660096
rect 279234 660084 279240 660096
rect 279292 660084 279298 660136
rect 48222 660016 48228 660068
rect 48280 660056 48286 660068
rect 279878 660056 279884 660068
rect 48280 660028 279884 660056
rect 48280 660016 48286 660028
rect 279878 660016 279884 660028
rect 279936 660016 279942 660068
rect 50246 659948 50252 660000
rect 50304 659988 50310 660000
rect 521654 659988 521660 660000
rect 50304 659960 521660 659988
rect 50304 659948 50310 659960
rect 521654 659948 521660 659960
rect 521712 659948 521718 660000
rect 3418 659880 3424 659932
rect 3476 659920 3482 659932
rect 478966 659920 478972 659932
rect 3476 659892 478972 659920
rect 3476 659880 3482 659892
rect 478966 659880 478972 659892
rect 479024 659880 479030 659932
rect 3326 659812 3332 659864
rect 3384 659852 3390 659864
rect 520366 659852 520372 659864
rect 3384 659824 520372 659852
rect 3384 659812 3390 659824
rect 520366 659812 520372 659824
rect 520424 659812 520430 659864
rect 49970 657976 49976 658028
rect 50028 658016 50034 658028
rect 50246 658016 50252 658028
rect 50028 657988 50252 658016
rect 50028 657976 50034 657988
rect 50246 657976 50252 657988
rect 50304 657976 50310 658028
rect 50522 657500 50528 657552
rect 50580 657540 50586 657552
rect 50890 657540 50896 657552
rect 50580 657512 50896 657540
rect 50580 657500 50586 657512
rect 50890 657500 50896 657512
rect 50948 657500 50954 657552
rect 49326 655052 49332 655104
rect 49384 655092 49390 655104
rect 49602 655092 49608 655104
rect 49384 655064 49608 655092
rect 49384 655052 49390 655064
rect 49602 655052 49608 655064
rect 49660 655052 49666 655104
rect 48682 652740 48688 652792
rect 48740 652780 48746 652792
rect 50154 652780 50160 652792
rect 48740 652752 50160 652780
rect 48740 652740 48746 652752
rect 50154 652740 50160 652752
rect 50212 652740 50218 652792
rect 50982 651380 50988 651432
rect 51040 651420 51046 651432
rect 52178 651420 52184 651432
rect 51040 651392 52184 651420
rect 51040 651380 51046 651392
rect 52178 651380 52184 651392
rect 52236 651380 52242 651432
rect 49418 648524 49424 648576
rect 49476 648564 49482 648576
rect 50062 648564 50068 648576
rect 49476 648536 50068 648564
rect 49476 648524 49482 648536
rect 50062 648524 50068 648536
rect 50120 648524 50126 648576
rect 254302 645872 254308 645924
rect 254360 645912 254366 645924
rect 257338 645912 257344 645924
rect 254360 645884 257344 645912
rect 254360 645872 254366 645884
rect 257338 645872 257344 645884
rect 257396 645872 257402 645924
rect 282914 643696 282920 643748
rect 282972 643736 282978 643748
rect 477034 643736 477040 643748
rect 282972 643708 477040 643736
rect 282972 643696 282978 643708
rect 477034 643696 477040 643708
rect 477092 643696 477098 643748
rect 534718 643084 534724 643136
rect 534776 643124 534782 643136
rect 580166 643124 580172 643136
rect 534776 643096 580172 643124
rect 534776 643084 534782 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 360930 642676 360936 642728
rect 360988 642716 360994 642728
rect 379422 642716 379428 642728
rect 360988 642688 379428 642716
rect 360988 642676 360994 642688
rect 379422 642676 379428 642688
rect 379480 642676 379486 642728
rect 370038 642608 370044 642660
rect 370096 642648 370102 642660
rect 403802 642648 403808 642660
rect 370096 642620 403808 642648
rect 370096 642608 370102 642620
rect 403802 642608 403808 642620
rect 403860 642608 403866 642660
rect 359550 642540 359556 642592
rect 359608 642580 359614 642592
rect 376110 642580 376116 642592
rect 359608 642552 376116 642580
rect 359608 642540 359614 642552
rect 376110 642540 376116 642552
rect 376168 642540 376174 642592
rect 392670 642540 392676 642592
rect 392728 642580 392734 642592
rect 400766 642580 400772 642592
rect 392728 642552 400772 642580
rect 392728 642540 392734 642552
rect 400766 642540 400772 642552
rect 400824 642540 400830 642592
rect 327718 642472 327724 642524
rect 327776 642512 327782 642524
rect 377766 642512 377772 642524
rect 327776 642484 377772 642512
rect 327776 642472 327782 642484
rect 377766 642472 377772 642484
rect 377824 642472 377830 642524
rect 389910 642472 389916 642524
rect 389968 642512 389974 642524
rect 399478 642512 399484 642524
rect 389968 642484 399484 642512
rect 389968 642472 389974 642484
rect 399478 642472 399484 642484
rect 399536 642472 399542 642524
rect 371142 642404 371148 642456
rect 371200 642444 371206 642456
rect 405366 642444 405372 642456
rect 371200 642416 405372 642444
rect 371200 642404 371206 642416
rect 405366 642404 405372 642416
rect 405424 642404 405430 642456
rect 287606 642336 287612 642388
rect 287664 642376 287670 642388
rect 349890 642376 349896 642388
rect 287664 642348 349896 642376
rect 287664 642336 287670 642348
rect 349890 642336 349896 642348
rect 349948 642336 349954 642388
rect 360838 642336 360844 642388
rect 360896 642376 360902 642388
rect 396534 642376 396540 642388
rect 360896 642348 396540 642376
rect 360896 642336 360902 642348
rect 396534 642336 396540 642348
rect 396592 642336 396598 642388
rect 293770 642268 293776 642320
rect 293828 642308 293834 642320
rect 321186 642308 321192 642320
rect 293828 642280 321192 642308
rect 293828 642268 293834 642280
rect 321186 642268 321192 642280
rect 321244 642268 321250 642320
rect 359458 642268 359464 642320
rect 359516 642308 359522 642320
rect 373350 642308 373356 642320
rect 359516 642280 373356 642308
rect 359516 642268 359522 642280
rect 373350 642268 373356 642280
rect 373408 642268 373414 642320
rect 373902 642268 373908 642320
rect 373960 642308 373966 642320
rect 400858 642308 400864 642320
rect 373960 642280 400864 642308
rect 373960 642268 373966 642280
rect 400858 642268 400864 642280
rect 400916 642268 400922 642320
rect 300762 642200 300768 642252
rect 300820 642240 300826 642252
rect 331858 642240 331864 642252
rect 300820 642212 331864 642240
rect 300820 642200 300826 642212
rect 331858 642200 331864 642212
rect 331916 642200 331922 642252
rect 358814 642200 358820 642252
rect 358872 642240 358878 642252
rect 388254 642240 388260 642252
rect 358872 642212 388260 642240
rect 358872 642200 358878 642212
rect 388254 642200 388260 642212
rect 388312 642200 388318 642252
rect 394326 642200 394332 642252
rect 394384 642240 394390 642252
rect 405182 642240 405188 642252
rect 394384 642212 405188 642240
rect 394384 642200 394390 642212
rect 405182 642200 405188 642212
rect 405240 642200 405246 642252
rect 295242 642132 295248 642184
rect 295300 642172 295306 642184
rect 329098 642172 329104 642184
rect 295300 642144 329104 642172
rect 295300 642132 295306 642144
rect 329098 642132 329104 642144
rect 329156 642132 329162 642184
rect 359734 642132 359740 642184
rect 359792 642172 359798 642184
rect 390462 642172 390468 642184
rect 359792 642144 390468 642172
rect 359792 642132 359798 642144
rect 390462 642132 390468 642144
rect 390520 642132 390526 642184
rect 393222 642132 393228 642184
rect 393280 642172 393286 642184
rect 400674 642172 400680 642184
rect 393280 642144 400680 642172
rect 393280 642132 393286 642144
rect 400674 642132 400680 642144
rect 400732 642132 400738 642184
rect 286502 642064 286508 642116
rect 286560 642104 286566 642116
rect 322290 642104 322296 642116
rect 286560 642076 322296 642104
rect 286560 642064 286566 642076
rect 322290 642064 322296 642076
rect 322348 642064 322354 642116
rect 357342 642064 357348 642116
rect 357400 642104 357406 642116
rect 388806 642104 388812 642116
rect 357400 642076 388812 642104
rect 357400 642064 357406 642076
rect 388806 642064 388812 642076
rect 388864 642064 388870 642116
rect 392118 642064 392124 642116
rect 392176 642104 392182 642116
rect 400398 642104 400404 642116
rect 392176 642076 400404 642104
rect 392176 642064 392182 642076
rect 400398 642064 400404 642076
rect 400456 642064 400462 642116
rect 282086 641996 282092 642048
rect 282144 642036 282150 642048
rect 319530 642036 319536 642048
rect 282144 642008 319536 642036
rect 282144 641996 282150 642008
rect 319530 641996 319536 642008
rect 319588 641996 319594 642048
rect 353110 641996 353116 642048
rect 353168 642036 353174 642048
rect 386598 642036 386604 642048
rect 353168 642008 386604 642036
rect 353168 641996 353174 642008
rect 386598 641996 386604 642008
rect 386656 641996 386662 642048
rect 387702 641996 387708 642048
rect 387760 642036 387766 642048
rect 399570 642036 399576 642048
rect 387760 642008 399576 642036
rect 387760 641996 387766 642008
rect 399570 641996 399576 642008
rect 399628 641996 399634 642048
rect 282730 641928 282736 641980
rect 282788 641968 282794 641980
rect 321002 641968 321008 641980
rect 282788 641940 321008 641968
rect 282788 641928 282794 641940
rect 321002 641928 321008 641940
rect 321060 641928 321066 641980
rect 355962 641928 355968 641980
rect 356020 641968 356026 641980
rect 391014 641968 391020 641980
rect 356020 641940 391020 641968
rect 356020 641928 356026 641940
rect 391014 641928 391020 641940
rect 391072 641928 391078 641980
rect 284202 641860 284208 641912
rect 284260 641900 284266 641912
rect 327810 641900 327816 641912
rect 284260 641872 327816 641900
rect 284260 641860 284266 641872
rect 327810 641860 327816 641872
rect 327868 641860 327874 641912
rect 360010 641860 360016 641912
rect 360068 641900 360074 641912
rect 371694 641900 371700 641912
rect 360068 641872 371700 641900
rect 360068 641860 360074 641872
rect 371694 641860 371700 641872
rect 371752 641860 371758 641912
rect 375282 641860 375288 641912
rect 375340 641900 375346 641912
rect 389358 641900 389364 641912
rect 375340 641872 389364 641900
rect 375340 641860 375346 641872
rect 389358 641860 389364 641872
rect 389416 641860 389422 641912
rect 394878 641860 394884 641912
rect 394936 641900 394942 641912
rect 400582 641900 400588 641912
rect 394936 641872 400588 641900
rect 394936 641860 394942 641872
rect 400582 641860 400588 641872
rect 400640 641860 400646 641912
rect 297542 641792 297548 641844
rect 297600 641832 297606 641844
rect 352926 641832 352932 641844
rect 297600 641804 352932 641832
rect 297600 641792 297606 641804
rect 352926 641792 352932 641804
rect 352984 641792 352990 641844
rect 358906 641792 358912 641844
rect 358964 641832 358970 641844
rect 366726 641832 366732 641844
rect 358964 641804 366732 641832
rect 358964 641792 358970 641804
rect 366726 641792 366732 641804
rect 366784 641792 366790 641844
rect 379514 641792 379520 641844
rect 379572 641832 379578 641844
rect 386046 641832 386052 641844
rect 379572 641804 386052 641832
rect 379572 641792 379578 641804
rect 386046 641792 386052 641804
rect 386104 641792 386110 641844
rect 393774 641792 393780 641844
rect 393832 641832 393838 641844
rect 399294 641832 399300 641844
rect 393832 641804 399300 641832
rect 393832 641792 393838 641804
rect 399294 641792 399300 641804
rect 399352 641792 399358 641844
rect 475378 641792 475384 641844
rect 475436 641832 475442 641844
rect 493226 641832 493232 641844
rect 475436 641804 493232 641832
rect 475436 641792 475442 641804
rect 493226 641792 493232 641804
rect 493284 641792 493290 641844
rect 49142 641724 49148 641776
rect 49200 641764 49206 641776
rect 50246 641764 50252 641776
rect 49200 641736 50252 641764
rect 49200 641724 49206 641736
rect 50246 641724 50252 641736
rect 50304 641724 50310 641776
rect 299290 641724 299296 641776
rect 299348 641764 299354 641776
rect 321094 641764 321100 641776
rect 299348 641736 321100 641764
rect 299348 641724 299354 641736
rect 321094 641724 321100 641736
rect 321152 641724 321158 641776
rect 349982 641724 349988 641776
rect 350040 641764 350046 641776
rect 363414 641764 363420 641776
rect 350040 641736 363420 641764
rect 350040 641724 350046 641736
rect 363414 641724 363420 641736
rect 363472 641724 363478 641776
rect 367002 641724 367008 641776
rect 367060 641764 367066 641776
rect 372246 641764 372252 641776
rect 367060 641736 372252 641764
rect 367060 641724 367066 641736
rect 372246 641724 372252 641736
rect 372304 641724 372310 641776
rect 378042 641724 378048 641776
rect 378100 641764 378106 641776
rect 384390 641764 384396 641776
rect 378100 641736 384396 641764
rect 378100 641724 378106 641736
rect 384390 641724 384396 641736
rect 384448 641724 384454 641776
rect 395430 641724 395436 641776
rect 395488 641764 395494 641776
rect 399662 641764 399668 641776
rect 395488 641736 399668 641764
rect 395488 641724 395494 641736
rect 399662 641724 399668 641736
rect 399720 641724 399726 641776
rect 406378 641724 406384 641776
rect 406436 641764 406442 641776
rect 510614 641764 510620 641776
rect 406436 641736 510620 641764
rect 406436 641724 406442 641736
rect 510614 641724 510620 641736
rect 510672 641724 510678 641776
rect 278682 640976 278688 641028
rect 278740 641016 278746 641028
rect 310054 641016 310060 641028
rect 278740 640988 310060 641016
rect 278740 640976 278746 640988
rect 310054 640976 310060 640988
rect 310112 640976 310118 641028
rect 315850 640976 315856 641028
rect 315908 641016 315914 641028
rect 523678 641016 523684 641028
rect 315908 640988 523684 641016
rect 315908 640976 315914 640988
rect 523678 640976 523684 640988
rect 523736 640976 523742 641028
rect 314102 640908 314108 640960
rect 314160 640948 314166 640960
rect 527818 640948 527824 640960
rect 314160 640920 527824 640948
rect 314160 640908 314166 640920
rect 527818 640908 527824 640920
rect 527876 640908 527882 640960
rect 359826 640840 359832 640892
rect 359884 640880 359890 640892
rect 381630 640880 381636 640892
rect 359884 640852 381636 640880
rect 359884 640840 359890 640852
rect 381630 640840 381636 640852
rect 381688 640840 381694 640892
rect 355502 640772 355508 640824
rect 355560 640812 355566 640824
rect 378318 640812 378324 640824
rect 355560 640784 378324 640812
rect 355560 640772 355566 640784
rect 378318 640772 378324 640784
rect 378376 640772 378382 640824
rect 357066 640704 357072 640756
rect 357124 640744 357130 640756
rect 384942 640744 384948 640756
rect 357124 640716 384948 640744
rect 357124 640704 357130 640716
rect 384942 640704 384948 640716
rect 385000 640704 385006 640756
rect 312998 640636 313004 640688
rect 313056 640676 313062 640688
rect 338758 640676 338764 640688
rect 313056 640648 338764 640676
rect 313056 640636 313062 640648
rect 338758 640636 338764 640648
rect 338816 640636 338822 640688
rect 372798 640636 372804 640688
rect 372856 640676 372862 640688
rect 400306 640676 400312 640688
rect 372856 640648 400312 640676
rect 372856 640636 372862 640648
rect 400306 640636 400312 640648
rect 400364 640636 400370 640688
rect 309686 640568 309692 640620
rect 309744 640608 309750 640620
rect 356974 640608 356980 640620
rect 309744 640580 356980 640608
rect 309744 640568 309750 640580
rect 356974 640568 356980 640580
rect 357032 640568 357038 640620
rect 357158 640568 357164 640620
rect 357216 640608 357222 640620
rect 385494 640608 385500 640620
rect 357216 640580 385500 640608
rect 357216 640568 357222 640580
rect 385494 640568 385500 640580
rect 385552 640568 385558 640620
rect 304810 640500 304816 640552
rect 304868 640540 304874 640552
rect 354030 640540 354036 640552
rect 304868 640512 354036 640540
rect 304868 640500 304874 640512
rect 354030 640500 354036 640512
rect 354088 640500 354094 640552
rect 354122 640500 354128 640552
rect 354180 640540 354186 640552
rect 383838 640540 383844 640552
rect 354180 640512 383844 640540
rect 354180 640500 354186 640512
rect 383838 640500 383844 640512
rect 383896 640500 383902 640552
rect 387150 640500 387156 640552
rect 387208 640540 387214 640552
rect 402330 640540 402336 640552
rect 387208 640512 402336 640540
rect 387208 640500 387214 640512
rect 402330 640500 402336 640512
rect 402388 640500 402394 640552
rect 254302 640432 254308 640484
rect 254360 640472 254366 640484
rect 257430 640472 257436 640484
rect 254360 640444 257436 640472
rect 254360 640432 254366 640444
rect 257430 640432 257436 640444
rect 257488 640432 257494 640484
rect 301958 640432 301964 640484
rect 302016 640472 302022 640484
rect 356790 640472 356796 640484
rect 302016 640444 356796 640472
rect 302016 640432 302022 640444
rect 356790 640432 356796 640444
rect 356848 640432 356854 640484
rect 364518 640432 364524 640484
rect 364576 640472 364582 640484
rect 400214 640472 400220 640484
rect 364576 640444 400220 640472
rect 364576 640432 364582 640444
rect 400214 640432 400220 640444
rect 400272 640432 400278 640484
rect 315206 640364 315212 640416
rect 315264 640404 315270 640416
rect 322382 640404 322388 640416
rect 315264 640376 322388 640404
rect 315264 640364 315270 640376
rect 322382 640364 322388 640376
rect 322440 640364 322446 640416
rect 361206 640364 361212 640416
rect 361264 640404 361270 640416
rect 379974 640404 379980 640416
rect 361264 640376 379980 640404
rect 361264 640364 361270 640376
rect 379974 640364 379980 640376
rect 380032 640364 380038 640416
rect 310330 640296 310336 640348
rect 310388 640336 310394 640348
rect 320818 640336 320824 640348
rect 310388 640308 320824 640336
rect 310388 640296 310394 640308
rect 320818 640296 320824 640308
rect 320876 640296 320882 640348
rect 361114 640296 361120 640348
rect 361172 640336 361178 640348
rect 382734 640336 382740 640348
rect 361172 640308 382740 640336
rect 361172 640296 361178 640308
rect 382734 640296 382740 640308
rect 382792 640296 382798 640348
rect 364978 639888 364984 639940
rect 365036 639928 365042 639940
rect 365254 639928 365260 639940
rect 365036 639900 365260 639928
rect 365036 639888 365042 639900
rect 365254 639888 365260 639900
rect 365312 639888 365318 639940
rect 367002 639860 367008 639872
rect 360166 639832 367008 639860
rect 358630 639752 358636 639804
rect 358688 639792 358694 639804
rect 360166 639792 360194 639832
rect 367002 639820 367008 639832
rect 367060 639820 367066 639872
rect 375282 639792 375288 639804
rect 358688 639764 360194 639792
rect 361592 639764 375288 639792
rect 358688 639752 358694 639764
rect 358446 639684 358452 639736
rect 358504 639724 358510 639736
rect 361592 639724 361620 639764
rect 375282 639752 375288 639764
rect 375340 639752 375346 639804
rect 358504 639696 361620 639724
rect 358504 639684 358510 639696
rect 362218 639684 362224 639736
rect 362276 639724 362282 639736
rect 374638 639724 374644 639736
rect 362276 639696 374644 639724
rect 362276 639684 362282 639696
rect 374638 639684 374644 639696
rect 374696 639684 374702 639736
rect 367554 639616 367560 639668
rect 367612 639656 367618 639668
rect 372522 639656 372528 639668
rect 367612 639628 372528 639656
rect 367612 639616 367618 639628
rect 372522 639616 372528 639628
rect 372580 639616 372586 639668
rect 399110 639656 399116 639668
rect 389146 639628 399116 639656
rect 357802 639548 357808 639600
rect 357860 639588 357866 639600
rect 376294 639588 376300 639600
rect 357860 639560 376300 639588
rect 357860 639548 357866 639560
rect 376294 639548 376300 639560
rect 376352 639548 376358 639600
rect 361482 639480 361488 639532
rect 361540 639520 361546 639532
rect 370222 639520 370228 639532
rect 361540 639492 370228 639520
rect 361540 639480 361546 639492
rect 370222 639480 370228 639492
rect 370280 639480 370286 639532
rect 302206 639424 307432 639452
rect 296438 639276 296444 639328
rect 296496 639316 296502 639328
rect 296496 639288 296714 639316
rect 296496 639276 296502 639288
rect 296686 639112 296714 639288
rect 302206 639112 302234 639424
rect 303062 639344 303068 639396
rect 303120 639384 303126 639396
rect 303120 639356 307340 639384
rect 303120 639344 303126 639356
rect 306282 639276 306288 639328
rect 306340 639276 306346 639328
rect 296686 639084 302234 639112
rect 306300 639044 306328 639276
rect 307312 639112 307340 639356
rect 307404 639180 307432 639424
rect 360102 639412 360108 639464
rect 360160 639452 360166 639464
rect 368198 639452 368204 639464
rect 360160 639424 368204 639452
rect 360160 639412 360166 639424
rect 368198 639412 368204 639424
rect 368256 639412 368262 639464
rect 369504 639424 372476 639452
rect 358538 639344 358544 639396
rect 358596 639384 358602 639396
rect 362218 639384 362224 639396
rect 358596 639356 362224 639384
rect 358596 639344 358602 639356
rect 362218 639344 362224 639356
rect 362276 639344 362282 639396
rect 364978 639344 364984 639396
rect 365036 639344 365042 639396
rect 365346 639344 365352 639396
rect 365404 639344 365410 639396
rect 366450 639344 366456 639396
rect 366508 639344 366514 639396
rect 311710 639276 311716 639328
rect 311768 639316 311774 639328
rect 324958 639316 324964 639328
rect 311768 639288 324964 639316
rect 311768 639276 311774 639288
rect 324958 639276 324964 639288
rect 325016 639276 325022 639328
rect 322198 639180 322204 639192
rect 307404 639152 322204 639180
rect 322198 639140 322204 639152
rect 322256 639140 322262 639192
rect 353938 639112 353944 639124
rect 307312 639084 353944 639112
rect 353938 639072 353944 639084
rect 353996 639072 354002 639124
rect 356882 639044 356888 639056
rect 306300 639016 356888 639044
rect 356882 639004 356888 639016
rect 356940 639004 356946 639056
rect 278774 638936 278780 638988
rect 278832 638976 278838 638988
rect 361574 638976 361580 638988
rect 278832 638948 361580 638976
rect 278832 638936 278838 638948
rect 361574 638936 361580 638948
rect 361632 638936 361638 638988
rect 364996 638976 365024 639344
rect 365364 639044 365392 639344
rect 366468 639248 366496 639344
rect 366468 639220 367094 639248
rect 367066 639112 367094 639220
rect 369504 639112 369532 639424
rect 369670 639344 369676 639396
rect 369728 639344 369734 639396
rect 369688 639316 369716 639344
rect 369688 639288 372292 639316
rect 367066 639084 369532 639112
rect 372264 639112 372292 639288
rect 372448 639180 372476 639424
rect 374730 639412 374736 639464
rect 374788 639452 374794 639464
rect 374788 639424 377444 639452
rect 374788 639412 374794 639424
rect 372522 639344 372528 639396
rect 372580 639344 372586 639396
rect 375834 639344 375840 639396
rect 375892 639344 375898 639396
rect 377416 639384 377444 639424
rect 377490 639412 377496 639464
rect 377548 639452 377554 639464
rect 389146 639452 389174 639628
rect 399110 639616 399116 639628
rect 399168 639616 399174 639668
rect 396166 639548 396172 639600
rect 396224 639588 396230 639600
rect 399018 639588 399024 639600
rect 396224 639560 399024 639588
rect 396224 639548 396230 639560
rect 399018 639548 399024 639560
rect 399076 639548 399082 639600
rect 391198 639480 391204 639532
rect 391256 639520 391262 639532
rect 404630 639520 404636 639532
rect 391256 639492 404636 639520
rect 391256 639480 391262 639492
rect 404630 639480 404636 639492
rect 404688 639480 404694 639532
rect 377548 639424 389174 639452
rect 390296 639424 396074 639452
rect 377548 639412 377554 639424
rect 390296 639384 390324 639424
rect 377416 639356 390324 639384
rect 391198 639344 391204 639396
rect 391256 639344 391262 639396
rect 372540 639248 372568 639344
rect 375852 639316 375880 639344
rect 391216 639316 391244 639344
rect 375852 639288 391244 639316
rect 396046 639316 396074 639424
rect 397914 639412 397920 639464
rect 397972 639452 397978 639464
rect 398926 639452 398932 639464
rect 397972 639424 398932 639452
rect 397972 639412 397978 639424
rect 398926 639412 398932 639424
rect 398984 639412 398990 639464
rect 403158 639316 403164 639328
rect 396046 639288 403164 639316
rect 403158 639276 403164 639288
rect 403216 639276 403222 639328
rect 399938 639248 399944 639260
rect 372540 639220 399944 639248
rect 399938 639208 399944 639220
rect 399996 639208 400002 639260
rect 400490 639180 400496 639192
rect 372448 639152 400496 639180
rect 400490 639140 400496 639152
rect 400548 639140 400554 639192
rect 403894 639112 403900 639124
rect 372264 639084 403900 639112
rect 403894 639072 403900 639084
rect 403952 639072 403958 639124
rect 402146 639044 402152 639056
rect 365364 639016 402152 639044
rect 402146 639004 402152 639016
rect 402204 639004 402210 639056
rect 401778 638976 401784 638988
rect 364996 638948 401784 638976
rect 401778 638936 401784 638948
rect 401836 638936 401842 638988
rect 403618 634788 403624 634840
rect 403676 634828 403682 634840
rect 477678 634828 477684 634840
rect 403676 634800 477684 634828
rect 403676 634788 403682 634800
rect 477678 634788 477684 634800
rect 477736 634788 477742 634840
rect 254670 633428 254676 633480
rect 254728 633468 254734 633480
rect 269850 633468 269856 633480
rect 254728 633440 269856 633468
rect 254728 633428 254734 633440
rect 269850 633428 269856 633440
rect 269908 633428 269914 633480
rect 523678 632000 523684 632052
rect 523736 632040 523742 632052
rect 580166 632040 580172 632052
rect 523736 632012 580172 632040
rect 523736 632000 523742 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 49326 629688 49332 629740
rect 49384 629728 49390 629740
rect 52086 629728 52092 629740
rect 49384 629700 52092 629728
rect 49384 629688 49390 629700
rect 52086 629688 52092 629700
rect 52144 629688 52150 629740
rect 254670 627920 254676 627972
rect 254728 627960 254734 627972
rect 275370 627960 275376 627972
rect 254728 627932 275376 627960
rect 254728 627920 254734 627932
rect 275370 627920 275376 627932
rect 275428 627920 275434 627972
rect 48866 618944 48872 618996
rect 48924 618984 48930 618996
rect 51994 618984 52000 618996
rect 48924 618956 52000 618984
rect 48924 618944 48930 618956
rect 51994 618944 52000 618956
rect 52052 618944 52058 618996
rect 254394 616836 254400 616888
rect 254452 616876 254458 616888
rect 264238 616876 264244 616888
rect 254452 616848 264244 616876
rect 254452 616836 254458 616848
rect 264238 616836 264244 616848
rect 264296 616836 264302 616888
rect 538858 616836 538864 616888
rect 538916 616876 538922 616888
rect 580166 616876 580172 616888
rect 538916 616848 580172 616876
rect 538916 616836 538922 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 48774 612756 48780 612808
rect 48832 612796 48838 612808
rect 51902 612796 51908 612808
rect 48832 612768 51908 612796
rect 48832 612756 48838 612768
rect 51902 612756 51908 612768
rect 51960 612756 51966 612808
rect 254486 611328 254492 611380
rect 254544 611368 254550 611380
rect 273898 611368 273904 611380
rect 254544 611340 273904 611368
rect 254544 611328 254550 611340
rect 273898 611328 273904 611340
rect 273956 611328 273962 611380
rect 254210 604460 254216 604512
rect 254268 604500 254274 604512
rect 271138 604500 271144 604512
rect 254268 604472 271144 604500
rect 254268 604460 254274 604472
rect 271138 604460 271144 604472
rect 271196 604460 271202 604512
rect 398374 600244 398380 600296
rect 398432 600284 398438 600296
rect 403618 600284 403624 600296
rect 398432 600256 403624 600284
rect 398432 600244 398438 600256
rect 403618 600244 403624 600256
rect 403676 600244 403682 600296
rect 391934 599972 391940 600024
rect 391992 600012 391998 600024
rect 392302 600012 392308 600024
rect 391992 599984 392308 600012
rect 391992 599972 391998 599984
rect 392302 599972 392308 599984
rect 392360 599972 392366 600024
rect 301958 599904 301964 599956
rect 302016 599944 302022 599956
rect 302188 599944 302194 599956
rect 302016 599916 302194 599944
rect 302016 599904 302022 599916
rect 302188 599904 302194 599916
rect 302246 599904 302252 599956
rect 296714 599836 296720 599888
rect 296772 599876 296778 599888
rect 297772 599876 297778 599888
rect 296772 599848 297778 599876
rect 296772 599836 296778 599848
rect 297772 599836 297778 599848
rect 297830 599836 297836 599888
rect 298094 599836 298100 599888
rect 298152 599876 298158 599888
rect 299428 599876 299434 599888
rect 298152 599848 299434 599876
rect 298152 599836 298158 599848
rect 299428 599836 299434 599848
rect 299486 599836 299492 599888
rect 392302 599836 392308 599888
rect 392360 599876 392366 599888
rect 399202 599876 399208 599888
rect 392360 599848 399208 599876
rect 392360 599836 392366 599848
rect 399202 599836 399208 599848
rect 399260 599836 399266 599888
rect 382274 599768 382280 599820
rect 382332 599808 382338 599820
rect 400582 599808 400588 599820
rect 382332 599780 400588 599808
rect 382332 599768 382338 599780
rect 400582 599768 400588 599780
rect 400640 599768 400646 599820
rect 378502 599700 378508 599752
rect 378560 599740 378566 599752
rect 400766 599740 400772 599752
rect 378560 599712 400772 599740
rect 378560 599700 378566 599712
rect 400766 599700 400772 599712
rect 400824 599700 400830 599752
rect 372614 599632 372620 599684
rect 372672 599672 372678 599684
rect 399294 599672 399300 599684
rect 372672 599644 399300 599672
rect 372672 599632 372678 599644
rect 399294 599632 399300 599644
rect 399352 599632 399358 599684
rect 254578 599564 254584 599616
rect 254636 599604 254642 599616
rect 320174 599604 320180 599616
rect 254636 599576 320180 599604
rect 254636 599564 254642 599576
rect 320174 599564 320180 599576
rect 320232 599564 320238 599616
rect 365714 599564 365720 599616
rect 365772 599604 365778 599616
rect 400674 599604 400680 599616
rect 365772 599576 400680 599604
rect 365772 599564 365778 599576
rect 400674 599564 400680 599576
rect 400732 599564 400738 599616
rect 297818 599224 297824 599276
rect 297876 599264 297882 599276
rect 327718 599264 327724 599276
rect 297876 599236 327724 599264
rect 297876 599224 297882 599236
rect 327718 599224 327724 599236
rect 327776 599224 327782 599276
rect 300854 599156 300860 599208
rect 300912 599196 300918 599208
rect 301958 599196 301964 599208
rect 300912 599168 301964 599196
rect 300912 599156 300918 599168
rect 301958 599156 301964 599168
rect 302016 599196 302022 599208
rect 331950 599196 331956 599208
rect 302016 599168 331956 599196
rect 302016 599156 302022 599168
rect 331950 599156 331956 599168
rect 332008 599156 332014 599208
rect 306374 599088 306380 599140
rect 306432 599128 306438 599140
rect 306742 599128 306748 599140
rect 306432 599100 306748 599128
rect 306432 599088 306438 599100
rect 306742 599088 306748 599100
rect 306800 599128 306806 599140
rect 353110 599128 353116 599140
rect 306800 599100 353116 599128
rect 306800 599088 306806 599100
rect 353110 599088 353116 599100
rect 353168 599088 353174 599140
rect 387702 599088 387708 599140
rect 387760 599128 387766 599140
rect 406378 599128 406384 599140
rect 387760 599100 406384 599128
rect 387760 599088 387766 599100
rect 406378 599088 406384 599100
rect 406436 599088 406442 599140
rect 299382 599020 299388 599072
rect 299440 599060 299446 599072
rect 360930 599060 360936 599072
rect 299440 599032 360936 599060
rect 299440 599020 299446 599032
rect 360930 599020 360936 599032
rect 360988 599020 360994 599072
rect 361758 599020 361764 599072
rect 361816 599060 361822 599072
rect 475378 599060 475384 599072
rect 361816 599032 475384 599060
rect 361816 599020 361822 599032
rect 475378 599020 475384 599032
rect 475436 599020 475442 599072
rect 283006 598952 283012 599004
rect 283064 598992 283070 599004
rect 349982 598992 349988 599004
rect 283064 598964 349988 598992
rect 283064 598952 283070 598964
rect 349982 598952 349988 598964
rect 350040 598952 350046 599004
rect 254762 598884 254768 598936
rect 254820 598924 254826 598936
rect 361776 598924 361804 599020
rect 386598 598952 386604 599004
rect 386656 598992 386662 599004
rect 387702 598992 387708 599004
rect 386656 598964 387708 598992
rect 386656 598952 386662 598964
rect 387702 598952 387708 598964
rect 387760 598952 387766 599004
rect 254820 598896 361804 598924
rect 254820 598884 254826 598896
rect 388254 598884 388260 598936
rect 388312 598924 388318 598936
rect 521746 598924 521752 598936
rect 388312 598896 521752 598924
rect 388312 598884 388318 598896
rect 521746 598884 521752 598896
rect 521804 598884 521810 598936
rect 302142 598816 302148 598868
rect 302200 598856 302206 598868
rect 302200 598828 311204 598856
rect 302200 598816 302206 598828
rect 303522 598748 303528 598800
rect 303580 598788 303586 598800
rect 311176 598788 311204 598828
rect 311250 598816 311256 598868
rect 311308 598856 311314 598868
rect 361206 598856 361212 598868
rect 311308 598828 361212 598856
rect 311308 598816 311314 598828
rect 361206 598816 361212 598828
rect 361264 598816 361270 598868
rect 386414 598816 386420 598868
rect 386472 598856 386478 598868
rect 387150 598856 387156 598868
rect 386472 598828 387156 598856
rect 386472 598816 386478 598828
rect 387150 598816 387156 598828
rect 387208 598856 387214 598868
rect 513834 598856 513840 598868
rect 387208 598828 513840 598856
rect 387208 598816 387214 598828
rect 513834 598816 513840 598828
rect 513892 598816 513898 598868
rect 359826 598788 359832 598800
rect 303580 598760 311112 598788
rect 311176 598760 359832 598788
rect 303580 598748 303586 598760
rect 311084 598720 311112 598760
rect 359826 598748 359832 598760
rect 359884 598748 359890 598800
rect 388438 598748 388444 598800
rect 388496 598788 388502 598800
rect 478138 598788 478144 598800
rect 388496 598760 478144 598788
rect 388496 598748 388502 598760
rect 478138 598748 478144 598760
rect 478196 598748 478202 598800
rect 361114 598720 361120 598732
rect 311084 598692 361120 598720
rect 361114 598680 361120 598692
rect 361172 598680 361178 598732
rect 286870 598612 286876 598664
rect 286928 598652 286934 598664
rect 289170 598652 289176 598664
rect 286928 598624 289176 598652
rect 286928 598612 286934 598624
rect 289170 598612 289176 598624
rect 289228 598612 289234 598664
rect 292482 598612 292488 598664
rect 292540 598652 292546 598664
rect 297450 598652 297456 598664
rect 292540 598624 297456 598652
rect 292540 598612 292546 598624
rect 297450 598612 297456 598624
rect 297508 598612 297514 598664
rect 304902 598612 304908 598664
rect 304960 598652 304966 598664
rect 357066 598652 357072 598664
rect 304960 598624 357072 598652
rect 304960 598612 304966 598624
rect 357066 598612 357072 598624
rect 357124 598612 357130 598664
rect 361022 598612 361028 598664
rect 361080 598652 361086 598664
rect 380526 598652 380532 598664
rect 361080 598624 380532 598652
rect 361080 598612 361086 598624
rect 380526 598612 380532 598624
rect 380584 598612 380590 598664
rect 289786 598556 302234 598584
rect 285122 598408 285128 598460
rect 285180 598448 285186 598460
rect 289786 598448 289814 598556
rect 285180 598420 289814 598448
rect 302206 598448 302234 598556
rect 305822 598544 305828 598596
rect 305880 598584 305886 598596
rect 306282 598584 306288 598596
rect 305880 598556 306288 598584
rect 305880 598544 305886 598556
rect 306282 598544 306288 598556
rect 306340 598584 306346 598596
rect 357158 598584 357164 598596
rect 306340 598556 357164 598584
rect 306340 598544 306346 598556
rect 357158 598544 357164 598556
rect 357216 598544 357222 598596
rect 359642 598544 359648 598596
rect 359700 598584 359706 598596
rect 382182 598584 382188 598596
rect 359700 598556 382188 598584
rect 359700 598544 359706 598556
rect 382182 598544 382188 598556
rect 382240 598544 382246 598596
rect 388254 598544 388260 598596
rect 388312 598584 388318 598596
rect 388530 598584 388536 598596
rect 388312 598556 388536 598584
rect 388312 598544 388318 598556
rect 388530 598544 388536 598556
rect 388588 598544 388594 598596
rect 304166 598476 304172 598528
rect 304224 598516 304230 598528
rect 354122 598516 354128 598528
rect 304224 598488 354128 598516
rect 304224 598476 304230 598488
rect 354122 598476 354128 598488
rect 354180 598476 354186 598528
rect 360930 598476 360936 598528
rect 360988 598516 360994 598528
rect 391566 598516 391572 598528
rect 360988 598488 391572 598516
rect 360988 598476 360994 598488
rect 391566 598476 391572 598488
rect 391624 598476 391630 598528
rect 320910 598448 320916 598460
rect 302206 598420 320916 598448
rect 285180 598408 285186 598420
rect 320910 598408 320916 598420
rect 320968 598408 320974 598460
rect 366174 598408 366180 598460
rect 366232 598448 366238 598460
rect 397730 598448 397736 598460
rect 366232 598420 397736 598448
rect 366232 598408 366238 598420
rect 397730 598408 397736 598420
rect 397788 598408 397794 598460
rect 288986 598340 288992 598392
rect 289044 598380 289050 598392
rect 289044 598352 297404 598380
rect 289044 598340 289050 598352
rect 290090 598204 290096 598256
rect 290148 598244 290154 598256
rect 297376 598244 297404 598352
rect 297450 598340 297456 598392
rect 297508 598380 297514 598392
rect 297508 598352 302234 598380
rect 297508 598340 297514 598352
rect 302206 598312 302234 598352
rect 303062 598340 303068 598392
rect 303120 598380 303126 598392
rect 303522 598380 303528 598392
rect 303120 598352 303528 598380
rect 303120 598340 303126 598352
rect 303522 598340 303528 598352
rect 303580 598340 303586 598392
rect 303614 598340 303620 598392
rect 303672 598380 303678 598392
rect 355502 598380 355508 598392
rect 303672 598352 355508 598380
rect 303672 598340 303678 598352
rect 355502 598340 355508 598352
rect 355560 598340 355566 598392
rect 363414 598340 363420 598392
rect 363472 598380 363478 598392
rect 398098 598380 398104 598392
rect 363472 598352 398104 598380
rect 363472 598340 363478 598352
rect 398098 598340 398104 598352
rect 398156 598340 398162 598392
rect 404722 598312 404728 598324
rect 302206 598284 404728 598312
rect 404722 598272 404728 598284
rect 404780 598272 404786 598324
rect 404814 598244 404820 598256
rect 290148 598216 292574 598244
rect 297376 598216 404820 598244
rect 290148 598204 290154 598216
rect 287054 598136 287060 598188
rect 287112 598176 287118 598188
rect 287514 598176 287520 598188
rect 287112 598148 287520 598176
rect 287112 598136 287118 598148
rect 287514 598136 287520 598148
rect 287572 598136 287578 598188
rect 291102 598136 291108 598188
rect 291160 598176 291166 598188
rect 291838 598176 291844 598188
rect 291160 598148 291844 598176
rect 291160 598136 291166 598148
rect 291838 598136 291844 598148
rect 291896 598136 291902 598188
rect 292546 598176 292574 598216
rect 404814 598204 404820 598216
rect 404872 598204 404878 598256
rect 472802 598204 472808 598256
rect 472860 598244 472866 598256
rect 496446 598244 496452 598256
rect 472860 598216 496452 598244
rect 472860 598204 472866 598216
rect 496446 598204 496452 598216
rect 496504 598204 496510 598256
rect 323670 598176 323676 598188
rect 292546 598148 323676 598176
rect 323670 598136 323676 598148
rect 323728 598136 323734 598188
rect 369854 598136 369860 598188
rect 369912 598176 369918 598188
rect 370222 598176 370228 598188
rect 369912 598148 370228 598176
rect 369912 598136 369918 598148
rect 370222 598136 370228 598148
rect 370280 598136 370286 598188
rect 372706 598136 372712 598188
rect 372764 598176 372770 598188
rect 373534 598176 373540 598188
rect 372764 598148 373540 598176
rect 372764 598136 372770 598148
rect 373534 598136 373540 598148
rect 373592 598136 373598 598188
rect 378410 598136 378416 598188
rect 378468 598176 378474 598188
rect 379054 598176 379060 598188
rect 378468 598148 379060 598176
rect 378468 598136 378474 598148
rect 379054 598136 379060 598148
rect 379112 598136 379118 598188
rect 380986 598136 380992 598188
rect 381044 598176 381050 598188
rect 381262 598176 381268 598188
rect 381044 598148 381268 598176
rect 381044 598136 381050 598148
rect 381262 598136 381268 598148
rect 381320 598136 381326 598188
rect 389266 598136 389272 598188
rect 389324 598176 389330 598188
rect 389542 598176 389548 598188
rect 389324 598148 389548 598176
rect 389324 598136 389330 598148
rect 389542 598136 389548 598148
rect 389600 598136 389606 598188
rect 393314 598136 393320 598188
rect 393372 598176 393378 598188
rect 393958 598176 393964 598188
rect 393372 598148 393964 598176
rect 393372 598136 393378 598148
rect 393958 598136 393964 598148
rect 394016 598136 394022 598188
rect 396074 598136 396080 598188
rect 396132 598176 396138 598188
rect 396718 598176 396724 598188
rect 396132 598148 396724 598176
rect 396132 598136 396138 598148
rect 396718 598136 396724 598148
rect 396776 598136 396782 598188
rect 298646 598068 298652 598120
rect 298704 598108 298710 598120
rect 300670 598108 300676 598120
rect 298704 598080 300676 598108
rect 298704 598068 298710 598080
rect 300670 598068 300676 598080
rect 300728 598108 300734 598120
rect 303614 598108 303620 598120
rect 300728 598080 303620 598108
rect 300728 598068 300734 598080
rect 303614 598068 303620 598080
rect 303672 598068 303678 598120
rect 304166 598068 304172 598120
rect 304224 598108 304230 598120
rect 304810 598108 304816 598120
rect 304224 598080 304816 598108
rect 304224 598068 304230 598080
rect 304810 598068 304816 598080
rect 304868 598068 304874 598120
rect 306466 598068 306472 598120
rect 306524 598108 306530 598120
rect 307386 598108 307392 598120
rect 306524 598080 307392 598108
rect 306524 598068 306530 598080
rect 307386 598068 307392 598080
rect 307444 598068 307450 598120
rect 309134 598068 309140 598120
rect 309192 598108 309198 598120
rect 310146 598108 310152 598120
rect 309192 598080 310152 598108
rect 309192 598068 309198 598080
rect 310146 598068 310152 598080
rect 310204 598068 310210 598120
rect 311894 598068 311900 598120
rect 311952 598108 311958 598120
rect 312354 598108 312360 598120
rect 311952 598080 312360 598108
rect 311952 598068 311958 598080
rect 312354 598068 312360 598080
rect 312412 598068 312418 598120
rect 313274 598068 313280 598120
rect 313332 598108 313338 598120
rect 314010 598108 314016 598120
rect 313332 598080 314016 598108
rect 313332 598068 313338 598080
rect 314010 598068 314016 598080
rect 314068 598068 314074 598120
rect 314654 598068 314660 598120
rect 314712 598108 314718 598120
rect 315114 598108 315120 598120
rect 314712 598080 315120 598108
rect 314712 598068 314718 598080
rect 315114 598068 315120 598080
rect 315172 598068 315178 598120
rect 389174 598068 389180 598120
rect 389232 598108 389238 598120
rect 390094 598108 390100 598120
rect 389232 598080 390100 598108
rect 389232 598068 389238 598080
rect 390094 598068 390100 598080
rect 390152 598068 390158 598120
rect 392026 598068 392032 598120
rect 392084 598108 392090 598120
rect 392854 598108 392860 598120
rect 392084 598080 392860 598108
rect 392084 598068 392090 598080
rect 392854 598068 392860 598080
rect 392912 598068 392918 598120
rect 300302 598000 300308 598052
rect 300360 598040 300366 598052
rect 300578 598040 300584 598052
rect 300360 598012 300584 598040
rect 300360 598000 300366 598012
rect 300578 598000 300584 598012
rect 300636 598040 300642 598052
rect 311250 598040 311256 598052
rect 300636 598012 311256 598040
rect 300636 598000 300642 598012
rect 311250 598000 311256 598012
rect 311308 598000 311314 598052
rect 314746 598000 314752 598052
rect 314804 598040 314810 598052
rect 315666 598040 315672 598052
rect 314804 598012 315672 598040
rect 314804 598000 314810 598012
rect 315666 598000 315672 598012
rect 315724 598000 315730 598052
rect 308306 597932 308312 597984
rect 308364 597972 308370 597984
rect 323578 597972 323584 597984
rect 308364 597944 323584 597972
rect 308364 597932 308370 597944
rect 323578 597932 323584 597944
rect 323636 597932 323642 597984
rect 395430 597796 395436 597848
rect 395488 597836 395494 597848
rect 400582 597836 400588 597848
rect 395488 597808 400588 597836
rect 395488 597796 395494 597808
rect 400582 597796 400588 597808
rect 400640 597796 400646 597848
rect 362862 597524 362868 597576
rect 362920 597564 362926 597576
rect 368658 597564 368664 597576
rect 362920 597536 368664 597564
rect 362920 597524 362926 597536
rect 368658 597524 368664 597536
rect 368716 597524 368722 597576
rect 383654 597184 383660 597236
rect 383712 597224 383718 597236
rect 384574 597224 384580 597236
rect 383712 597196 384580 597224
rect 383712 597184 383718 597196
rect 384574 597184 384580 597196
rect 384632 597184 384638 597236
rect 282914 597048 282920 597100
rect 282972 597088 282978 597100
rect 283650 597088 283656 597100
rect 282972 597060 283656 597088
rect 282972 597048 282978 597060
rect 283650 597048 283656 597060
rect 283708 597048 283714 597100
rect 313182 596912 313188 596964
rect 313240 596952 313246 596964
rect 337470 596952 337476 596964
rect 313240 596924 337476 596952
rect 313240 596912 313246 596924
rect 337470 596912 337476 596924
rect 337528 596912 337534 596964
rect 347682 596912 347688 596964
rect 347740 596952 347746 596964
rect 375558 596952 375564 596964
rect 347740 596924 375564 596952
rect 347740 596912 347746 596924
rect 375558 596912 375564 596924
rect 375616 596912 375622 596964
rect 253382 596844 253388 596896
rect 253440 596884 253446 596896
rect 502334 596884 502340 596896
rect 253440 596856 502340 596884
rect 253440 596844 253446 596856
rect 502334 596844 502340 596856
rect 502392 596844 502398 596896
rect 325602 596776 325608 596828
rect 325660 596816 325666 596828
rect 398190 596816 398196 596828
rect 325660 596788 398196 596816
rect 325660 596776 325666 596788
rect 398190 596776 398196 596788
rect 398248 596776 398254 596828
rect 468662 596776 468668 596828
rect 468720 596816 468726 596828
rect 479702 596816 479708 596828
rect 468720 596788 479708 596816
rect 468720 596776 468726 596788
rect 479702 596776 479708 596788
rect 479760 596776 479766 596828
rect 367278 596368 367284 596420
rect 367336 596368 367342 596420
rect 367296 596216 367324 596368
rect 367278 596164 367284 596216
rect 367336 596164 367342 596216
rect 320174 596096 320180 596148
rect 320232 596136 320238 596148
rect 325602 596136 325608 596148
rect 320232 596108 325608 596136
rect 320232 596096 320238 596108
rect 325602 596096 325608 596108
rect 325660 596096 325666 596148
rect 292574 596028 292580 596080
rect 292632 596068 292638 596080
rect 293586 596068 293592 596080
rect 292632 596040 293592 596068
rect 292632 596028 292638 596040
rect 293586 596028 293592 596040
rect 293644 596028 293650 596080
rect 364426 596028 364432 596080
rect 364484 596068 364490 596080
rect 365254 596068 365260 596080
rect 364484 596040 365260 596068
rect 364484 596028 364490 596040
rect 365254 596028 365260 596040
rect 365312 596028 365318 596080
rect 367094 596028 367100 596080
rect 367152 596068 367158 596080
rect 368014 596068 368020 596080
rect 367152 596040 368020 596068
rect 367152 596028 367158 596040
rect 368014 596028 368020 596040
rect 368072 596028 368078 596080
rect 297542 595484 297548 595536
rect 297600 595524 297606 595536
rect 341518 595524 341524 595536
rect 297600 595496 341524 595524
rect 297600 595484 297606 595496
rect 341518 595484 341524 595496
rect 341576 595484 341582 595536
rect 349982 595484 349988 595536
rect 350040 595524 350046 595536
rect 363966 595524 363972 595536
rect 350040 595496 363972 595524
rect 350040 595484 350046 595496
rect 363966 595484 363972 595496
rect 364024 595484 364030 595536
rect 372890 595484 372896 595536
rect 372948 595524 372954 595536
rect 383838 595524 383844 595536
rect 372948 595496 383844 595524
rect 372948 595484 372954 595496
rect 383838 595484 383844 595496
rect 383896 595484 383902 595536
rect 253290 595416 253296 595468
rect 253348 595456 253354 595468
rect 503714 595456 503720 595468
rect 253348 595428 503720 595456
rect 253348 595416 253354 595428
rect 503714 595416 503720 595428
rect 503772 595416 503778 595468
rect 383930 595212 383936 595264
rect 383988 595252 383994 595264
rect 392578 595252 392584 595264
rect 383988 595224 392584 595252
rect 383988 595212 383994 595224
rect 392578 595212 392584 595224
rect 392636 595212 392642 595264
rect 49510 594804 49516 594856
rect 49568 594844 49574 594856
rect 51718 594844 51724 594856
rect 49568 594816 51724 594844
rect 49568 594804 49574 594816
rect 51718 594804 51724 594816
rect 51776 594804 51782 594856
rect 307018 594124 307024 594176
rect 307076 594164 307082 594176
rect 327718 594164 327724 594176
rect 307076 594136 327724 594164
rect 307076 594124 307082 594136
rect 327718 594124 327724 594136
rect 327776 594124 327782 594176
rect 343542 594124 343548 594176
rect 343600 594164 343606 594176
rect 371786 594164 371792 594176
rect 343600 594136 371792 594164
rect 343600 594124 343606 594136
rect 371786 594124 371792 594136
rect 371844 594124 371850 594176
rect 288434 594056 288440 594108
rect 288492 594096 288498 594108
rect 345658 594096 345664 594108
rect 288492 594068 345664 594096
rect 288492 594056 288498 594068
rect 345658 594056 345664 594068
rect 345716 594056 345722 594108
rect 371878 594056 371884 594108
rect 371936 594096 371942 594108
rect 391934 594096 391940 594108
rect 371936 594068 391940 594096
rect 371936 594056 371942 594068
rect 391934 594056 391940 594068
rect 391992 594056 391998 594108
rect 254486 593376 254492 593428
rect 254544 593416 254550 593428
rect 275278 593416 275284 593428
rect 254544 593388 275284 593416
rect 254544 593376 254550 593388
rect 275278 593376 275284 593388
rect 275336 593376 275342 593428
rect 311986 592696 311992 592748
rect 312044 592736 312050 592748
rect 322474 592736 322480 592748
rect 312044 592708 322480 592736
rect 312044 592696 312050 592708
rect 322474 592696 322480 592708
rect 322532 592696 322538 592748
rect 254854 592628 254860 592680
rect 254912 592668 254918 592680
rect 269758 592668 269764 592680
rect 254912 592640 269764 592668
rect 254912 592628 254918 592640
rect 269758 592628 269764 592640
rect 269816 592628 269822 592680
rect 293494 592628 293500 592680
rect 293552 592668 293558 592680
rect 347038 592668 347044 592680
rect 293552 592640 347044 592668
rect 293552 592628 293558 592640
rect 347038 592628 347044 592640
rect 347096 592628 347102 592680
rect 385678 592016 385684 592068
rect 385736 592056 385742 592068
rect 389174 592056 389180 592068
rect 385736 592028 389180 592056
rect 385736 592016 385742 592028
rect 389174 592016 389180 592028
rect 389232 592016 389238 592068
rect 306834 591336 306840 591388
rect 306892 591376 306898 591388
rect 334618 591376 334624 591388
rect 306892 591348 334624 591376
rect 306892 591336 306898 591348
rect 334618 591336 334624 591348
rect 334676 591336 334682 591388
rect 336090 591336 336096 591388
rect 336148 591376 336154 591388
rect 396166 591376 396172 591388
rect 336148 591348 396172 591376
rect 336148 591336 336154 591348
rect 396166 591336 396172 591348
rect 396224 591336 396230 591388
rect 260098 591268 260104 591320
rect 260156 591308 260162 591320
rect 480254 591308 480260 591320
rect 260156 591280 480260 591308
rect 260156 591268 260162 591280
rect 480254 591268 480260 591280
rect 480312 591268 480318 591320
rect 478782 590656 478788 590708
rect 478840 590696 478846 590708
rect 579798 590696 579804 590708
rect 478840 590668 579804 590696
rect 478840 590656 478846 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 47854 590588 47860 590640
rect 47912 590628 47918 590640
rect 48958 590628 48964 590640
rect 47912 590600 48964 590628
rect 47912 590588 47918 590600
rect 48958 590588 48964 590600
rect 49016 590588 49022 590640
rect 329742 589976 329748 590028
rect 329800 590016 329806 590028
rect 364702 590016 364708 590028
rect 329800 589988 364708 590016
rect 329800 589976 329806 589988
rect 364702 589976 364708 589988
rect 364760 589976 364766 590028
rect 381538 589976 381544 590028
rect 381596 590016 381602 590028
rect 386414 590016 386420 590028
rect 381596 589988 386420 590016
rect 381596 589976 381602 589988
rect 386414 589976 386420 589988
rect 386472 589976 386478 590028
rect 294598 589908 294604 589960
rect 294656 589948 294662 589960
rect 386782 589948 386788 589960
rect 294656 589920 386788 589948
rect 294656 589908 294662 589920
rect 386782 589908 386788 589920
rect 386840 589908 386846 589960
rect 367186 589432 367192 589484
rect 367244 589472 367250 589484
rect 367370 589472 367376 589484
rect 367244 589444 367376 589472
rect 367244 589432 367250 589444
rect 367370 589432 367376 589444
rect 367428 589432 367434 589484
rect 314838 588616 314844 588668
rect 314896 588656 314902 588668
rect 338850 588656 338856 588668
rect 314896 588628 338856 588656
rect 314896 588616 314902 588628
rect 338850 588616 338856 588628
rect 338908 588616 338914 588668
rect 342162 588616 342168 588668
rect 342220 588656 342226 588668
rect 367186 588656 367192 588668
rect 342220 588628 367192 588656
rect 342220 588616 342226 588628
rect 367186 588616 367192 588628
rect 367244 588616 367250 588668
rect 291378 588548 291384 588600
rect 291436 588588 291442 588600
rect 350074 588588 350080 588600
rect 291436 588560 350080 588588
rect 291436 588548 291442 588560
rect 350074 588548 350080 588560
rect 350132 588548 350138 588600
rect 254578 587936 254584 587988
rect 254636 587976 254642 587988
rect 260098 587976 260104 587988
rect 254636 587948 260104 587976
rect 254636 587936 254642 587948
rect 260098 587936 260104 587948
rect 260156 587936 260162 587988
rect 333882 587188 333888 587240
rect 333940 587228 333946 587240
rect 368566 587228 368572 587240
rect 333940 587200 368572 587228
rect 333940 587188 333946 587200
rect 368566 587188 368572 587200
rect 368624 587188 368630 587240
rect 287974 587120 287980 587172
rect 288032 587160 288038 587172
rect 342898 587160 342904 587172
rect 288032 587132 342904 587160
rect 288032 587120 288038 587132
rect 342898 587120 342904 587132
rect 342956 587120 342962 587172
rect 304718 585828 304724 585880
rect 304776 585868 304782 585880
rect 340138 585868 340144 585880
rect 304776 585840 340144 585868
rect 304776 585828 304782 585840
rect 340138 585828 340144 585840
rect 340196 585828 340202 585880
rect 361114 585828 361120 585880
rect 361172 585868 361178 585880
rect 392118 585868 392124 585880
rect 361172 585840 392124 585868
rect 361172 585828 361178 585840
rect 392118 585828 392124 585840
rect 392176 585828 392182 585880
rect 331950 585760 331956 585812
rect 332008 585800 332014 585812
rect 372798 585800 372804 585812
rect 332008 585772 372804 585800
rect 332008 585760 332014 585772
rect 372798 585760 372804 585772
rect 372856 585760 372862 585812
rect 310606 584400 310612 584452
rect 310664 584440 310670 584452
rect 345750 584440 345756 584452
rect 310664 584412 345756 584440
rect 310664 584400 310670 584412
rect 345750 584400 345756 584412
rect 345808 584400 345814 584452
rect 293954 581612 293960 581664
rect 294012 581652 294018 581664
rect 367186 581652 367192 581664
rect 294012 581624 367192 581652
rect 294012 581612 294018 581624
rect 367186 581612 367192 581624
rect 367244 581612 367250 581664
rect 253934 581272 253940 581324
rect 253992 581312 253998 581324
rect 255958 581312 255964 581324
rect 253992 581284 255964 581312
rect 253992 581272 253998 581284
rect 255958 581272 255964 581284
rect 256016 581272 256022 581324
rect 319438 580252 319444 580304
rect 319496 580292 319502 580304
rect 475562 580292 475568 580304
rect 319496 580264 475568 580292
rect 319496 580252 319502 580264
rect 475562 580252 475568 580264
rect 475620 580252 475626 580304
rect 329098 578892 329104 578944
rect 329156 578932 329162 578944
rect 382458 578932 382464 578944
rect 329156 578904 382464 578932
rect 329156 578892 329162 578904
rect 382458 578892 382464 578904
rect 382516 578892 382522 578944
rect 322382 578144 322388 578196
rect 322440 578184 322446 578196
rect 580166 578184 580172 578196
rect 322440 578156 580172 578184
rect 322440 578144 322446 578156
rect 580166 578144 580172 578156
rect 580224 578144 580230 578196
rect 303430 577532 303436 577584
rect 303488 577572 303494 577584
rect 335998 577572 336004 577584
rect 303488 577544 336004 577572
rect 303488 577532 303494 577544
rect 335998 577532 336004 577544
rect 336056 577532 336062 577584
rect 321186 577464 321192 577516
rect 321244 577504 321250 577516
rect 379514 577504 379520 577516
rect 321244 577476 379520 577504
rect 321244 577464 321250 577476
rect 379514 577464 379520 577476
rect 379572 577464 379578 577516
rect 287054 576172 287060 576224
rect 287112 576212 287118 576224
rect 354214 576212 354220 576224
rect 287112 576184 354220 576212
rect 287112 576172 287118 576184
rect 354214 576172 354220 576184
rect 354272 576172 354278 576224
rect 306466 576104 306472 576156
rect 306524 576144 306530 576156
rect 389266 576144 389272 576156
rect 306524 576116 389272 576144
rect 306524 576104 306530 576116
rect 389266 576104 389272 576116
rect 389324 576104 389330 576156
rect 254210 575492 254216 575544
rect 254268 575532 254274 575544
rect 278038 575532 278044 575544
rect 254268 575504 278044 575532
rect 254268 575492 254274 575504
rect 278038 575492 278044 575504
rect 278096 575492 278102 575544
rect 327810 574812 327816 574864
rect 327868 574852 327874 574864
rect 396166 574852 396172 574864
rect 327868 574824 396172 574852
rect 327868 574812 327874 574824
rect 396166 574812 396172 574824
rect 396224 574812 396230 574864
rect 304810 574744 304816 574796
rect 304868 574784 304874 574796
rect 394878 574784 394884 574796
rect 304868 574756 394884 574784
rect 304868 574744 304874 574756
rect 394878 574744 394884 574756
rect 394936 574744 394942 574796
rect 296714 573384 296720 573436
rect 296772 573424 296778 573436
rect 367370 573424 367376 573436
rect 296772 573396 367376 573424
rect 296772 573384 296778 573396
rect 367370 573384 367376 573396
rect 367428 573384 367434 573436
rect 314746 573316 314752 573368
rect 314804 573356 314810 573368
rect 390646 573356 390652 573368
rect 314804 573328 390652 573356
rect 314804 573316 314810 573328
rect 390646 573316 390652 573328
rect 390704 573316 390710 573368
rect 285674 572024 285680 572076
rect 285732 572064 285738 572076
rect 353110 572064 353116 572076
rect 285732 572036 353116 572064
rect 285732 572024 285738 572036
rect 353110 572024 353116 572036
rect 353168 572024 353174 572076
rect 319530 571956 319536 572008
rect 319588 571996 319594 572008
rect 522114 571996 522120 572008
rect 319588 571968 522120 571996
rect 319588 571956 319594 571968
rect 522114 571956 522120 571968
rect 522172 571956 522178 572008
rect 310514 570664 310520 570716
rect 310572 570704 310578 570716
rect 374270 570704 374276 570716
rect 310572 570676 374276 570704
rect 310572 570664 310578 570676
rect 374270 570664 374276 570676
rect 374328 570664 374334 570716
rect 284386 570596 284392 570648
rect 284444 570636 284450 570648
rect 386598 570636 386604 570648
rect 284444 570608 386604 570636
rect 284444 570596 284450 570608
rect 386598 570596 386604 570608
rect 386656 570596 386662 570648
rect 253934 569984 253940 570036
rect 253992 570024 253998 570036
rect 256050 570024 256056 570036
rect 253992 569996 256056 570024
rect 253992 569984 253998 569996
rect 256050 569984 256056 569996
rect 256108 569984 256114 570036
rect 292574 569168 292580 569220
rect 292632 569208 292638 569220
rect 357066 569208 357072 569220
rect 292632 569180 357072 569208
rect 292632 569168 292638 569180
rect 357066 569168 357072 569180
rect 357124 569168 357130 569220
rect 307754 567876 307760 567928
rect 307812 567916 307818 567928
rect 368566 567916 368572 567928
rect 307812 567888 368572 567916
rect 307812 567876 307818 567888
rect 368566 567876 368572 567888
rect 368624 567876 368630 567928
rect 289078 567808 289084 567860
rect 289136 567848 289142 567860
rect 386690 567848 386696 567860
rect 289136 567820 386696 567848
rect 289136 567808 289142 567820
rect 386690 567808 386696 567820
rect 386748 567808 386754 567860
rect 388530 567196 388536 567248
rect 388588 567236 388594 567248
rect 393406 567236 393412 567248
rect 388588 567208 393412 567236
rect 388588 567196 388594 567208
rect 393406 567196 393412 567208
rect 393464 567196 393470 567248
rect 3326 567128 3332 567180
rect 3384 567168 3390 567180
rect 50430 567168 50436 567180
rect 3384 567140 50436 567168
rect 3384 567128 3390 567140
rect 50430 567128 50436 567140
rect 50488 567128 50494 567180
rect 313366 566448 313372 566500
rect 313424 566488 313430 566500
rect 376846 566488 376852 566500
rect 313424 566460 376852 566488
rect 313424 566448 313430 566460
rect 376846 566448 376852 566460
rect 376904 566448 376910 566500
rect 372706 565836 372712 565888
rect 372764 565876 372770 565888
rect 404906 565876 404912 565888
rect 372764 565848 404912 565876
rect 372764 565836 372770 565848
rect 404906 565836 404912 565848
rect 404964 565836 404970 565888
rect 350442 565224 350448 565276
rect 350500 565264 350506 565276
rect 372706 565264 372712 565276
rect 350500 565236 372712 565264
rect 350500 565224 350506 565236
rect 372706 565224 372712 565236
rect 372764 565224 372770 565276
rect 306190 565156 306196 565208
rect 306248 565196 306254 565208
rect 365898 565196 365904 565208
rect 306248 565168 365904 565196
rect 306248 565156 306254 565168
rect 365898 565156 365904 565168
rect 365956 565156 365962 565208
rect 283006 565088 283012 565140
rect 283064 565128 283070 565140
rect 354306 565128 354312 565140
rect 283064 565100 354312 565128
rect 283064 565088 283070 565100
rect 354306 565088 354312 565100
rect 354364 565088 354370 565140
rect 358262 565088 358268 565140
rect 358320 565128 358326 565140
rect 396074 565128 396080 565140
rect 358320 565100 396080 565128
rect 358320 565088 358326 565100
rect 396074 565088 396080 565100
rect 396132 565088 396138 565140
rect 254578 564408 254584 564460
rect 254636 564448 254642 564460
rect 279418 564448 279424 564460
rect 254636 564420 279424 564448
rect 254636 564408 254642 564420
rect 279418 564408 279424 564420
rect 279476 564408 279482 564460
rect 359090 563796 359096 563848
rect 359148 563836 359154 563848
rect 386506 563836 386512 563848
rect 359148 563808 386512 563836
rect 359148 563796 359154 563808
rect 386506 563796 386512 563808
rect 386564 563796 386570 563848
rect 358354 563728 358360 563780
rect 358412 563768 358418 563780
rect 394694 563768 394700 563780
rect 358412 563740 394700 563768
rect 358412 563728 358418 563740
rect 394694 563728 394700 563740
rect 394752 563728 394758 563780
rect 300762 563660 300768 563712
rect 300820 563700 300826 563712
rect 362954 563700 362960 563712
rect 300820 563672 362960 563700
rect 300820 563660 300826 563672
rect 362954 563660 362960 563672
rect 363012 563660 363018 563712
rect 321094 562368 321100 562420
rect 321152 562408 321158 562420
rect 401962 562408 401968 562420
rect 321152 562380 401968 562408
rect 321152 562368 321158 562380
rect 401962 562368 401968 562380
rect 402020 562368 402026 562420
rect 253198 562300 253204 562352
rect 253256 562340 253262 562352
rect 381078 562340 381084 562352
rect 253256 562312 381084 562340
rect 253256 562300 253262 562312
rect 381078 562300 381084 562312
rect 381136 562300 381142 562352
rect 321002 560940 321008 560992
rect 321060 560980 321066 560992
rect 402054 560980 402060 560992
rect 321060 560952 402060 560980
rect 321060 560940 321066 560952
rect 402054 560940 402060 560952
rect 402112 560940 402118 560992
rect 384298 560736 384304 560788
rect 384356 560776 384362 560788
rect 390738 560776 390744 560788
rect 384356 560748 390744 560776
rect 384356 560736 384362 560748
rect 390738 560736 390744 560748
rect 390796 560736 390802 560788
rect 363230 559648 363236 559700
rect 363288 559688 363294 559700
rect 374086 559688 374092 559700
rect 363288 559660 374092 559688
rect 363288 559648 363294 559660
rect 374086 559648 374092 559660
rect 374144 559648 374150 559700
rect 364426 559580 364432 559632
rect 364484 559620 364490 559632
rect 376662 559620 376668 559632
rect 364484 559592 376668 559620
rect 364484 559580 364490 559592
rect 376662 559580 376668 559592
rect 376720 559620 376726 559632
rect 396074 559620 396080 559632
rect 376720 559592 396080 559620
rect 376720 559580 376726 559592
rect 396074 559580 396080 559592
rect 396132 559580 396138 559632
rect 316126 559512 316132 559564
rect 316184 559552 316190 559564
rect 400950 559552 400956 559564
rect 316184 559524 400956 559552
rect 316184 559512 316190 559524
rect 400950 559512 400956 559524
rect 401008 559512 401014 559564
rect 358998 558220 359004 558272
rect 359056 558260 359062 558272
rect 380986 558260 380992 558272
rect 359056 558232 380992 558260
rect 359056 558220 359062 558232
rect 380986 558220 380992 558232
rect 381044 558220 381050 558272
rect 291838 558152 291844 558204
rect 291896 558192 291902 558204
rect 375466 558192 375472 558204
rect 291896 558164 375472 558192
rect 291896 558152 291902 558164
rect 375466 558152 375472 558164
rect 375524 558152 375530 558204
rect 376754 558152 376760 558204
rect 376812 558192 376818 558204
rect 377122 558192 377128 558204
rect 376812 558164 377128 558192
rect 376812 558152 376818 558164
rect 377122 558152 377128 558164
rect 377180 558152 377186 558204
rect 254578 557540 254584 557592
rect 254636 557580 254642 557592
rect 265618 557580 265624 557592
rect 254636 557552 265624 557580
rect 254636 557540 254642 557552
rect 265618 557540 265624 557552
rect 265676 557540 265682 557592
rect 357894 556860 357900 556912
rect 357952 556900 357958 556912
rect 381170 556900 381176 556912
rect 357952 556872 381176 556900
rect 357952 556860 357958 556872
rect 381170 556860 381176 556872
rect 381228 556860 381234 556912
rect 362586 556792 362592 556844
rect 362644 556832 362650 556844
rect 373994 556832 374000 556844
rect 362644 556804 374000 556832
rect 362644 556792 362650 556804
rect 373994 556792 374000 556804
rect 374052 556792 374058 556844
rect 378042 556792 378048 556844
rect 378100 556832 378106 556844
rect 538858 556832 538864 556844
rect 378100 556804 538864 556832
rect 378100 556792 378106 556804
rect 538858 556792 538864 556804
rect 538916 556792 538922 556844
rect 365806 556180 365812 556232
rect 365864 556220 365870 556232
rect 371326 556220 371332 556232
rect 365864 556192 371332 556220
rect 365864 556180 365870 556192
rect 371326 556180 371332 556192
rect 371384 556180 371390 556232
rect 359182 555500 359188 555552
rect 359240 555540 359246 555552
rect 385126 555540 385132 555552
rect 359240 555512 385132 555540
rect 359240 555500 359246 555512
rect 385126 555500 385132 555512
rect 385184 555500 385190 555552
rect 284294 555432 284300 555484
rect 284352 555472 284358 555484
rect 399846 555472 399852 555484
rect 284352 555444 399852 555472
rect 284352 555432 284358 555444
rect 399846 555432 399852 555444
rect 399904 555432 399910 555484
rect 369946 554820 369952 554872
rect 370004 554860 370010 554872
rect 402974 554860 402980 554872
rect 370004 554832 402980 554860
rect 370004 554820 370010 554832
rect 402974 554820 402980 554832
rect 403032 554820 403038 554872
rect 367094 554752 367100 554804
rect 367152 554792 367158 554804
rect 404538 554792 404544 554804
rect 367152 554764 404544 554792
rect 367152 554752 367158 554764
rect 404538 554752 404544 554764
rect 404596 554752 404602 554804
rect 2958 554684 2964 554736
rect 3016 554724 3022 554736
rect 50338 554724 50344 554736
rect 3016 554696 50344 554724
rect 3016 554684 3022 554696
rect 50338 554684 50344 554696
rect 50396 554684 50402 554736
rect 355594 554208 355600 554260
rect 355652 554248 355658 554260
rect 367094 554248 367100 554260
rect 355652 554220 367100 554248
rect 355652 554208 355658 554220
rect 367094 554208 367100 554220
rect 367152 554208 367158 554260
rect 355778 554140 355784 554192
rect 355836 554180 355842 554192
rect 369946 554180 369952 554192
rect 355836 554152 369952 554180
rect 355836 554140 355842 554152
rect 369946 554140 369952 554152
rect 370004 554140 370010 554192
rect 322290 554072 322296 554124
rect 322348 554112 322354 554124
rect 401870 554112 401876 554124
rect 322348 554084 401876 554112
rect 322348 554072 322354 554084
rect 401870 554072 401876 554084
rect 401928 554072 401934 554124
rect 314654 554004 314660 554056
rect 314712 554044 314718 554056
rect 401226 554044 401232 554056
rect 314712 554016 401232 554044
rect 314712 554004 314718 554016
rect 401226 554004 401232 554016
rect 401284 554004 401290 554056
rect 392578 553324 392584 553376
rect 392636 553364 392642 553376
rect 394142 553364 394148 553376
rect 392636 553336 394148 553364
rect 392636 553324 392642 553336
rect 394142 553324 394148 553336
rect 394200 553324 394206 553376
rect 385034 553256 385040 553308
rect 385092 553296 385098 553308
rect 392210 553296 392216 553308
rect 385092 553268 392216 553296
rect 385092 553256 385098 553268
rect 392210 553256 392216 553268
rect 392268 553256 392274 553308
rect 389266 553052 389272 553104
rect 389324 553092 389330 553104
rect 399110 553092 399116 553104
rect 389324 553064 399116 553092
rect 389324 553052 389330 553064
rect 399110 553052 399116 553064
rect 399168 553052 399174 553104
rect 360102 552916 360108 552968
rect 360160 552956 360166 552968
rect 378686 552956 378692 552968
rect 360160 552928 378692 552956
rect 360160 552916 360166 552928
rect 378686 552916 378692 552928
rect 378744 552916 378750 552968
rect 383746 552916 383752 552968
rect 383804 552956 383810 552968
rect 400030 552956 400036 552968
rect 383804 552928 400036 552956
rect 383804 552916 383810 552928
rect 400030 552916 400036 552928
rect 400088 552916 400094 552968
rect 368658 552888 368664 552900
rect 354646 552860 368664 552888
rect 347130 552780 347136 552832
rect 347188 552820 347194 552832
rect 354646 552820 354674 552860
rect 368658 552848 368664 552860
rect 368716 552888 368722 552900
rect 388346 552888 388352 552900
rect 368716 552860 388352 552888
rect 368716 552848 368722 552860
rect 388346 552848 388352 552860
rect 388404 552848 388410 552900
rect 347188 552792 354674 552820
rect 347188 552780 347194 552792
rect 379974 552780 379980 552832
rect 380032 552820 380038 552832
rect 400398 552820 400404 552832
rect 380032 552792 400404 552820
rect 380032 552780 380038 552792
rect 400398 552780 400404 552792
rect 400456 552780 400462 552832
rect 356698 552712 356704 552764
rect 356756 552752 356762 552764
rect 396718 552752 396724 552764
rect 356756 552724 396724 552752
rect 356756 552712 356762 552724
rect 396718 552712 396724 552724
rect 396776 552712 396782 552764
rect 309226 552644 309232 552696
rect 309284 552684 309290 552696
rect 360654 552684 360660 552696
rect 309284 552656 360660 552684
rect 309284 552644 309290 552656
rect 360654 552644 360660 552656
rect 360712 552644 360718 552696
rect 361482 552644 361488 552696
rect 361540 552684 361546 552696
rect 374178 552684 374184 552696
rect 361540 552656 374184 552684
rect 361540 552644 361546 552656
rect 374178 552644 374184 552656
rect 374236 552644 374242 552696
rect 376110 552644 376116 552696
rect 376168 552684 376174 552696
rect 399018 552684 399024 552696
rect 376168 552656 399024 552684
rect 376168 552644 376174 552656
rect 399018 552644 399024 552656
rect 399076 552644 399082 552696
rect 399478 552644 399484 552696
rect 399536 552684 399542 552696
rect 402422 552684 402428 552696
rect 399536 552656 402428 552684
rect 399536 552644 399542 552656
rect 402422 552644 402428 552656
rect 402480 552644 402486 552696
rect 393498 552508 393504 552560
rect 393556 552548 393562 552560
rect 400490 552548 400496 552560
rect 393556 552520 400496 552548
rect 393556 552508 393562 552520
rect 400490 552508 400496 552520
rect 400548 552508 400554 552560
rect 355226 552304 355232 552356
rect 355284 552344 355290 552356
rect 361114 552344 361120 552356
rect 355284 552316 361120 552344
rect 355284 552304 355290 552316
rect 361114 552304 361120 552316
rect 361172 552304 361178 552356
rect 375650 552304 375656 552356
rect 375708 552344 375714 552356
rect 403434 552344 403440 552356
rect 375708 552316 403440 552344
rect 375708 552304 375714 552316
rect 403434 552304 403440 552316
rect 403492 552304 403498 552356
rect 356606 552236 356612 552288
rect 356664 552276 356670 552288
rect 385678 552276 385684 552288
rect 356664 552248 385684 552276
rect 356664 552236 356670 552248
rect 385678 552236 385684 552248
rect 385736 552236 385742 552288
rect 398650 552236 398656 552288
rect 398708 552276 398714 552288
rect 409138 552276 409144 552288
rect 398708 552248 409144 552276
rect 398708 552236 398714 552248
rect 409138 552236 409144 552248
rect 409196 552236 409202 552288
rect 354398 552168 354404 552220
rect 354456 552208 354462 552220
rect 384298 552208 384304 552220
rect 354456 552180 384304 552208
rect 354456 552168 354462 552180
rect 384298 552168 384304 552180
rect 384356 552168 384362 552220
rect 394786 552168 394792 552220
rect 394844 552208 394850 552220
rect 430574 552208 430580 552220
rect 394844 552180 430580 552208
rect 394844 552168 394850 552180
rect 430574 552168 430580 552180
rect 430632 552168 430638 552220
rect 357158 552100 357164 552152
rect 357216 552140 357222 552152
rect 371878 552140 371884 552152
rect 357216 552112 371884 552140
rect 357216 552100 357222 552112
rect 371878 552100 371884 552112
rect 371936 552100 371942 552152
rect 373534 552100 373540 552152
rect 373592 552140 373598 552152
rect 498838 552140 498844 552152
rect 373592 552112 498844 552140
rect 373592 552100 373598 552112
rect 498838 552100 498844 552112
rect 498896 552100 498902 552152
rect 254578 552032 254584 552084
rect 254636 552072 254642 552084
rect 268378 552072 268384 552084
rect 254636 552044 268384 552072
rect 254636 552032 254642 552044
rect 268378 552032 268384 552044
rect 268436 552032 268442 552084
rect 348418 552032 348424 552084
rect 348476 552072 348482 552084
rect 381538 552072 381544 552084
rect 348476 552044 381544 552072
rect 348476 552032 348482 552044
rect 381538 552032 381544 552044
rect 381596 552032 381602 552084
rect 391198 552032 391204 552084
rect 391256 552072 391262 552084
rect 391566 552072 391572 552084
rect 391256 552044 391572 552072
rect 391256 552032 391262 552044
rect 391566 552032 391572 552044
rect 391624 552072 391630 552084
rect 520550 552072 520556 552084
rect 391624 552044 520556 552072
rect 391624 552032 391630 552044
rect 520550 552032 520556 552044
rect 520608 552032 520614 552084
rect 398098 551964 398104 552016
rect 398156 552004 398162 552016
rect 401594 552004 401600 552016
rect 398156 551976 401600 552004
rect 398156 551964 398162 551976
rect 401594 551964 401600 551976
rect 401652 551964 401658 552016
rect 375006 551896 375012 551948
rect 375064 551936 375070 551948
rect 375650 551936 375656 551948
rect 375064 551908 375656 551936
rect 375064 551896 375070 551908
rect 375650 551896 375656 551908
rect 375708 551896 375714 551948
rect 358078 551692 358084 551744
rect 358136 551732 358142 551744
rect 360930 551732 360936 551744
rect 358136 551704 360936 551732
rect 358136 551692 358142 551704
rect 360930 551692 360936 551704
rect 360988 551692 360994 551744
rect 389450 551692 389456 551744
rect 389508 551732 389514 551744
rect 399754 551732 399760 551744
rect 389508 551704 399760 551732
rect 389508 551692 389514 551704
rect 399754 551692 399760 551704
rect 399812 551692 399818 551744
rect 355134 551624 355140 551676
rect 355192 551664 355198 551676
rect 377122 551664 377128 551676
rect 355192 551636 377128 551664
rect 355192 551624 355198 551636
rect 377122 551624 377128 551636
rect 377180 551664 377186 551676
rect 400766 551664 400772 551676
rect 377180 551636 400772 551664
rect 377180 551624 377186 551636
rect 400766 551624 400772 551636
rect 400824 551624 400830 551676
rect 322382 551556 322388 551608
rect 322440 551596 322446 551608
rect 376662 551596 376668 551608
rect 322440 551568 376668 551596
rect 322440 551556 322446 551568
rect 376662 551556 376668 551568
rect 376720 551556 376726 551608
rect 383654 551556 383660 551608
rect 383712 551596 383718 551608
rect 399478 551596 399484 551608
rect 383712 551568 399484 551596
rect 383712 551556 383718 551568
rect 399478 551556 399484 551568
rect 399536 551556 399542 551608
rect 304626 551488 304632 551540
rect 304684 551528 304690 551540
rect 403066 551528 403072 551540
rect 304684 551500 403072 551528
rect 304684 551488 304690 551500
rect 403066 551488 403072 551500
rect 403124 551488 403130 551540
rect 295518 551420 295524 551472
rect 295576 551460 295582 551472
rect 403342 551460 403348 551472
rect 295576 551432 403348 551460
rect 295576 551420 295582 551432
rect 403342 551420 403348 551432
rect 403400 551420 403406 551472
rect 295334 551352 295340 551404
rect 295392 551392 295398 551404
rect 403526 551392 403532 551404
rect 295392 551364 403532 551392
rect 295392 551352 295398 551364
rect 403526 551352 403532 551364
rect 403584 551352 403590 551404
rect 295426 551284 295432 551336
rect 295484 551324 295490 551336
rect 404446 551324 404452 551336
rect 295484 551296 404452 551324
rect 295484 551284 295490 551296
rect 404446 551284 404452 551296
rect 404504 551284 404510 551336
rect 358170 551216 358176 551268
rect 358228 551256 358234 551268
rect 361022 551256 361028 551268
rect 358228 551228 361028 551256
rect 358228 551216 358234 551228
rect 361022 551216 361028 551228
rect 361080 551216 361086 551268
rect 363138 551216 363144 551268
rect 363196 551256 363202 551268
rect 363598 551256 363604 551268
rect 363196 551228 363604 551256
rect 363196 551216 363202 551228
rect 363598 551216 363604 551228
rect 363656 551216 363662 551268
rect 382274 551216 382280 551268
rect 382332 551256 382338 551268
rect 382918 551256 382924 551268
rect 382332 551228 382924 551256
rect 382332 551216 382338 551228
rect 382918 551216 382924 551228
rect 382976 551216 382982 551268
rect 364334 551080 364340 551132
rect 364392 551120 364398 551132
rect 365162 551120 365168 551132
rect 364392 551092 365168 551120
rect 364392 551080 364398 551092
rect 365162 551080 365168 551092
rect 365220 551080 365226 551132
rect 351270 550808 351276 550860
rect 351328 550848 351334 550860
rect 388530 550848 388536 550860
rect 351328 550820 388536 550848
rect 351328 550808 351334 550820
rect 388530 550808 388536 550820
rect 388588 550848 388594 550860
rect 388990 550848 388996 550860
rect 388588 550820 388996 550848
rect 388588 550808 388594 550820
rect 388990 550808 388996 550820
rect 389048 550808 389054 550860
rect 358722 550740 358728 550792
rect 358780 550780 358786 550792
rect 360838 550780 360844 550792
rect 358780 550752 360844 550780
rect 358780 550740 358786 550752
rect 360838 550740 360844 550752
rect 360896 550740 360902 550792
rect 367094 550740 367100 550792
rect 367152 550780 367158 550792
rect 419534 550780 419540 550792
rect 367152 550752 419540 550780
rect 367152 550740 367158 550752
rect 419534 550740 419540 550752
rect 419592 550740 419598 550792
rect 341610 550672 341616 550724
rect 341668 550712 341674 550724
rect 342162 550712 342168 550724
rect 341668 550684 342168 550712
rect 341668 550672 341674 550684
rect 342162 550672 342168 550684
rect 342220 550712 342226 550724
rect 404354 550712 404360 550724
rect 342220 550684 404360 550712
rect 342220 550672 342226 550684
rect 404354 550672 404360 550684
rect 404412 550672 404418 550724
rect 351178 550604 351184 550656
rect 351236 550644 351242 550656
rect 364334 550644 364340 550656
rect 351236 550616 364340 550644
rect 351236 550604 351242 550616
rect 364334 550604 364340 550616
rect 364392 550604 364398 550656
rect 369026 550604 369032 550656
rect 369084 550644 369090 550656
rect 448514 550644 448520 550656
rect 369084 550616 448520 550644
rect 369084 550604 369090 550616
rect 448514 550604 448520 550616
rect 448572 550604 448578 550656
rect 386598 550536 386604 550588
rect 386656 550576 386662 550588
rect 387058 550576 387064 550588
rect 386656 550548 387064 550576
rect 386656 550536 386662 550548
rect 387058 550536 387064 550548
rect 387116 550536 387122 550588
rect 399662 550536 399668 550588
rect 399720 550576 399726 550588
rect 401686 550576 401692 550588
rect 399720 550548 401692 550576
rect 399720 550536 399726 550548
rect 401686 550536 401692 550548
rect 401744 550536 401750 550588
rect 393314 550468 393320 550520
rect 393372 550508 393378 550520
rect 400490 550508 400496 550520
rect 393372 550480 400496 550508
rect 393372 550468 393378 550480
rect 400490 550468 400496 550480
rect 400548 550468 400554 550520
rect 375346 550140 385034 550168
rect 375006 550100 375012 550112
rect 354646 550072 375012 550100
rect 353202 549992 353208 550044
rect 353260 550032 353266 550044
rect 354646 550032 354674 550072
rect 375006 550060 375012 550072
rect 375064 550060 375070 550112
rect 353260 550004 354674 550032
rect 353260 549992 353266 550004
rect 355870 549992 355876 550044
rect 355928 550032 355934 550044
rect 362954 550032 362960 550044
rect 355928 550004 362960 550032
rect 355928 549992 355934 550004
rect 362954 549992 362960 550004
rect 363012 549992 363018 550044
rect 355686 549924 355692 549976
rect 355744 549964 355750 549976
rect 375346 549964 375374 550140
rect 380158 550060 380164 550112
rect 380216 550100 380222 550112
rect 383930 550100 383936 550112
rect 380216 550072 383936 550100
rect 380216 550060 380222 550072
rect 383930 550060 383936 550072
rect 383988 550060 383994 550112
rect 355744 549936 375374 549964
rect 355744 549924 355750 549936
rect 378778 549924 378784 549976
rect 378836 549964 378842 549976
rect 380986 549964 380992 549976
rect 378836 549936 380992 549964
rect 378836 549924 378842 549936
rect 380986 549924 380992 549936
rect 381044 549924 381050 549976
rect 385006 549964 385034 550140
rect 397638 550100 397644 550112
rect 393286 550072 397644 550100
rect 393286 549964 393314 550072
rect 397638 550060 397644 550072
rect 397696 550060 397702 550112
rect 397546 549992 397552 550044
rect 397604 549992 397610 550044
rect 385006 549936 393314 549964
rect 352374 549856 352380 549908
rect 352432 549896 352438 549908
rect 380158 549896 380164 549908
rect 352432 549868 380164 549896
rect 352432 549856 352438 549868
rect 380158 549856 380164 549868
rect 380216 549856 380222 549908
rect 383562 549896 383568 549908
rect 380820 549868 383568 549896
rect 359918 549788 359924 549840
rect 359976 549828 359982 549840
rect 362310 549828 362316 549840
rect 359976 549800 362316 549828
rect 359976 549788 359982 549800
rect 362310 549788 362316 549800
rect 362368 549788 362374 549840
rect 371326 549828 371332 549840
rect 369826 549800 371332 549828
rect 359826 549652 359832 549704
rect 359884 549692 359890 549704
rect 359884 549664 367094 549692
rect 359884 549652 359890 549664
rect 367066 549624 367094 549664
rect 369826 549624 369854 549800
rect 371326 549788 371332 549800
rect 371384 549788 371390 549840
rect 378778 549828 378784 549840
rect 373966 549800 378784 549828
rect 373966 549624 373994 549800
rect 378778 549788 378784 549800
rect 378836 549788 378842 549840
rect 354646 549596 365116 549624
rect 367066 549596 369854 549624
rect 371896 549596 373994 549624
rect 352466 549516 352472 549568
rect 352524 549556 352530 549568
rect 354646 549556 354674 549596
rect 352524 549528 354674 549556
rect 365088 549556 365116 549596
rect 371896 549556 371924 549596
rect 365088 549528 371924 549556
rect 352524 549516 352530 549528
rect 324222 549380 324228 549432
rect 324280 549420 324286 549432
rect 359918 549420 359924 549432
rect 324280 549392 359924 549420
rect 324280 549380 324286 549392
rect 359918 549380 359924 549392
rect 359976 549380 359982 549432
rect 327810 549312 327816 549364
rect 327868 549352 327874 549364
rect 359826 549352 359832 549364
rect 327868 549324 359832 549352
rect 327868 549312 327874 549324
rect 359826 549312 359832 549324
rect 359884 549312 359890 549364
rect 325510 549244 325516 549296
rect 325568 549284 325574 549296
rect 380820 549284 380848 549868
rect 383562 549856 383568 549868
rect 383620 549856 383626 549908
rect 383930 549856 383936 549908
rect 383988 549896 383994 549908
rect 397564 549896 397592 549992
rect 400674 549896 400680 549908
rect 383988 549868 400680 549896
rect 383988 549856 383994 549868
rect 400674 549856 400680 549868
rect 400732 549856 400738 549908
rect 380986 549788 380992 549840
rect 381044 549788 381050 549840
rect 383626 549800 383884 549828
rect 381004 549692 381032 549788
rect 383626 549692 383654 549800
rect 383856 549760 383884 549800
rect 383856 549732 385034 549760
rect 381004 549664 383654 549692
rect 385006 549556 385034 549732
rect 400582 549720 400588 549772
rect 400640 549760 400646 549772
rect 401042 549760 401048 549772
rect 400640 549732 401048 549760
rect 400640 549720 400646 549732
rect 401042 549720 401048 549732
rect 401100 549720 401106 549772
rect 400582 549556 400588 549568
rect 385006 549528 400588 549556
rect 400582 549516 400588 549528
rect 400640 549516 400646 549568
rect 325568 549256 380848 549284
rect 325568 549244 325574 549256
rect 322290 548564 322296 548616
rect 322348 548604 322354 548616
rect 356606 548604 356612 548616
rect 322348 548576 356612 548604
rect 322348 548564 322354 548576
rect 356606 548564 356612 548576
rect 356664 548564 356670 548616
rect 302142 548496 302148 548548
rect 302200 548536 302206 548548
rect 357066 548536 357072 548548
rect 302200 548508 357072 548536
rect 302200 548496 302206 548508
rect 357066 548496 357072 548508
rect 357124 548496 357130 548548
rect 281534 547816 281540 547868
rect 281592 547856 281598 547868
rect 357434 547856 357440 547868
rect 281592 547828 357440 547856
rect 281592 547816 281598 547828
rect 357434 547816 357440 547828
rect 357492 547816 357498 547868
rect 254578 546456 254584 546508
rect 254636 546496 254642 546508
rect 261478 546496 261484 546508
rect 254636 546468 261484 546496
rect 254636 546456 254642 546468
rect 261478 546456 261484 546468
rect 261536 546456 261542 546508
rect 399570 546456 399576 546508
rect 399628 546496 399634 546508
rect 402514 546496 402520 546508
rect 399628 546468 402520 546496
rect 399628 546456 399634 546468
rect 402514 546456 402520 546468
rect 402572 546456 402578 546508
rect 322474 546388 322480 546440
rect 322532 546428 322538 546440
rect 357434 546428 357440 546440
rect 322532 546400 357440 546428
rect 322532 546388 322538 546400
rect 357434 546388 357440 546400
rect 357492 546388 357498 546440
rect 276842 545844 276848 545896
rect 276900 545884 276906 545896
rect 301866 545884 301872 545896
rect 276900 545856 301872 545884
rect 276900 545844 276906 545856
rect 301866 545844 301872 545856
rect 301924 545844 301930 545896
rect 279694 545776 279700 545828
rect 279752 545816 279758 545828
rect 312906 545816 312912 545828
rect 279752 545788 312912 545816
rect 279752 545776 279758 545788
rect 312906 545776 312912 545788
rect 312964 545776 312970 545828
rect 279602 545708 279608 545760
rect 279660 545748 279666 545760
rect 313642 545748 313648 545760
rect 279660 545720 313648 545748
rect 279660 545708 279666 545720
rect 313642 545708 313648 545720
rect 313700 545708 313706 545760
rect 317414 545708 317420 545760
rect 317472 545748 317478 545760
rect 332594 545748 332600 545760
rect 317472 545720 332600 545748
rect 317472 545708 317478 545720
rect 332594 545708 332600 545720
rect 332652 545708 332658 545760
rect 254670 545028 254676 545080
rect 254728 545068 254734 545080
rect 260190 545068 260196 545080
rect 254728 545040 260196 545068
rect 254728 545028 254734 545040
rect 260190 545028 260196 545040
rect 260248 545028 260254 545080
rect 306374 545028 306380 545080
rect 306432 545068 306438 545080
rect 357434 545068 357440 545080
rect 306432 545040 357440 545068
rect 306432 545028 306438 545040
rect 357434 545028 357440 545040
rect 357492 545028 357498 545080
rect 309134 544348 309140 544400
rect 309192 544388 309198 544400
rect 355502 544388 355508 544400
rect 309192 544360 355508 544388
rect 309192 544348 309198 544360
rect 355502 544348 355508 544360
rect 355560 544348 355566 544400
rect 482186 544348 482192 544400
rect 482244 544388 482250 544400
rect 525058 544388 525064 544400
rect 482244 544360 525064 544388
rect 482244 544348 482250 544360
rect 525058 544348 525064 544360
rect 525116 544348 525122 544400
rect 357618 543736 357624 543788
rect 357676 543776 357682 543788
rect 359642 543776 359648 543788
rect 357676 543748 359648 543776
rect 357676 543736 357682 543748
rect 359642 543736 359648 543748
rect 359700 543736 359706 543788
rect 279878 543668 279884 543720
rect 279936 543708 279942 543720
rect 298186 543708 298192 543720
rect 279936 543680 298192 543708
rect 279936 543668 279942 543680
rect 298186 543668 298192 543680
rect 298244 543668 298250 543720
rect 279326 543532 279332 543584
rect 279384 543572 279390 543584
rect 298922 543572 298928 543584
rect 279384 543544 298928 543572
rect 279384 543532 279390 543544
rect 298922 543532 298928 543544
rect 298980 543532 298986 543584
rect 401778 543532 401784 543584
rect 401836 543572 401842 543584
rect 402054 543572 402060 543584
rect 401836 543544 402060 543572
rect 401836 543532 401842 543544
rect 402054 543532 402060 543544
rect 402112 543532 402118 543584
rect 478966 543532 478972 543584
rect 479024 543572 479030 543584
rect 479702 543572 479708 543584
rect 479024 543544 479708 543572
rect 479024 543532 479030 543544
rect 479702 543532 479708 543544
rect 479760 543532 479766 543584
rect 279234 543464 279240 543516
rect 279292 543504 279298 543516
rect 299658 543504 299664 543516
rect 279292 543476 299664 543504
rect 279292 543464 279298 543476
rect 299658 543464 299664 543476
rect 299716 543464 299722 543516
rect 279510 543396 279516 543448
rect 279568 543436 279574 543448
rect 302602 543436 302608 543448
rect 279568 543408 302608 543436
rect 279568 543396 279574 543408
rect 302602 543396 302608 543408
rect 302660 543396 302666 543448
rect 401778 543396 401784 543448
rect 401836 543436 401842 543448
rect 404538 543436 404544 543448
rect 401836 543408 404544 543436
rect 401836 543396 401842 543408
rect 404538 543396 404544 543408
rect 404596 543396 404602 543448
rect 276750 543328 276756 543380
rect 276808 543368 276814 543380
rect 304074 543368 304080 543380
rect 276808 543340 304080 543368
rect 276808 543328 276814 543340
rect 304074 543328 304080 543340
rect 304132 543328 304138 543380
rect 279142 543260 279148 543312
rect 279200 543300 279206 543312
rect 316310 543300 316316 543312
rect 279200 543272 316316 543300
rect 279200 543260 279206 543272
rect 316310 543260 316316 543272
rect 316368 543260 316374 543312
rect 280062 543192 280068 543244
rect 280120 543232 280126 543244
rect 315114 543232 315120 543244
rect 280120 543204 315120 543232
rect 280120 543192 280126 543204
rect 315114 543192 315120 543204
rect 315172 543192 315178 543244
rect 278130 543124 278136 543176
rect 278188 543164 278194 543176
rect 316586 543164 316592 543176
rect 278188 543136 316592 543164
rect 278188 543124 278194 543136
rect 316586 543124 316592 543136
rect 316644 543124 316650 543176
rect 427814 543124 427820 543176
rect 427872 543164 427878 543176
rect 509418 543164 509424 543176
rect 427872 543136 509424 543164
rect 427872 543124 427878 543136
rect 509418 543124 509424 543136
rect 509476 543124 509482 543176
rect 276658 543056 276664 543108
rect 276716 543096 276722 543108
rect 303614 543096 303620 543108
rect 276716 543068 303620 543096
rect 276716 543056 276722 543068
rect 303614 543056 303620 543068
rect 303672 543056 303678 543108
rect 326338 543056 326344 543108
rect 326396 543096 326402 543108
rect 357710 543096 357716 543108
rect 326396 543068 357716 543096
rect 326396 543056 326402 543068
rect 357710 543056 357716 543068
rect 357768 543056 357774 543108
rect 420914 543056 420920 543108
rect 420972 543096 420978 543108
rect 513374 543096 513380 543108
rect 420972 543068 513380 543096
rect 420972 543056 420978 543068
rect 513374 543056 513380 543068
rect 513432 543056 513438 543108
rect 279970 542988 279976 543040
rect 280028 543028 280034 543040
rect 314838 543028 314844 543040
rect 280028 543000 314844 543028
rect 280028 542988 280034 543000
rect 314838 542988 314844 543000
rect 314896 542988 314902 543040
rect 316034 542988 316040 543040
rect 316092 543028 316098 543040
rect 354122 543028 354128 543040
rect 316092 543000 354128 543028
rect 316092 542988 316098 543000
rect 354122 542988 354128 543000
rect 354180 542988 354186 543040
rect 416774 542988 416780 543040
rect 416832 543028 416838 543040
rect 482278 543028 482284 543040
rect 416832 543000 482284 543028
rect 416832 542988 416838 543000
rect 482278 542988 482284 543000
rect 482336 542988 482342 543040
rect 498838 542988 498844 543040
rect 498896 543028 498902 543040
rect 511994 543028 512000 543040
rect 498896 543000 512000 543028
rect 498896 542988 498902 543000
rect 511994 542988 512000 543000
rect 512052 542988 512058 543040
rect 470594 542920 470600 542972
rect 470652 542960 470658 542972
rect 499022 542960 499028 542972
rect 470652 542932 499028 542960
rect 470652 542920 470658 542932
rect 499022 542920 499028 542932
rect 499080 542920 499086 542972
rect 476758 542852 476764 542904
rect 476816 542892 476822 542904
rect 506106 542892 506112 542904
rect 476816 542864 506112 542892
rect 476816 542852 476822 542864
rect 506106 542852 506112 542864
rect 506164 542852 506170 542904
rect 473354 542784 473360 542836
rect 473412 542824 473418 542836
rect 510614 542824 510620 542836
rect 473412 542796 510620 542824
rect 473412 542784 473418 542796
rect 510614 542784 510620 542796
rect 510672 542784 510678 542836
rect 472618 542716 472624 542768
rect 472676 542756 472682 542768
rect 515766 542756 515772 542768
rect 472676 542728 515772 542756
rect 472676 542716 472682 542728
rect 515766 542716 515772 542728
rect 515824 542716 515830 542768
rect 438854 542648 438860 542700
rect 438912 542688 438918 542700
rect 494054 542688 494060 542700
rect 438912 542660 494060 542688
rect 438912 542648 438918 542660
rect 494054 542648 494060 542660
rect 494112 542648 494118 542700
rect 279694 542580 279700 542632
rect 279752 542620 279758 542632
rect 279752 542592 287054 542620
rect 279752 542580 279758 542592
rect 279602 542512 279608 542564
rect 279660 542552 279666 542564
rect 287026 542552 287054 542592
rect 475470 542580 475476 542632
rect 475528 542620 475534 542632
rect 514754 542620 514760 542632
rect 475528 542592 514760 542620
rect 475528 542580 475534 542592
rect 514754 542580 514760 542592
rect 514812 542580 514818 542632
rect 292758 542552 292764 542564
rect 279660 542524 285168 542552
rect 287026 542524 292764 542552
rect 279660 542512 279666 542524
rect 279786 542444 279792 542496
rect 279844 542484 279850 542496
rect 285140 542484 285168 542524
rect 292758 542512 292764 542524
rect 292816 542512 292822 542564
rect 423674 542512 423680 542564
rect 423732 542552 423738 542564
rect 500310 542552 500316 542564
rect 423732 542524 500316 542552
rect 423732 542512 423738 542524
rect 500310 542512 500316 542524
rect 500368 542512 500374 542564
rect 503990 542512 503996 542564
rect 504048 542552 504054 542564
rect 540238 542552 540244 542564
rect 504048 542524 540244 542552
rect 504048 542512 504054 542524
rect 540238 542512 540244 542524
rect 540296 542512 540302 542564
rect 293954 542484 293960 542496
rect 279844 542456 285076 542484
rect 285140 542456 293960 542484
rect 279844 542444 279850 542456
rect 278314 542376 278320 542428
rect 278372 542416 278378 542428
rect 284938 542416 284944 542428
rect 278372 542388 284944 542416
rect 278372 542376 278378 542388
rect 284938 542376 284944 542388
rect 284996 542376 285002 542428
rect 285048 542416 285076 542456
rect 293954 542444 293960 542456
rect 294012 542444 294018 542496
rect 478230 542444 478236 542496
rect 478288 542484 478294 542496
rect 488166 542484 488172 542496
rect 478288 542456 488172 542484
rect 478288 542444 478294 542456
rect 488166 542444 488172 542456
rect 488224 542444 488230 542496
rect 295334 542416 295340 542428
rect 285048 542388 295340 542416
rect 295334 542376 295340 542388
rect 295392 542376 295398 542428
rect 466454 542376 466460 542428
rect 466512 542416 466518 542428
rect 484854 542416 484860 542428
rect 466512 542388 484860 542416
rect 466512 542376 466518 542388
rect 484854 542376 484860 542388
rect 484912 542376 484918 542428
rect 313274 541628 313280 541680
rect 313332 541668 313338 541680
rect 350166 541668 350172 541680
rect 313332 541640 350172 541668
rect 313332 541628 313338 541640
rect 350166 541628 350172 541640
rect 350224 541628 350230 541680
rect 406378 541356 406384 541408
rect 406436 541396 406442 541408
rect 493226 541396 493232 541408
rect 406436 541368 493232 541396
rect 406436 541356 406442 541368
rect 493226 541356 493232 541368
rect 493284 541356 493290 541408
rect 403618 541288 403624 541340
rect 403676 541328 403682 541340
rect 495434 541328 495440 541340
rect 403676 541300 495440 541328
rect 403676 541288 403682 541300
rect 495434 541288 495440 541300
rect 495492 541288 495498 541340
rect 475378 541220 475384 541272
rect 475436 541260 475442 541272
rect 511258 541260 511264 541272
rect 475436 541232 511264 541260
rect 475436 541220 475442 541232
rect 511258 541220 511264 541232
rect 511316 541220 511322 541272
rect 440878 541152 440884 541204
rect 440936 541192 440942 541204
rect 483014 541192 483020 541204
rect 440936 541164 483020 541192
rect 440936 541152 440942 541164
rect 483014 541152 483020 541164
rect 483072 541152 483078 541204
rect 484762 541152 484768 541204
rect 484820 541192 484826 541204
rect 542998 541192 543004 541204
rect 484820 541164 543004 541192
rect 484820 541152 484826 541164
rect 542998 541152 543004 541164
rect 543056 541152 543062 541204
rect 436830 541084 436836 541136
rect 436888 541124 436894 541136
rect 508682 541124 508688 541136
rect 436888 541096 508688 541124
rect 436888 541084 436894 541096
rect 508682 541084 508688 541096
rect 508740 541084 508746 541136
rect 492582 541016 492588 541068
rect 492640 541056 492646 541068
rect 556154 541056 556160 541068
rect 492640 541028 556160 541056
rect 492640 541016 492646 541028
rect 556154 541016 556160 541028
rect 556212 541016 556218 541068
rect 254394 540948 254400 541000
rect 254452 540988 254458 541000
rect 266998 540988 267004 541000
rect 254452 540960 267004 540988
rect 254452 540948 254458 540960
rect 266998 540948 267004 540960
rect 267056 540948 267062 541000
rect 401778 540948 401784 541000
rect 401836 540988 401842 541000
rect 437474 540988 437480 541000
rect 401836 540960 437480 540988
rect 401836 540948 401842 540960
rect 437474 540948 437480 540960
rect 437532 540948 437538 541000
rect 488074 540948 488080 541000
rect 488132 540988 488138 541000
rect 545114 540988 545120 541000
rect 488132 540960 545120 540988
rect 488132 540948 488138 540960
rect 545114 540948 545120 540960
rect 545172 540948 545178 541000
rect 306282 540268 306288 540320
rect 306340 540308 306346 540320
rect 347222 540308 347228 540320
rect 306340 540280 347228 540308
rect 306340 540268 306346 540280
rect 347222 540268 347228 540280
rect 347280 540268 347286 540320
rect 303522 540200 303528 540252
rect 303580 540240 303586 540252
rect 353294 540240 353300 540252
rect 303580 540212 353300 540240
rect 303580 540200 303586 540212
rect 353294 540200 353300 540212
rect 353352 540200 353358 540252
rect 402974 539996 402980 540048
rect 403032 540036 403038 540048
rect 500954 540036 500960 540048
rect 403032 540008 500960 540036
rect 403032 539996 403038 540008
rect 500954 539996 500960 540008
rect 501012 539996 501018 540048
rect 489822 539928 489828 539980
rect 489880 539968 489886 539980
rect 520274 539968 520280 539980
rect 489880 539940 520280 539968
rect 489880 539928 489886 539940
rect 520274 539928 520280 539940
rect 520332 539928 520338 539980
rect 486970 539860 486976 539912
rect 487028 539900 487034 539912
rect 547874 539900 547880 539912
rect 487028 539872 547880 539900
rect 487028 539860 487034 539872
rect 547874 539860 547880 539872
rect 547932 539860 547938 539912
rect 490650 539792 490656 539844
rect 490708 539832 490714 539844
rect 565814 539832 565820 539844
rect 490708 539804 565820 539832
rect 490708 539792 490714 539804
rect 565814 539792 565820 539804
rect 565872 539792 565878 539844
rect 410518 539724 410524 539776
rect 410576 539764 410582 539776
rect 496446 539764 496452 539776
rect 410576 539736 496452 539764
rect 410576 539724 410582 539736
rect 496446 539724 496452 539736
rect 496504 539724 496510 539776
rect 498194 539724 498200 539776
rect 498252 539764 498258 539776
rect 544378 539764 544384 539776
rect 498252 539736 544384 539764
rect 498252 539724 498258 539736
rect 544378 539724 544384 539736
rect 544436 539724 544442 539776
rect 493226 539656 493232 539708
rect 493284 539696 493290 539708
rect 525058 539696 525064 539708
rect 493284 539668 525064 539696
rect 493284 539656 493290 539668
rect 525058 539656 525064 539668
rect 525116 539656 525122 539708
rect 276658 539588 276664 539640
rect 276716 539628 276722 539640
rect 286410 539628 286416 539640
rect 276716 539600 286416 539628
rect 276716 539588 276722 539600
rect 286410 539588 286416 539600
rect 286468 539588 286474 539640
rect 404998 539588 405004 539640
rect 405056 539628 405062 539640
rect 518342 539628 518348 539640
rect 405056 539600 518348 539628
rect 405056 539588 405062 539600
rect 518342 539588 518348 539600
rect 518400 539588 518406 539640
rect 280798 539520 280804 539572
rect 280856 539560 280862 539572
rect 284202 539560 284208 539572
rect 280856 539532 284208 539560
rect 280856 539520 280862 539532
rect 284202 539520 284208 539532
rect 284260 539520 284266 539572
rect 332594 539520 332600 539572
rect 332652 539560 332658 539572
rect 357434 539560 357440 539572
rect 332652 539532 357440 539560
rect 332652 539520 332658 539532
rect 357434 539520 357440 539532
rect 357492 539520 357498 539572
rect 519630 539520 519636 539572
rect 519688 539560 519694 539572
rect 523034 539560 523040 539572
rect 519688 539532 523040 539560
rect 519688 539520 519694 539532
rect 523034 539520 523040 539532
rect 523092 539520 523098 539572
rect 322934 537548 322940 537600
rect 322992 537588 322998 537600
rect 358262 537588 358268 537600
rect 322992 537560 358268 537588
rect 322992 537548 322998 537560
rect 358262 537548 358268 537560
rect 358320 537548 358326 537600
rect 320174 537480 320180 537532
rect 320232 537520 320238 537532
rect 356698 537520 356704 537532
rect 320232 537492 356704 537520
rect 320232 537480 320238 537492
rect 356698 537480 356704 537492
rect 356756 537480 356762 537532
rect 358262 536868 358268 536920
rect 358320 536908 358326 536920
rect 358906 536908 358912 536920
rect 358320 536880 358912 536908
rect 358320 536868 358326 536880
rect 358906 536868 358912 536880
rect 358964 536868 358970 536920
rect 358446 536800 358452 536852
rect 358504 536840 358510 536852
rect 359550 536840 359556 536852
rect 358504 536812 359556 536840
rect 358504 536800 358510 536812
rect 359550 536800 359556 536812
rect 359608 536800 359614 536852
rect 523678 536800 523684 536852
rect 523736 536840 523742 536852
rect 580166 536840 580172 536852
rect 523736 536812 580172 536840
rect 523736 536800 523742 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 347038 536732 347044 536784
rect 347096 536772 347102 536784
rect 357434 536772 357440 536784
rect 347096 536744 357440 536772
rect 347096 536732 347102 536744
rect 357434 536732 357440 536744
rect 357492 536732 357498 536784
rect 355410 536664 355416 536716
rect 355468 536704 355474 536716
rect 357894 536704 357900 536716
rect 355468 536676 357900 536704
rect 355468 536664 355474 536676
rect 357894 536664 357900 536676
rect 357952 536664 357958 536716
rect 522206 535644 522212 535696
rect 522264 535684 522270 535696
rect 525150 535684 525156 535696
rect 522264 535656 525156 535684
rect 522264 535644 522270 535656
rect 525150 535644 525156 535656
rect 525208 535644 525214 535696
rect 357526 535508 357532 535560
rect 357584 535548 357590 535560
rect 357584 535520 357664 535548
rect 357584 535508 357590 535520
rect 354214 535372 354220 535424
rect 354272 535412 354278 535424
rect 357526 535412 357532 535424
rect 354272 535384 357532 535412
rect 354272 535372 354278 535384
rect 357526 535372 357532 535384
rect 357584 535372 357590 535424
rect 357636 535412 357664 535520
rect 359642 535412 359648 535424
rect 357636 535384 359648 535412
rect 359642 535372 359648 535384
rect 359700 535372 359706 535424
rect 322106 535304 322112 535356
rect 322164 535344 322170 535356
rect 352374 535344 352380 535356
rect 322164 535316 352380 535344
rect 322164 535304 322170 535316
rect 352374 535304 352380 535316
rect 352432 535304 352438 535356
rect 354306 535304 354312 535356
rect 354364 535344 354370 535356
rect 357894 535344 357900 535356
rect 354364 535316 357900 535344
rect 354364 535304 354370 535316
rect 357894 535304 357900 535316
rect 357952 535304 357958 535356
rect 337470 535236 337476 535288
rect 337528 535276 337534 535288
rect 357434 535276 357440 535288
rect 337528 535248 357440 535276
rect 337528 535236 337534 535248
rect 357434 535236 357440 535248
rect 357492 535236 357498 535288
rect 322474 535168 322480 535220
rect 322532 535208 322538 535220
rect 355134 535208 355140 535220
rect 322532 535180 355140 535208
rect 322532 535168 322538 535180
rect 355134 535168 355140 535180
rect 355192 535168 355198 535220
rect 322566 534692 322572 534744
rect 322624 534732 322630 534744
rect 337930 534732 337936 534744
rect 322624 534704 337936 534732
rect 322624 534692 322630 534704
rect 337930 534692 337936 534704
rect 337988 534692 337994 534744
rect 254578 534080 254584 534132
rect 254636 534120 254642 534132
rect 278130 534120 278136 534132
rect 254636 534092 278136 534120
rect 254636 534080 254642 534092
rect 278130 534080 278136 534092
rect 278188 534080 278194 534132
rect 400858 534080 400864 534132
rect 400916 534120 400922 534132
rect 402054 534120 402060 534132
rect 400916 534092 402060 534120
rect 400916 534080 400922 534092
rect 402054 534080 402060 534092
rect 402112 534080 402118 534132
rect 401594 533876 401600 533928
rect 401652 533916 401658 533928
rect 404906 533916 404912 533928
rect 401652 533888 404912 533916
rect 401652 533876 401658 533888
rect 404906 533876 404912 533888
rect 404964 533876 404970 533928
rect 322474 533400 322480 533452
rect 322532 533440 322538 533452
rect 329558 533440 329564 533452
rect 322532 533412 329564 533440
rect 322532 533400 322538 533412
rect 329558 533400 329564 533412
rect 329616 533400 329622 533452
rect 338022 533400 338028 533452
rect 338080 533440 338086 533452
rect 357526 533440 357532 533452
rect 338080 533412 357532 533440
rect 338080 533400 338086 533412
rect 357526 533400 357532 533412
rect 357584 533400 357590 533452
rect 322842 533332 322848 533384
rect 322900 533372 322906 533384
rect 357158 533372 357164 533384
rect 322900 533344 357164 533372
rect 322900 533332 322906 533344
rect 357158 533332 357164 533344
rect 357216 533332 357222 533384
rect 423030 533332 423036 533384
rect 423088 533372 423094 533384
rect 477586 533372 477592 533384
rect 423088 533344 477592 533372
rect 423088 533332 423094 533344
rect 477586 533332 477592 533344
rect 477644 533332 477650 533384
rect 454770 532720 454776 532772
rect 454828 532760 454834 532772
rect 477586 532760 477592 532772
rect 454828 532732 477592 532760
rect 454828 532720 454834 532732
rect 477586 532720 477592 532732
rect 477644 532720 477650 532772
rect 321646 532652 321652 532704
rect 321704 532692 321710 532704
rect 352466 532692 352472 532704
rect 321704 532664 352472 532692
rect 321704 532652 321710 532664
rect 352466 532652 352472 532664
rect 352524 532652 352530 532704
rect 353294 532652 353300 532704
rect 353352 532692 353358 532704
rect 357526 532692 357532 532704
rect 353352 532664 357532 532692
rect 353352 532652 353358 532664
rect 357526 532652 357532 532664
rect 357584 532652 357590 532704
rect 522942 532652 522948 532704
rect 523000 532692 523006 532704
rect 534718 532692 534724 532704
rect 523000 532664 534724 532692
rect 523000 532652 523006 532664
rect 534718 532652 534724 532664
rect 534776 532652 534782 532704
rect 345750 532584 345756 532636
rect 345808 532624 345814 532636
rect 357434 532624 357440 532636
rect 345808 532596 357440 532624
rect 345808 532584 345814 532596
rect 357434 532584 357440 532596
rect 357492 532584 357498 532636
rect 329558 531972 329564 532024
rect 329616 532012 329622 532024
rect 336090 532012 336096 532024
rect 329616 531984 336096 532012
rect 329616 531972 329622 531984
rect 336090 531972 336096 531984
rect 336148 532012 336154 532024
rect 342990 532012 342996 532024
rect 336148 531984 342996 532012
rect 336148 531972 336154 531984
rect 342990 531972 342996 531984
rect 343048 531972 343054 532024
rect 463694 531292 463700 531344
rect 463752 531332 463758 531344
rect 477586 531332 477592 531344
rect 463752 531304 477592 531332
rect 463752 531292 463758 531304
rect 477586 531292 477592 531304
rect 477644 531292 477650 531344
rect 322474 531224 322480 531276
rect 322532 531264 322538 531276
rect 338022 531264 338028 531276
rect 322532 531236 338028 531264
rect 322532 531224 322538 531236
rect 338022 531224 338028 531236
rect 338080 531224 338086 531276
rect 458818 531224 458824 531276
rect 458876 531264 458882 531276
rect 478690 531264 478696 531276
rect 458876 531236 478696 531264
rect 458876 531224 458882 531236
rect 478690 531224 478696 531236
rect 478748 531224 478754 531276
rect 322658 530544 322664 530596
rect 322716 530584 322722 530596
rect 350534 530584 350540 530596
rect 322716 530556 350540 530584
rect 322716 530544 322722 530556
rect 350534 530544 350540 530556
rect 350592 530544 350598 530596
rect 401594 530204 401600 530256
rect 401652 530244 401658 530256
rect 403526 530244 403532 530256
rect 401652 530216 403532 530244
rect 401652 530204 401658 530216
rect 403526 530204 403532 530216
rect 403584 530204 403590 530256
rect 322566 529932 322572 529984
rect 322624 529972 322630 529984
rect 357158 529972 357164 529984
rect 322624 529944 357164 529972
rect 322624 529932 322630 529944
rect 357158 529932 357164 529944
rect 357216 529932 357222 529984
rect 401778 529932 401784 529984
rect 401836 529972 401842 529984
rect 458174 529972 458180 529984
rect 401836 529944 458180 529972
rect 401836 529932 401842 529944
rect 458174 529932 458180 529944
rect 458232 529932 458238 529984
rect 322474 529864 322480 529916
rect 322532 529904 322538 529916
rect 351270 529904 351276 529916
rect 322532 529876 351276 529904
rect 322532 529864 322538 529876
rect 351270 529864 351276 529876
rect 351328 529864 351334 529916
rect 338850 529796 338856 529848
rect 338908 529836 338914 529848
rect 357434 529836 357440 529848
rect 338908 529808 357440 529836
rect 338908 529796 338914 529808
rect 357434 529796 357440 529808
rect 357492 529796 357498 529848
rect 322474 529660 322480 529712
rect 322532 529700 322538 529712
rect 322842 529700 322848 529712
rect 322532 529672 322848 529700
rect 322532 529660 322538 529672
rect 322842 529660 322848 529672
rect 322900 529660 322906 529712
rect 401594 529116 401600 529168
rect 401652 529156 401658 529168
rect 403802 529156 403808 529168
rect 401652 529128 403808 529156
rect 401652 529116 401658 529128
rect 403802 529116 403808 529128
rect 403860 529116 403866 529168
rect 401778 528640 401784 528692
rect 401836 528680 401842 528692
rect 405090 528680 405096 528692
rect 401836 528652 405096 528680
rect 401836 528640 401842 528652
rect 405090 528640 405096 528652
rect 405148 528640 405154 528692
rect 254578 528572 254584 528624
rect 254636 528612 254642 528624
rect 273990 528612 273996 528624
rect 254636 528584 273996 528612
rect 254636 528572 254642 528584
rect 273990 528572 273996 528584
rect 274048 528572 274054 528624
rect 452654 528572 452660 528624
rect 452712 528612 452718 528624
rect 477586 528612 477592 528624
rect 452712 528584 477592 528612
rect 452712 528572 452718 528584
rect 477586 528572 477592 528584
rect 477644 528572 477650 528624
rect 322106 528504 322112 528556
rect 322164 528544 322170 528556
rect 355226 528544 355232 528556
rect 322164 528516 355232 528544
rect 322164 528504 322170 528516
rect 355226 528504 355232 528516
rect 355284 528504 355290 528556
rect 401594 528436 401600 528488
rect 401652 528476 401658 528488
rect 404446 528476 404452 528488
rect 401652 528448 404452 528476
rect 401652 528436 401658 528448
rect 404446 528436 404452 528448
rect 404504 528436 404510 528488
rect 322566 527144 322572 527196
rect 322624 527184 322630 527196
rect 322750 527184 322756 527196
rect 322624 527156 322756 527184
rect 322624 527144 322630 527156
rect 322750 527144 322756 527156
rect 322808 527144 322814 527196
rect 418798 527144 418804 527196
rect 418856 527184 418862 527196
rect 477586 527184 477592 527196
rect 418856 527156 477592 527184
rect 418856 527144 418862 527156
rect 477586 527144 477592 527156
rect 477644 527144 477650 527196
rect 322198 527076 322204 527128
rect 322256 527116 322262 527128
rect 357434 527116 357440 527128
rect 322256 527088 357440 527116
rect 322256 527076 322262 527088
rect 357434 527076 357440 527088
rect 357492 527076 357498 527128
rect 412634 527076 412640 527128
rect 412692 527116 412698 527128
rect 477678 527116 477684 527128
rect 412692 527088 477684 527116
rect 412692 527076 412698 527088
rect 477678 527076 477684 527088
rect 477736 527076 477742 527128
rect 322474 527008 322480 527060
rect 322532 527048 322538 527060
rect 354398 527048 354404 527060
rect 322532 527020 354404 527048
rect 322532 527008 322538 527020
rect 354398 527008 354404 527020
rect 354456 527008 354462 527060
rect 355318 527008 355324 527060
rect 355376 527048 355382 527060
rect 357526 527048 357532 527060
rect 355376 527020 357532 527048
rect 355376 527008 355382 527020
rect 357526 527008 357532 527020
rect 357584 527008 357590 527060
rect 322566 526940 322572 526992
rect 322624 526980 322630 526992
rect 326338 526980 326344 526992
rect 322624 526952 326344 526980
rect 322624 526940 322630 526952
rect 326338 526940 326344 526952
rect 326396 526940 326402 526992
rect 401594 526396 401600 526448
rect 401652 526436 401658 526448
rect 403250 526436 403256 526448
rect 401652 526408 403256 526436
rect 401652 526396 401658 526408
rect 403250 526396 403256 526408
rect 403308 526396 403314 526448
rect 358262 525784 358268 525836
rect 358320 525824 358326 525836
rect 359458 525824 359464 525836
rect 358320 525796 359464 525824
rect 358320 525784 358326 525796
rect 359458 525784 359464 525796
rect 359516 525784 359522 525836
rect 400398 525784 400404 525836
rect 400456 525824 400462 525836
rect 432598 525824 432604 525836
rect 400456 525796 432604 525824
rect 400456 525784 400462 525796
rect 432598 525784 432604 525796
rect 432656 525784 432662 525836
rect 460198 525784 460204 525836
rect 460256 525824 460262 525836
rect 477586 525824 477592 525836
rect 460256 525796 477592 525824
rect 460256 525784 460262 525796
rect 477586 525784 477592 525796
rect 477644 525784 477650 525836
rect 522942 525784 522948 525836
rect 523000 525824 523006 525836
rect 536098 525824 536104 525836
rect 523000 525796 536104 525824
rect 523000 525784 523006 525796
rect 536098 525784 536104 525796
rect 536156 525784 536162 525836
rect 401594 525716 401600 525768
rect 401652 525756 401658 525768
rect 404630 525756 404636 525768
rect 401652 525728 404636 525756
rect 401652 525716 401658 525728
rect 404630 525716 404636 525728
rect 404688 525716 404694 525768
rect 527818 525716 527824 525768
rect 527876 525756 527882 525768
rect 579798 525756 579804 525768
rect 527876 525728 579804 525756
rect 527876 525716 527882 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 401594 525240 401600 525292
rect 401652 525280 401658 525292
rect 404354 525280 404360 525292
rect 401652 525252 404360 525280
rect 401652 525240 401658 525252
rect 404354 525240 404360 525252
rect 404412 525240 404418 525292
rect 322842 525036 322848 525088
rect 322900 525076 322906 525088
rect 348510 525076 348516 525088
rect 322900 525048 348516 525076
rect 322900 525036 322906 525048
rect 348510 525036 348516 525048
rect 348568 525036 348574 525088
rect 422938 524424 422944 524476
rect 422996 524464 423002 524476
rect 478138 524464 478144 524476
rect 422996 524436 478144 524464
rect 422996 524424 423002 524436
rect 478138 524424 478144 524436
rect 478196 524424 478202 524476
rect 334618 524356 334624 524408
rect 334676 524396 334682 524408
rect 357434 524396 357440 524408
rect 334676 524368 357440 524396
rect 334676 524356 334682 524368
rect 357434 524356 357440 524368
rect 357492 524356 357498 524408
rect 401594 524356 401600 524408
rect 401652 524396 401658 524408
rect 404814 524396 404820 524408
rect 401652 524368 404820 524396
rect 401652 524356 401658 524368
rect 404814 524356 404820 524368
rect 404872 524356 404878 524408
rect 322658 523676 322664 523728
rect 322716 523716 322722 523728
rect 355226 523716 355232 523728
rect 322716 523688 355232 523716
rect 322716 523676 322722 523688
rect 355226 523676 355232 523688
rect 355284 523676 355290 523728
rect 254302 522996 254308 523048
rect 254360 523036 254366 523048
rect 274082 523036 274088 523048
rect 254360 523008 274088 523036
rect 254360 522996 254366 523008
rect 274082 522996 274088 523008
rect 274140 522996 274146 523048
rect 522942 522996 522948 523048
rect 523000 523036 523006 523048
rect 534718 523036 534724 523048
rect 523000 523008 534724 523036
rect 523000 522996 523006 523008
rect 534718 522996 534724 523008
rect 534776 522996 534782 523048
rect 322566 522928 322572 522980
rect 322624 522968 322630 522980
rect 348418 522968 348424 522980
rect 322624 522940 348424 522968
rect 322624 522928 322630 522940
rect 348418 522928 348424 522940
rect 348476 522928 348482 522980
rect 322474 522248 322480 522300
rect 322532 522288 322538 522300
rect 352466 522288 352472 522300
rect 322532 522260 352472 522288
rect 322532 522248 322538 522260
rect 352466 522248 352472 522260
rect 352524 522248 352530 522300
rect 322106 521908 322112 521960
rect 322164 521948 322170 521960
rect 322658 521948 322664 521960
rect 322164 521920 322664 521948
rect 322164 521908 322170 521920
rect 322658 521908 322664 521920
rect 322716 521908 322722 521960
rect 401594 521636 401600 521688
rect 401652 521676 401658 521688
rect 423766 521676 423772 521688
rect 401652 521648 423772 521676
rect 401652 521636 401658 521648
rect 423766 521636 423772 521648
rect 423824 521636 423830 521688
rect 322474 521568 322480 521620
rect 322532 521608 322538 521620
rect 353202 521608 353208 521620
rect 322532 521580 353208 521608
rect 322532 521568 322538 521580
rect 353202 521568 353208 521580
rect 353260 521568 353266 521620
rect 401594 521024 401600 521076
rect 401652 521064 401658 521076
rect 403434 521064 403440 521076
rect 401652 521036 403440 521064
rect 401652 521024 401658 521036
rect 403434 521024 403440 521036
rect 403492 521024 403498 521076
rect 322198 520888 322204 520940
rect 322256 520928 322262 520940
rect 351270 520928 351276 520940
rect 322256 520900 351276 520928
rect 322256 520888 322262 520900
rect 351270 520888 351276 520900
rect 351328 520888 351334 520940
rect 322198 520752 322204 520804
rect 322256 520792 322262 520804
rect 322382 520792 322388 520804
rect 322256 520764 322388 520792
rect 322256 520752 322262 520764
rect 322382 520752 322388 520764
rect 322440 520752 322446 520804
rect 522942 520616 522948 520668
rect 523000 520656 523006 520668
rect 530578 520656 530584 520668
rect 523000 520628 530584 520656
rect 523000 520616 523006 520628
rect 530578 520616 530584 520628
rect 530636 520616 530642 520668
rect 322014 520276 322020 520328
rect 322072 520316 322078 520328
rect 347038 520316 347044 520328
rect 322072 520288 347044 520316
rect 322072 520276 322078 520288
rect 347038 520276 347044 520288
rect 347096 520276 347102 520328
rect 321646 520208 321652 520260
rect 321704 520248 321710 520260
rect 321704 520220 335354 520248
rect 321704 520208 321710 520220
rect 335326 520180 335354 520220
rect 353018 520208 353024 520260
rect 353076 520248 353082 520260
rect 357434 520248 357440 520260
rect 353076 520220 357440 520248
rect 353076 520208 353082 520220
rect 357434 520208 357440 520220
rect 357492 520208 357498 520260
rect 347682 520180 347688 520192
rect 335326 520152 347688 520180
rect 347682 520140 347688 520152
rect 347740 520180 347746 520192
rect 354214 520180 354220 520192
rect 347740 520152 354220 520180
rect 347740 520140 347746 520152
rect 354214 520140 354220 520152
rect 354272 520140 354278 520192
rect 401594 520140 401600 520192
rect 401652 520180 401658 520192
rect 405274 520180 405280 520192
rect 401652 520152 405280 520180
rect 401652 520140 401658 520152
rect 405274 520140 405280 520152
rect 405332 520140 405338 520192
rect 322198 519256 322204 519308
rect 322256 519296 322262 519308
rect 325050 519296 325056 519308
rect 322256 519268 325056 519296
rect 322256 519256 322262 519268
rect 325050 519256 325056 519268
rect 325108 519256 325114 519308
rect 414014 518916 414020 518968
rect 414072 518956 414078 518968
rect 477586 518956 477592 518968
rect 414072 518928 477592 518956
rect 414072 518916 414078 518928
rect 477586 518916 477592 518928
rect 477644 518916 477650 518968
rect 350074 518848 350080 518900
rect 350132 518888 350138 518900
rect 357434 518888 357440 518900
rect 350132 518860 357440 518888
rect 350132 518848 350138 518860
rect 357434 518848 357440 518860
rect 357492 518848 357498 518900
rect 321738 518032 321744 518084
rect 321796 518072 321802 518084
rect 324222 518072 324228 518084
rect 321796 518044 324228 518072
rect 321796 518032 321802 518044
rect 324222 518032 324228 518044
rect 324280 518032 324286 518084
rect 254578 517760 254584 517812
rect 254636 517800 254642 517812
rect 258718 517800 258724 517812
rect 254636 517772 258724 517800
rect 254636 517760 254642 517772
rect 258718 517760 258724 517772
rect 258776 517760 258782 517812
rect 324314 517624 324320 517676
rect 324372 517664 324378 517676
rect 325510 517664 325516 517676
rect 324372 517636 325516 517664
rect 324372 517624 324378 517636
rect 325510 517624 325516 517636
rect 325568 517664 325574 517676
rect 350718 517664 350724 517676
rect 325568 517636 350724 517664
rect 325568 517624 325574 517636
rect 350718 517624 350724 517636
rect 350776 517624 350782 517676
rect 322290 517556 322296 517608
rect 322348 517596 322354 517608
rect 350626 517596 350632 517608
rect 322348 517568 350632 517596
rect 322348 517556 322354 517568
rect 350626 517556 350632 517568
rect 350684 517596 350690 517608
rect 355870 517596 355876 517608
rect 350684 517568 355876 517596
rect 350684 517556 350690 517568
rect 355870 517556 355876 517568
rect 355928 517556 355934 517608
rect 468478 517556 468484 517608
rect 468536 517596 468542 517608
rect 477586 517596 477592 517608
rect 468536 517568 477592 517596
rect 468536 517556 468542 517568
rect 477586 517556 477592 517568
rect 477644 517556 477650 517608
rect 329190 517488 329196 517540
rect 329248 517528 329254 517540
rect 357526 517528 357532 517540
rect 329248 517500 357532 517528
rect 329248 517488 329254 517500
rect 357526 517488 357532 517500
rect 357584 517488 357590 517540
rect 450538 517488 450544 517540
rect 450596 517528 450602 517540
rect 477678 517528 477684 517540
rect 450596 517500 477684 517528
rect 450596 517488 450602 517500
rect 477678 517488 477684 517500
rect 477736 517488 477742 517540
rect 322842 517420 322848 517472
rect 322900 517460 322906 517472
rect 324314 517460 324320 517472
rect 322900 517432 324320 517460
rect 322900 517420 322906 517432
rect 324314 517420 324320 517432
rect 324372 517420 324378 517472
rect 340138 517420 340144 517472
rect 340196 517460 340202 517472
rect 357434 517460 357440 517472
rect 340196 517432 357440 517460
rect 340196 517420 340202 517432
rect 357434 517420 357440 517432
rect 357492 517420 357498 517472
rect 427078 517420 427084 517472
rect 427136 517460 427142 517472
rect 477586 517460 477592 517472
rect 427136 517432 477592 517460
rect 427136 517420 427142 517432
rect 477586 517420 477592 517432
rect 477644 517420 477650 517472
rect 401594 516128 401600 516180
rect 401652 516168 401658 516180
rect 405734 516168 405740 516180
rect 401652 516140 405740 516168
rect 401652 516128 401658 516140
rect 405734 516128 405740 516140
rect 405792 516128 405798 516180
rect 322290 516060 322296 516112
rect 322348 516100 322354 516112
rect 342254 516100 342260 516112
rect 322348 516072 342260 516100
rect 322348 516060 322354 516072
rect 342254 516060 342260 516072
rect 342312 516060 342318 516112
rect 401686 516060 401692 516112
rect 401744 516100 401750 516112
rect 404722 516100 404728 516112
rect 401744 516072 404728 516100
rect 401744 516060 401750 516072
rect 404722 516060 404728 516072
rect 404780 516060 404786 516112
rect 322842 515380 322848 515432
rect 322900 515420 322906 515432
rect 324222 515420 324228 515432
rect 322900 515392 324228 515420
rect 322900 515380 322906 515392
rect 324222 515380 324228 515392
rect 324280 515420 324286 515432
rect 331950 515420 331956 515432
rect 324280 515392 331956 515420
rect 324280 515380 324286 515392
rect 331950 515380 331956 515392
rect 332008 515380 332014 515432
rect 342254 515380 342260 515432
rect 342312 515420 342318 515432
rect 343542 515420 343548 515432
rect 342312 515392 343548 515420
rect 342312 515380 342318 515392
rect 343542 515380 343548 515392
rect 343600 515420 343606 515432
rect 355410 515420 355416 515432
rect 343600 515392 355416 515420
rect 343600 515380 343606 515392
rect 355410 515380 355416 515392
rect 355468 515380 355474 515432
rect 457438 514836 457444 514888
rect 457496 514876 457502 514888
rect 477586 514876 477592 514888
rect 457496 514848 477592 514876
rect 457496 514836 457502 514848
rect 477586 514836 477592 514848
rect 477644 514836 477650 514888
rect 400858 514768 400864 514820
rect 400916 514808 400922 514820
rect 477678 514808 477684 514820
rect 400916 514780 477684 514808
rect 400916 514768 400922 514780
rect 477678 514768 477684 514780
rect 477736 514768 477742 514820
rect 342898 514700 342904 514752
rect 342956 514740 342962 514752
rect 357434 514740 357440 514752
rect 342956 514712 357440 514740
rect 342956 514700 342962 514712
rect 357434 514700 357440 514712
rect 357492 514700 357498 514752
rect 358630 514292 358636 514344
rect 358688 514332 358694 514344
rect 359826 514332 359832 514344
rect 358688 514304 359832 514332
rect 358688 514292 358694 514304
rect 359826 514292 359832 514304
rect 359884 514292 359890 514344
rect 322750 514020 322756 514072
rect 322808 514060 322814 514072
rect 322934 514060 322940 514072
rect 322808 514032 322940 514060
rect 322808 514020 322814 514032
rect 322934 514020 322940 514032
rect 322992 514060 322998 514072
rect 329098 514060 329104 514072
rect 322992 514032 329104 514060
rect 322992 514020 322998 514032
rect 329098 514020 329104 514032
rect 329156 514020 329162 514072
rect 322290 513408 322296 513460
rect 322348 513448 322354 513460
rect 355318 513448 355324 513460
rect 322348 513420 355324 513448
rect 322348 513408 322354 513420
rect 355318 513408 355324 513420
rect 355376 513408 355382 513460
rect 413278 513340 413284 513392
rect 413336 513380 413342 513392
rect 477586 513380 477592 513392
rect 413336 513352 477592 513380
rect 413336 513340 413342 513352
rect 477586 513340 477592 513352
rect 477644 513340 477650 513392
rect 331858 513272 331864 513324
rect 331916 513312 331922 513324
rect 357434 513312 357440 513324
rect 331916 513284 357440 513312
rect 331916 513272 331922 513284
rect 357434 513272 357440 513284
rect 357492 513272 357498 513324
rect 522850 513204 522856 513256
rect 522908 513244 522914 513256
rect 526438 513244 526444 513256
rect 522908 513216 526444 513244
rect 522908 513204 522914 513216
rect 526438 513204 526444 513216
rect 526496 513204 526502 513256
rect 402422 513068 402428 513120
rect 402480 513108 402486 513120
rect 405366 513108 405372 513120
rect 402480 513080 405372 513108
rect 402480 513068 402486 513080
rect 405366 513068 405372 513080
rect 405424 513068 405430 513120
rect 322198 512592 322204 512644
rect 322256 512632 322262 512644
rect 331214 512632 331220 512644
rect 322256 512604 331220 512632
rect 322256 512592 322262 512604
rect 331214 512592 331220 512604
rect 331272 512592 331278 512644
rect 476850 512048 476856 512100
rect 476908 512088 476914 512100
rect 478138 512088 478144 512100
rect 476908 512060 478144 512088
rect 476908 512048 476914 512060
rect 478138 512048 478144 512060
rect 478196 512048 478202 512100
rect 436738 511980 436744 512032
rect 436796 512020 436802 512032
rect 477678 512020 477684 512032
rect 436796 511992 477684 512020
rect 436796 511980 436802 511992
rect 477678 511980 477684 511992
rect 477736 511980 477742 512032
rect 322198 511912 322204 511964
rect 322256 511952 322262 511964
rect 355778 511952 355784 511964
rect 322256 511924 355784 511952
rect 322256 511912 322262 511924
rect 355778 511912 355784 511924
rect 355836 511912 355842 511964
rect 358078 511912 358084 511964
rect 358136 511952 358142 511964
rect 359458 511952 359464 511964
rect 358136 511924 359464 511952
rect 358136 511912 358142 511924
rect 359458 511912 359464 511924
rect 359516 511912 359522 511964
rect 432598 511912 432604 511964
rect 432656 511952 432662 511964
rect 477586 511952 477592 511964
rect 432656 511924 477592 511952
rect 432656 511912 432662 511924
rect 477586 511912 477592 511924
rect 477644 511912 477650 511964
rect 320082 511844 320088 511896
rect 320140 511884 320146 511896
rect 345842 511884 345848 511896
rect 320140 511856 345848 511884
rect 320140 511844 320146 511856
rect 345842 511844 345848 511856
rect 345900 511844 345906 511896
rect 347222 511844 347228 511896
rect 347280 511884 347286 511896
rect 357434 511884 357440 511896
rect 347280 511856 357440 511884
rect 347280 511844 347286 511856
rect 357434 511844 357440 511856
rect 357492 511844 357498 511896
rect 321554 511232 321560 511284
rect 321612 511272 321618 511284
rect 333882 511272 333888 511284
rect 321612 511244 333888 511272
rect 321612 511232 321618 511244
rect 333882 511232 333888 511244
rect 333940 511272 333946 511284
rect 357250 511272 357256 511284
rect 333940 511244 357256 511272
rect 333940 511232 333946 511244
rect 357250 511232 357256 511244
rect 357308 511232 357314 511284
rect 522942 510688 522948 510740
rect 523000 510728 523006 510740
rect 538858 510728 538864 510740
rect 523000 510700 538864 510728
rect 523000 510688 523006 510700
rect 538858 510688 538864 510700
rect 538916 510688 538922 510740
rect 254394 510620 254400 510672
rect 254452 510660 254458 510672
rect 271230 510660 271236 510672
rect 254452 510632 271236 510660
rect 254452 510620 254458 510632
rect 271230 510620 271236 510632
rect 271288 510620 271294 510672
rect 319070 510620 319076 510672
rect 319128 510660 319134 510672
rect 320082 510660 320088 510672
rect 319128 510632 320088 510660
rect 319128 510620 319134 510632
rect 320082 510620 320088 510632
rect 320140 510620 320146 510672
rect 402882 510620 402888 510672
rect 402940 510660 402946 510672
rect 451274 510660 451280 510672
rect 402940 510632 451280 510660
rect 402940 510620 402946 510632
rect 451274 510620 451280 510632
rect 451332 510620 451338 510672
rect 526438 510620 526444 510672
rect 526496 510660 526502 510672
rect 580166 510660 580172 510672
rect 526496 510632 580172 510660
rect 526496 510620 526502 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 320358 510552 320364 510604
rect 320416 510592 320422 510604
rect 341610 510592 341616 510604
rect 320416 510564 341616 510592
rect 320416 510552 320422 510564
rect 341610 510552 341616 510564
rect 341668 510552 341674 510604
rect 342990 510552 342996 510604
rect 343048 510592 343054 510604
rect 357434 510592 357440 510604
rect 343048 510564 357440 510592
rect 343048 510552 343054 510564
rect 357434 510552 357440 510564
rect 357492 510552 357498 510604
rect 476942 510484 476948 510536
rect 477000 510524 477006 510536
rect 478138 510524 478144 510536
rect 477000 510496 478144 510524
rect 477000 510484 477006 510496
rect 478138 510484 478144 510496
rect 478196 510484 478202 510536
rect 324222 509872 324228 509924
rect 324280 509912 324286 509924
rect 350074 509912 350080 509924
rect 324280 509884 350080 509912
rect 324280 509872 324286 509884
rect 350074 509872 350080 509884
rect 350132 509872 350138 509924
rect 427722 509872 427728 509924
rect 427780 509912 427786 509924
rect 468662 509912 468668 509924
rect 427780 509884 468668 509912
rect 427780 509872 427786 509884
rect 468662 509872 468668 509884
rect 468720 509872 468726 509924
rect 402882 509260 402888 509312
rect 402940 509300 402946 509312
rect 427722 509300 427728 509312
rect 402940 509272 427728 509300
rect 402940 509260 402946 509272
rect 427722 509260 427728 509272
rect 427780 509260 427786 509312
rect 468570 509260 468576 509312
rect 468628 509300 468634 509312
rect 477586 509300 477592 509312
rect 468628 509272 477592 509300
rect 468628 509260 468634 509272
rect 477586 509260 477592 509272
rect 477644 509260 477650 509312
rect 322290 509192 322296 509244
rect 322348 509232 322354 509244
rect 355594 509232 355600 509244
rect 322348 509204 355600 509232
rect 322348 509192 322354 509204
rect 355594 509192 355600 509204
rect 355652 509192 355658 509244
rect 327718 509124 327724 509176
rect 327776 509164 327782 509176
rect 357986 509164 357992 509176
rect 327776 509136 357992 509164
rect 327776 509124 327782 509136
rect 357986 509124 357992 509136
rect 358044 509124 358050 509176
rect 345658 509056 345664 509108
rect 345716 509096 345722 509108
rect 357434 509096 357440 509108
rect 345716 509068 357440 509096
rect 345716 509056 345722 509068
rect 357434 509056 357440 509068
rect 357492 509056 357498 509108
rect 50798 508716 50804 508768
rect 50856 508756 50862 508768
rect 51258 508756 51264 508768
rect 50856 508728 51264 508756
rect 50856 508716 50862 508728
rect 51258 508716 51264 508728
rect 51316 508716 51322 508768
rect 321646 508580 321652 508632
rect 321704 508620 321710 508632
rect 322290 508620 322296 508632
rect 321704 508592 322296 508620
rect 321704 508580 321710 508592
rect 322290 508580 322296 508592
rect 322348 508580 322354 508632
rect 318886 508240 318892 508292
rect 318944 508280 318950 508292
rect 319346 508280 319352 508292
rect 318944 508252 319352 508280
rect 318944 508240 318950 508252
rect 319346 508240 319352 508252
rect 319404 508240 319410 508292
rect 320266 508104 320272 508156
rect 320324 508144 320330 508156
rect 320634 508144 320640 508156
rect 320324 508116 320640 508144
rect 320324 508104 320330 508116
rect 320634 508104 320640 508116
rect 320692 508144 320698 508156
rect 327810 508144 327816 508156
rect 320692 508116 327816 508144
rect 320692 508104 320698 508116
rect 327810 508104 327816 508116
rect 327868 508104 327874 508156
rect 319346 507832 319352 507884
rect 319404 507872 319410 507884
rect 356606 507872 356612 507884
rect 319404 507844 356612 507872
rect 319404 507832 319410 507844
rect 356606 507832 356612 507844
rect 356664 507832 356670 507884
rect 445754 507832 445760 507884
rect 445812 507872 445818 507884
rect 478138 507872 478144 507884
rect 445812 507844 478144 507872
rect 445812 507832 445818 507844
rect 478138 507832 478144 507844
rect 478196 507832 478202 507884
rect 320266 507764 320272 507816
rect 320324 507804 320330 507816
rect 320542 507804 320548 507816
rect 320324 507776 320548 507804
rect 320324 507764 320330 507776
rect 320542 507764 320548 507776
rect 320600 507804 320606 507816
rect 355686 507804 355692 507816
rect 320600 507776 355692 507804
rect 320600 507764 320606 507776
rect 355686 507764 355692 507776
rect 355744 507764 355750 507816
rect 335998 507696 336004 507748
rect 336056 507736 336062 507748
rect 357434 507736 357440 507748
rect 336056 507708 357440 507736
rect 336056 507696 336062 507708
rect 357434 507696 357440 507708
rect 357492 507696 357498 507748
rect 318886 506472 318892 506524
rect 318944 506512 318950 506524
rect 319346 506512 319352 506524
rect 318944 506484 319352 506512
rect 318944 506472 318950 506484
rect 319346 506472 319352 506484
rect 319404 506472 319410 506524
rect 431954 506472 431960 506524
rect 432012 506512 432018 506524
rect 477494 506512 477500 506524
rect 432012 506484 477500 506512
rect 432012 506472 432018 506484
rect 477494 506472 477500 506484
rect 477552 506472 477558 506524
rect 522942 506472 522948 506524
rect 523000 506512 523006 506524
rect 527818 506512 527824 506524
rect 523000 506484 527824 506512
rect 523000 506472 523006 506484
rect 527818 506472 527824 506484
rect 527876 506472 527882 506524
rect 320266 506404 320272 506456
rect 320324 506444 320330 506456
rect 351178 506444 351184 506456
rect 320324 506416 351184 506444
rect 320324 506404 320330 506416
rect 351178 506404 351184 506416
rect 351236 506404 351242 506456
rect 353110 506404 353116 506456
rect 353168 506444 353174 506456
rect 357434 506444 357440 506456
rect 353168 506416 357440 506444
rect 353168 506404 353174 506416
rect 357434 506404 357440 506416
rect 357492 506404 357498 506456
rect 401594 506404 401600 506456
rect 401652 506444 401658 506456
rect 403342 506444 403348 506456
rect 401652 506416 403348 506444
rect 401652 506404 401658 506416
rect 403342 506404 403348 506416
rect 403400 506404 403406 506456
rect 318978 506336 318984 506388
rect 319036 506376 319042 506388
rect 320082 506376 320088 506388
rect 319036 506348 320088 506376
rect 319036 506336 319042 506348
rect 320082 506336 320088 506348
rect 320140 506376 320146 506388
rect 329742 506376 329748 506388
rect 320140 506348 329748 506376
rect 320140 506336 320146 506348
rect 329742 506336 329748 506348
rect 329800 506336 329806 506388
rect 350166 506336 350172 506388
rect 350224 506376 350230 506388
rect 357618 506376 357624 506388
rect 350224 506348 357624 506376
rect 350224 506336 350230 506348
rect 357618 506336 357624 506348
rect 357676 506336 357682 506388
rect 329742 505724 329748 505776
rect 329800 505764 329806 505776
rect 359274 505764 359280 505776
rect 329800 505736 359280 505764
rect 329800 505724 329806 505736
rect 359274 505724 359280 505736
rect 359332 505724 359338 505776
rect 322566 505248 322572 505300
rect 322624 505288 322630 505300
rect 322750 505288 322756 505300
rect 322624 505260 322756 505288
rect 322624 505248 322630 505260
rect 322750 505248 322756 505260
rect 322808 505248 322814 505300
rect 254302 505112 254308 505164
rect 254360 505152 254366 505164
rect 269942 505152 269948 505164
rect 254360 505124 269948 505152
rect 254360 505112 254366 505124
rect 269942 505112 269948 505124
rect 270000 505112 270006 505164
rect 322474 505044 322480 505096
rect 322532 505084 322538 505096
rect 329190 505084 329196 505096
rect 322532 505056 329196 505084
rect 322532 505044 322538 505056
rect 329190 505044 329196 505056
rect 329248 505044 329254 505096
rect 341518 505044 341524 505096
rect 341576 505084 341582 505096
rect 357434 505084 357440 505096
rect 341576 505056 357440 505084
rect 341576 505044 341582 505056
rect 357434 505044 357440 505056
rect 357492 505044 357498 505096
rect 357618 504364 357624 504416
rect 357676 504404 357682 504416
rect 357894 504404 357900 504416
rect 357676 504376 357900 504404
rect 357676 504364 357682 504376
rect 357894 504364 357900 504376
rect 357952 504364 357958 504416
rect 349062 504160 349068 504212
rect 349120 504200 349126 504212
rect 349982 504200 349988 504212
rect 349120 504172 349988 504200
rect 349120 504160 349126 504172
rect 349982 504160 349988 504172
rect 350040 504160 350046 504212
rect 320266 503820 320272 503872
rect 320324 503860 320330 503872
rect 320542 503860 320548 503872
rect 320324 503832 320548 503860
rect 320324 503820 320330 503832
rect 320542 503820 320548 503832
rect 320600 503820 320606 503872
rect 321554 503684 321560 503736
rect 321612 503724 321618 503736
rect 349062 503724 349068 503736
rect 321612 503696 349068 503724
rect 321612 503684 321618 503696
rect 349062 503684 349068 503696
rect 349120 503684 349126 503736
rect 322474 503616 322480 503668
rect 322532 503656 322538 503668
rect 347130 503656 347136 503668
rect 322532 503628 347136 503656
rect 322532 503616 322538 503628
rect 347130 503616 347136 503628
rect 347188 503616 347194 503668
rect 401594 503616 401600 503668
rect 401652 503656 401658 503668
rect 407114 503656 407120 503668
rect 401652 503628 407120 503656
rect 401652 503616 401658 503628
rect 407114 503616 407120 503628
rect 407172 503616 407178 503668
rect 322658 502936 322664 502988
rect 322716 502976 322722 502988
rect 359366 502976 359372 502988
rect 322716 502948 359372 502976
rect 322716 502936 322722 502948
rect 359366 502936 359372 502948
rect 359424 502936 359430 502988
rect 462958 502324 462964 502376
rect 463016 502364 463022 502376
rect 477494 502364 477500 502376
rect 463016 502336 477500 502364
rect 463016 502324 463022 502336
rect 477494 502324 477500 502336
rect 477552 502324 477558 502376
rect 337378 502256 337384 502308
rect 337436 502296 337442 502308
rect 357434 502296 357440 502308
rect 337436 502268 357440 502296
rect 337436 502256 337442 502268
rect 357434 502256 357440 502268
rect 357492 502256 357498 502308
rect 434714 500964 434720 501016
rect 434772 501004 434778 501016
rect 477494 501004 477500 501016
rect 434772 500976 477500 501004
rect 434772 500964 434778 500976
rect 477494 500964 477500 500976
rect 477552 500964 477558 501016
rect 322566 500896 322572 500948
rect 322624 500936 322630 500948
rect 399570 500936 399576 500948
rect 322624 500908 399576 500936
rect 322624 500896 322630 500908
rect 399570 500896 399576 500908
rect 399628 500896 399634 500948
rect 478782 500896 478788 500948
rect 478840 500936 478846 500948
rect 519722 500936 519728 500948
rect 478840 500908 519728 500936
rect 478840 500896 478846 500908
rect 519722 500896 519728 500908
rect 519780 500896 519786 500948
rect 347038 500828 347044 500880
rect 347096 500868 347102 500880
rect 401962 500868 401968 500880
rect 347096 500840 401968 500868
rect 347096 500828 347102 500840
rect 401962 500828 401968 500840
rect 402020 500828 402026 500880
rect 359274 500760 359280 500812
rect 359332 500800 359338 500812
rect 359918 500800 359924 500812
rect 359332 500772 359924 500800
rect 359332 500760 359338 500772
rect 359918 500760 359924 500772
rect 359976 500760 359982 500812
rect 295242 500352 295248 500404
rect 295300 500392 295306 500404
rect 322934 500392 322940 500404
rect 295300 500364 322940 500392
rect 295300 500352 295306 500364
rect 322934 500352 322940 500364
rect 322992 500352 322998 500404
rect 322474 500284 322480 500336
rect 322532 500324 322538 500336
rect 359734 500324 359740 500336
rect 322532 500296 359740 500324
rect 322532 500284 322538 500296
rect 359734 500284 359740 500296
rect 359792 500284 359798 500336
rect 296622 500216 296628 500268
rect 296680 500256 296686 500268
rect 321738 500256 321744 500268
rect 296680 500228 321744 500256
rect 296680 500216 296686 500228
rect 321738 500216 321744 500228
rect 321796 500216 321802 500268
rect 322750 500216 322756 500268
rect 322808 500256 322814 500268
rect 322808 500228 354674 500256
rect 322808 500216 322814 500228
rect 354646 499984 354674 500228
rect 462314 500216 462320 500268
rect 462372 500256 462378 500268
rect 477402 500256 477408 500268
rect 462372 500228 477408 500256
rect 462372 500216 462378 500228
rect 477402 500216 477408 500228
rect 477460 500216 477466 500268
rect 360470 499984 360476 499996
rect 354646 499956 360476 499984
rect 360470 499944 360476 499956
rect 360528 499944 360534 499996
rect 359734 499876 359740 499928
rect 359792 499916 359798 499928
rect 362954 499916 362960 499928
rect 359792 499888 362960 499916
rect 359792 499876 359798 499888
rect 362954 499876 362960 499888
rect 363012 499916 363018 499928
rect 363874 499916 363880 499928
rect 363012 499888 363880 499916
rect 363012 499876 363018 499888
rect 363874 499876 363880 499888
rect 363932 499876 363938 499928
rect 254578 499536 254584 499588
rect 254636 499576 254642 499588
rect 262858 499576 262864 499588
rect 254636 499548 262864 499576
rect 254636 499536 254642 499548
rect 262858 499536 262864 499548
rect 262916 499536 262922 499588
rect 401594 499536 401600 499588
rect 401652 499576 401658 499588
rect 433334 499576 433340 499588
rect 401652 499548 433340 499576
rect 401652 499536 401658 499548
rect 433334 499536 433340 499548
rect 433392 499536 433398 499588
rect 454678 499536 454684 499588
rect 454736 499576 454742 499588
rect 477494 499576 477500 499588
rect 454736 499548 477500 499576
rect 454736 499536 454742 499548
rect 477494 499536 477500 499548
rect 477552 499536 477558 499588
rect 352926 499468 352932 499520
rect 352984 499508 352990 499520
rect 379330 499508 379336 499520
rect 352984 499480 379336 499508
rect 352984 499468 352990 499480
rect 379330 499468 379336 499480
rect 379388 499468 379394 499520
rect 394142 499468 394148 499520
rect 394200 499508 394206 499520
rect 403710 499508 403716 499520
rect 394200 499480 403716 499508
rect 394200 499468 394206 499480
rect 403710 499468 403716 499480
rect 403768 499468 403774 499520
rect 472710 499468 472716 499520
rect 472768 499508 472774 499520
rect 485774 499508 485780 499520
rect 472768 499480 485780 499508
rect 472768 499468 472774 499480
rect 485774 499468 485780 499480
rect 485832 499468 485838 499520
rect 358906 499400 358912 499452
rect 358964 499440 358970 499452
rect 478414 499440 478420 499452
rect 358964 499412 478420 499440
rect 358964 499400 358970 499412
rect 478414 499400 478420 499412
rect 478472 499400 478478 499452
rect 481358 499400 481364 499452
rect 481416 499440 481422 499452
rect 520826 499440 520832 499452
rect 481416 499412 520832 499440
rect 481416 499400 481422 499412
rect 520826 499400 520832 499412
rect 520884 499400 520890 499452
rect 323670 499332 323676 499384
rect 323728 499372 323734 499384
rect 369670 499372 369676 499384
rect 323728 499344 369676 499372
rect 323728 499332 323734 499344
rect 369670 499332 369676 499344
rect 369728 499332 369734 499384
rect 373534 499332 373540 499384
rect 373592 499372 373598 499384
rect 472802 499372 472808 499384
rect 373592 499344 472808 499372
rect 373592 499332 373598 499344
rect 472802 499332 472808 499344
rect 472860 499332 472866 499384
rect 477678 499332 477684 499384
rect 477736 499372 477742 499384
rect 492214 499372 492220 499384
rect 477736 499344 492220 499372
rect 477736 499332 477742 499344
rect 492214 499332 492220 499344
rect 492272 499332 492278 499384
rect 493594 499332 493600 499384
rect 493652 499372 493658 499384
rect 523678 499372 523684 499384
rect 493652 499344 523684 499372
rect 493652 499332 493658 499344
rect 523678 499332 523684 499344
rect 523736 499332 523742 499384
rect 323578 499264 323584 499316
rect 323636 499304 323642 499316
rect 397362 499304 397368 499316
rect 323636 499276 397368 499304
rect 323636 499264 323642 499276
rect 397362 499264 397368 499276
rect 397420 499264 397426 499316
rect 406470 499264 406476 499316
rect 406528 499304 406534 499316
rect 505738 499304 505744 499316
rect 406528 499276 505744 499304
rect 406528 499264 406534 499276
rect 505738 499264 505744 499276
rect 505796 499264 505802 499316
rect 352834 499196 352840 499248
rect 352892 499236 352898 499248
rect 399478 499236 399484 499248
rect 352892 499208 399484 499236
rect 352892 499196 352898 499208
rect 399478 499196 399484 499208
rect 399536 499196 399542 499248
rect 409230 499196 409236 499248
rect 409288 499236 409294 499248
rect 494790 499236 494796 499248
rect 409288 499208 494796 499236
rect 409288 499196 409294 499208
rect 494790 499196 494796 499208
rect 494848 499196 494854 499248
rect 357158 499128 357164 499180
rect 357216 499168 357222 499180
rect 402330 499168 402336 499180
rect 357216 499140 402336 499168
rect 357216 499128 357222 499140
rect 402330 499128 402336 499140
rect 402388 499128 402394 499180
rect 355410 499060 355416 499112
rect 355468 499100 355474 499112
rect 398006 499100 398012 499112
rect 355468 499072 398012 499100
rect 355468 499060 355474 499072
rect 398006 499060 398012 499072
rect 398064 499060 398070 499112
rect 357250 498992 357256 499044
rect 357308 499032 357314 499044
rect 389634 499032 389640 499044
rect 357308 499004 389640 499032
rect 357308 498992 357314 499004
rect 389634 498992 389640 499004
rect 389692 498992 389698 499044
rect 518250 498992 518256 499044
rect 518308 499032 518314 499044
rect 522390 499032 522396 499044
rect 518308 499004 522396 499032
rect 518308 498992 518314 499004
rect 522390 498992 522396 499004
rect 522448 498992 522454 499044
rect 359918 498924 359924 498976
rect 359976 498964 359982 498976
rect 381906 498964 381912 498976
rect 359976 498936 381912 498964
rect 359976 498924 359982 498936
rect 381906 498924 381912 498936
rect 381964 498924 381970 498976
rect 518158 498924 518164 498976
rect 518216 498964 518222 498976
rect 522482 498964 522488 498976
rect 518216 498936 522488 498964
rect 518216 498924 518222 498936
rect 522482 498924 522488 498936
rect 522540 498924 522546 498976
rect 357342 498856 357348 498908
rect 357400 498896 357406 498908
rect 367094 498896 367100 498908
rect 357400 498868 367100 498896
rect 357400 498856 357406 498868
rect 367094 498856 367100 498868
rect 367152 498856 367158 498908
rect 516778 498856 516784 498908
rect 516836 498896 516842 498908
rect 522298 498896 522304 498908
rect 516836 498868 522304 498896
rect 516836 498856 516842 498868
rect 522298 498856 522304 498868
rect 522356 498856 522362 498908
rect 278774 498788 278780 498840
rect 278832 498828 278838 498840
rect 320634 498828 320640 498840
rect 278832 498800 320640 498828
rect 278832 498788 278838 498800
rect 320634 498788 320640 498800
rect 320692 498788 320698 498840
rect 325050 498788 325056 498840
rect 325108 498828 325114 498840
rect 353478 498828 353484 498840
rect 325108 498800 353484 498828
rect 325108 498788 325114 498800
rect 353478 498788 353484 498800
rect 353536 498828 353542 498840
rect 367738 498828 367744 498840
rect 353536 498800 367744 498828
rect 353536 498788 353542 498800
rect 367738 498788 367744 498800
rect 367796 498788 367802 498840
rect 506474 498788 506480 498840
rect 506532 498828 506538 498840
rect 519814 498828 519820 498840
rect 506532 498800 519820 498828
rect 506532 498788 506538 498800
rect 519814 498788 519820 498800
rect 519872 498788 519878 498840
rect 320910 498720 320916 498772
rect 320968 498760 320974 498772
rect 370314 498760 370320 498772
rect 320968 498732 370320 498760
rect 320968 498720 320974 498732
rect 370314 498720 370320 498732
rect 370372 498720 370378 498772
rect 375466 498720 375472 498772
rect 375524 498760 375530 498772
rect 526438 498760 526444 498772
rect 375524 498732 526444 498760
rect 375524 498720 375530 498732
rect 526438 498720 526444 498732
rect 526496 498720 526502 498772
rect 354214 498176 354220 498228
rect 354272 498216 354278 498228
rect 354272 498188 354674 498216
rect 354272 498176 354278 498188
rect 354646 498080 354674 498188
rect 355410 498176 355416 498228
rect 355468 498216 355474 498228
rect 355594 498216 355600 498228
rect 355468 498188 355600 498216
rect 355468 498176 355474 498188
rect 355594 498176 355600 498188
rect 355652 498176 355658 498228
rect 357066 498108 357072 498160
rect 357124 498148 357130 498160
rect 361942 498148 361948 498160
rect 357124 498120 361948 498148
rect 357124 498108 357130 498120
rect 361942 498108 361948 498120
rect 362000 498108 362006 498160
rect 399294 498108 399300 498160
rect 399352 498148 399358 498160
rect 403894 498148 403900 498160
rect 399352 498120 403900 498148
rect 399352 498108 399358 498120
rect 403894 498108 403900 498120
rect 403952 498108 403958 498160
rect 479518 498108 479524 498160
rect 479576 498148 479582 498160
rect 483842 498148 483848 498160
rect 479576 498120 483848 498148
rect 479576 498108 479582 498120
rect 483842 498108 483848 498120
rect 483900 498108 483906 498160
rect 355410 498080 355416 498092
rect 354646 498052 355416 498080
rect 355410 498040 355416 498052
rect 355468 498080 355474 498092
rect 361298 498080 361304 498092
rect 355468 498052 361304 498080
rect 355468 498040 355474 498052
rect 361298 498040 361304 498052
rect 361356 498040 361362 498092
rect 396718 498040 396724 498092
rect 396776 498080 396782 498092
rect 403158 498080 403164 498092
rect 396776 498052 403164 498080
rect 396776 498040 396782 498052
rect 403158 498040 403164 498052
rect 403216 498040 403222 498092
rect 475562 498040 475568 498092
rect 475620 498080 475626 498092
rect 512178 498080 512184 498092
rect 475620 498052 512184 498080
rect 475620 498040 475626 498052
rect 512178 498040 512184 498052
rect 512236 498040 512242 498092
rect 355962 497972 355968 498024
rect 356020 498012 356026 498024
rect 364518 498012 364524 498024
rect 356020 497984 364524 498012
rect 356020 497972 356026 497984
rect 364518 497972 364524 497984
rect 364576 497972 364582 498024
rect 477034 497972 477040 498024
rect 477092 498012 477098 498024
rect 489638 498012 489644 498024
rect 477092 497984 489644 498012
rect 477092 497972 477098 497984
rect 489638 497972 489644 497984
rect 489696 497972 489702 498024
rect 498838 497972 498844 498024
rect 498896 498012 498902 498024
rect 499298 498012 499304 498024
rect 498896 497984 499304 498012
rect 498896 497972 498902 497984
rect 499298 497972 499304 497984
rect 499356 498012 499362 498024
rect 513466 498012 513472 498024
rect 499356 497984 513472 498012
rect 499356 497972 499362 497984
rect 513466 497972 513472 497984
rect 513524 497972 513530 498024
rect 296530 497904 296536 497956
rect 296588 497944 296594 497956
rect 305546 497944 305552 497956
rect 296588 497916 305552 497944
rect 296588 497904 296594 497916
rect 305546 497904 305552 497916
rect 305604 497904 305610 497956
rect 355502 497904 355508 497956
rect 355560 497944 355566 497956
rect 383838 497944 383844 497956
rect 355560 497916 383844 497944
rect 355560 497904 355566 497916
rect 383838 497904 383844 497916
rect 383896 497904 383902 497956
rect 388346 497904 388352 497956
rect 388404 497944 388410 497956
rect 405182 497944 405188 497956
rect 388404 497916 405188 497944
rect 388404 497904 388410 497916
rect 405182 497904 405188 497916
rect 405240 497904 405246 497956
rect 477402 497904 477408 497956
rect 477460 497944 477466 497956
rect 516042 497944 516048 497956
rect 477460 497916 516048 497944
rect 477460 497904 477466 497916
rect 516042 497904 516048 497916
rect 516100 497904 516106 497956
rect 298738 497836 298744 497888
rect 298796 497876 298802 497888
rect 312170 497876 312176 497888
rect 298796 497848 312176 497876
rect 298796 497836 298802 497848
rect 312170 497836 312176 497848
rect 312228 497836 312234 497888
rect 352558 497836 352564 497888
rect 352616 497876 352622 497888
rect 379974 497876 379980 497888
rect 352616 497848 379980 497876
rect 352616 497836 352622 497848
rect 379974 497836 379980 497848
rect 380032 497836 380038 497888
rect 291930 497768 291936 497820
rect 291988 497808 291994 497820
rect 315114 497808 315120 497820
rect 291988 497780 315120 497808
rect 291988 497768 291994 497780
rect 315114 497768 315120 497780
rect 315172 497768 315178 497820
rect 352466 497768 352472 497820
rect 352524 497808 352530 497820
rect 376110 497808 376116 497820
rect 352524 497780 376116 497808
rect 352524 497768 352530 497780
rect 376110 497768 376116 497780
rect 376168 497768 376174 497820
rect 376386 497768 376392 497820
rect 376444 497808 376450 497820
rect 393498 497808 393504 497820
rect 376444 497780 393504 497808
rect 376444 497768 376450 497780
rect 393498 497768 393504 497780
rect 393556 497768 393562 497820
rect 286042 497700 286048 497752
rect 286100 497740 286106 497752
rect 292022 497740 292028 497752
rect 286100 497712 292028 497740
rect 286100 497700 286106 497712
rect 292022 497700 292028 497712
rect 292080 497700 292086 497752
rect 293218 497700 293224 497752
rect 293276 497740 293282 497752
rect 316034 497740 316040 497752
rect 293276 497712 316040 497740
rect 293276 497700 293282 497712
rect 316034 497700 316040 497712
rect 316092 497700 316098 497752
rect 354122 497700 354128 497752
rect 354180 497740 354186 497752
rect 378042 497740 378048 497752
rect 354180 497712 378048 497740
rect 354180 497700 354186 497712
rect 378042 497700 378048 497712
rect 378100 497700 378106 497752
rect 258810 497632 258816 497684
rect 258868 497672 258874 497684
rect 301866 497672 301872 497684
rect 258868 497644 301872 497672
rect 258868 497632 258874 497644
rect 301866 497632 301872 497644
rect 301924 497632 301930 497684
rect 355318 497632 355324 497684
rect 355376 497672 355382 497684
rect 371602 497672 371608 497684
rect 355376 497644 371608 497672
rect 355376 497632 355382 497644
rect 371602 497632 371608 497644
rect 371660 497632 371666 497684
rect 459554 497632 459560 497684
rect 459612 497672 459618 497684
rect 486418 497672 486424 497684
rect 459612 497644 486424 497672
rect 459612 497632 459618 497644
rect 486418 497632 486424 497644
rect 486476 497632 486482 497684
rect 510338 497632 510344 497684
rect 510396 497672 510402 497684
rect 526438 497672 526444 497684
rect 510396 497644 526444 497672
rect 510396 497632 510402 497644
rect 526438 497632 526444 497644
rect 526496 497632 526502 497684
rect 267090 497564 267096 497616
rect 267148 497604 267154 497616
rect 316586 497604 316592 497616
rect 267148 497576 316592 497604
rect 267148 497564 267154 497576
rect 316586 497564 316592 497576
rect 316644 497564 316650 497616
rect 349062 497564 349068 497616
rect 349120 497604 349126 497616
rect 401686 497604 401692 497616
rect 349120 497576 401692 497604
rect 349120 497564 349126 497576
rect 401686 497564 401692 497576
rect 401744 497564 401750 497616
rect 456794 497564 456800 497616
rect 456852 497604 456858 497616
rect 488994 497604 489000 497616
rect 456852 497576 489000 497604
rect 456852 497564 456858 497576
rect 488994 497564 489000 497576
rect 489052 497564 489058 497616
rect 489178 497564 489184 497616
rect 489236 497604 489242 497616
rect 512822 497604 512828 497616
rect 489236 497576 512828 497604
rect 489236 497564 489242 497576
rect 512822 497564 512828 497576
rect 512880 497564 512886 497616
rect 256142 497496 256148 497548
rect 256200 497536 256206 497548
rect 314654 497536 314660 497548
rect 256200 497508 314660 497536
rect 256200 497496 256206 497508
rect 314654 497496 314660 497508
rect 314712 497496 314718 497548
rect 352742 497496 352748 497548
rect 352800 497536 352806 497548
rect 366450 497536 366456 497548
rect 352800 497508 366456 497536
rect 352800 497496 352806 497508
rect 366450 497496 366456 497508
rect 366508 497496 366514 497548
rect 398834 497496 398840 497548
rect 398892 497536 398898 497548
rect 480622 497536 480628 497548
rect 398892 497508 480628 497536
rect 398892 497496 398898 497508
rect 480622 497496 480628 497508
rect 480680 497496 480686 497548
rect 491938 497496 491944 497548
rect 491996 497536 492002 497548
rect 517330 497536 517336 497548
rect 491996 497508 517336 497536
rect 491996 497496 492002 497508
rect 517330 497496 517336 497508
rect 517388 497496 517394 497548
rect 257614 497428 257620 497480
rect 257672 497468 257678 497480
rect 317414 497468 317420 497480
rect 257672 497440 317420 497468
rect 257672 497428 257678 497440
rect 317414 497428 317420 497440
rect 317472 497428 317478 497480
rect 350074 497428 350080 497480
rect 350132 497468 350138 497480
rect 402054 497468 402060 497480
rect 350132 497440 402060 497468
rect 350132 497428 350138 497440
rect 402054 497428 402060 497440
rect 402112 497428 402118 497480
rect 409874 497428 409880 497480
rect 409932 497468 409938 497480
rect 514754 497468 514760 497480
rect 409932 497440 514760 497468
rect 409932 497428 409938 497440
rect 514754 497428 514760 497440
rect 514812 497428 514818 497480
rect 349890 497360 349896 497412
rect 349948 497400 349954 497412
rect 394786 497400 394792 497412
rect 349948 497372 394792 497400
rect 349948 497360 349954 497372
rect 394786 497360 394792 497372
rect 394844 497360 394850 497412
rect 352650 497292 352656 497344
rect 352708 497332 352714 497344
rect 372246 497332 372252 497344
rect 352708 497304 372252 497332
rect 352708 497292 352714 497304
rect 372246 497292 372252 497304
rect 372304 497292 372310 497344
rect 349798 497224 349804 497276
rect 349856 497264 349862 497276
rect 363230 497264 363236 497276
rect 349856 497236 363236 497264
rect 349856 497224 349862 497236
rect 363230 497224 363236 497236
rect 363288 497224 363294 497276
rect 486418 496816 486424 496868
rect 486476 496856 486482 496868
rect 490926 496856 490932 496868
rect 486476 496828 490932 496856
rect 486476 496816 486482 496828
rect 490926 496816 490932 496828
rect 490984 496816 490990 496868
rect 493318 496816 493324 496868
rect 493376 496856 493382 496868
rect 497366 496856 497372 496868
rect 493376 496828 497372 496856
rect 493376 496816 493382 496828
rect 497366 496816 497372 496828
rect 497424 496816 497430 496868
rect 479058 496748 479064 496800
rect 479116 496788 479122 496800
rect 481634 496788 481640 496800
rect 479116 496760 481640 496788
rect 479116 496748 479122 496760
rect 481634 496748 481640 496760
rect 481692 496748 481698 496800
rect 294138 496340 294144 496392
rect 294196 496380 294202 496392
rect 295978 496380 295984 496392
rect 294196 496352 295984 496380
rect 294196 496340 294202 496352
rect 295978 496340 295984 496352
rect 296036 496340 296042 496392
rect 357526 496340 357532 496392
rect 357584 496380 357590 496392
rect 362218 496380 362224 496392
rect 357584 496352 362224 496380
rect 357584 496340 357590 496352
rect 362218 496340 362224 496352
rect 362276 496340 362282 496392
rect 488442 496340 488448 496392
rect 488500 496380 488506 496392
rect 490558 496380 490564 496392
rect 488500 496352 490564 496380
rect 488500 496340 488506 496352
rect 490558 496340 490564 496352
rect 490616 496340 490622 496392
rect 501322 496204 501328 496256
rect 501380 496244 501386 496256
rect 516870 496244 516876 496256
rect 501380 496216 516876 496244
rect 501380 496204 501386 496216
rect 516870 496204 516876 496216
rect 516928 496204 516934 496256
rect 297266 496136 297272 496188
rect 297324 496176 297330 496188
rect 311894 496176 311900 496188
rect 297324 496148 311900 496176
rect 297324 496136 297330 496148
rect 311894 496136 311900 496148
rect 311952 496136 311958 496188
rect 358170 496136 358176 496188
rect 358228 496176 358234 496188
rect 408494 496176 408500 496188
rect 358228 496148 408500 496176
rect 358228 496136 358234 496148
rect 408494 496136 408500 496148
rect 408552 496136 408558 496188
rect 498194 496136 498200 496188
rect 498252 496176 498258 496188
rect 520090 496176 520096 496188
rect 498252 496148 520096 496176
rect 498252 496136 498258 496148
rect 520090 496136 520096 496148
rect 520148 496136 520154 496188
rect 285674 496068 285680 496120
rect 285732 496108 285738 496120
rect 320358 496108 320364 496120
rect 285732 496080 320364 496108
rect 285732 496068 285738 496080
rect 320358 496068 320364 496080
rect 320416 496068 320422 496120
rect 373994 496068 374000 496120
rect 374052 496108 374058 496120
rect 479702 496108 479708 496120
rect 374052 496080 479708 496108
rect 374052 496068 374058 496080
rect 479702 496068 479708 496080
rect 479760 496068 479766 496120
rect 491294 496068 491300 496120
rect 491352 496108 491358 496120
rect 520918 496108 520924 496120
rect 491352 496080 520924 496108
rect 491352 496068 491358 496080
rect 520918 496068 520924 496080
rect 520976 496068 520982 496120
rect 299382 494980 299388 495032
rect 299440 495020 299446 495032
rect 302326 495020 302332 495032
rect 299440 494992 302332 495020
rect 299440 494980 299446 494992
rect 302326 494980 302332 494992
rect 302384 494980 302390 495032
rect 484394 494776 484400 494828
rect 484452 494816 484458 494828
rect 520366 494816 520372 494828
rect 484452 494788 520372 494816
rect 484452 494776 484458 494788
rect 520366 494776 520372 494788
rect 520424 494776 520430 494828
rect 284294 494708 284300 494760
rect 284352 494748 284358 494760
rect 284938 494748 284944 494760
rect 284352 494720 284944 494748
rect 284352 494708 284358 494720
rect 284938 494708 284944 494720
rect 284996 494708 285002 494760
rect 287054 494708 287060 494760
rect 287112 494748 287118 494760
rect 287882 494748 287888 494760
rect 287112 494720 287888 494748
rect 287112 494708 287118 494720
rect 287882 494708 287888 494720
rect 287940 494708 287946 494760
rect 289814 494708 289820 494760
rect 289872 494748 289878 494760
rect 290826 494748 290832 494760
rect 289872 494720 290832 494748
rect 289872 494708 289878 494720
rect 290826 494708 290832 494720
rect 290884 494708 290890 494760
rect 292574 494708 292580 494760
rect 292632 494748 292638 494760
rect 319070 494748 319076 494760
rect 292632 494720 319076 494748
rect 292632 494708 292638 494720
rect 319070 494708 319076 494720
rect 319128 494708 319134 494760
rect 358354 494708 358360 494760
rect 358412 494748 358418 494760
rect 376018 494748 376024 494760
rect 358412 494720 376024 494748
rect 358412 494708 358418 494720
rect 376018 494708 376024 494720
rect 376076 494708 376082 494760
rect 478506 494708 478512 494760
rect 478564 494748 478570 494760
rect 563054 494748 563060 494760
rect 478564 494720 563060 494748
rect 478564 494708 478570 494720
rect 563054 494708 563060 494720
rect 563112 494708 563118 494760
rect 299474 494640 299480 494692
rect 299532 494680 299538 494692
rect 300394 494680 300400 494692
rect 299532 494652 300400 494680
rect 299532 494640 299538 494652
rect 300394 494640 300400 494652
rect 300452 494640 300458 494692
rect 307754 494096 307760 494148
rect 307812 494136 307818 494148
rect 308490 494136 308496 494148
rect 307812 494108 308496 494136
rect 307812 494096 307818 494108
rect 308490 494096 308496 494108
rect 308548 494096 308554 494148
rect 254578 494028 254584 494080
rect 254636 494068 254642 494080
rect 261570 494068 261576 494080
rect 254636 494040 261576 494068
rect 254636 494028 254642 494040
rect 261570 494028 261576 494040
rect 261628 494028 261634 494080
rect 478966 493484 478972 493536
rect 479024 493524 479030 493536
rect 488534 493524 488540 493536
rect 479024 493496 488540 493524
rect 479024 493484 479030 493496
rect 488534 493484 488540 493496
rect 488592 493484 488598 493536
rect 378686 493416 378692 493468
rect 378744 493456 378750 493468
rect 455414 493456 455420 493468
rect 378744 493428 455420 493456
rect 378744 493416 378750 493428
rect 455414 493416 455420 493428
rect 455472 493416 455478 493468
rect 483290 493416 483296 493468
rect 483348 493456 483354 493468
rect 552014 493456 552020 493468
rect 483348 493428 552020 493456
rect 483348 493416 483354 493428
rect 552014 493416 552020 493428
rect 552072 493416 552078 493468
rect 441614 493348 441620 493400
rect 441672 493388 441678 493400
rect 522206 493388 522212 493400
rect 441672 493360 522212 493388
rect 441672 493348 441678 493360
rect 522206 493348 522212 493360
rect 522264 493348 522270 493400
rect 264974 493280 264980 493332
rect 265032 493320 265038 493332
rect 320450 493320 320456 493332
rect 265032 493292 320456 493320
rect 265032 493280 265038 493292
rect 320450 493280 320456 493292
rect 320508 493280 320514 493332
rect 396074 493280 396080 493332
rect 396132 493320 396138 493332
rect 522022 493320 522028 493332
rect 396132 493292 522028 493320
rect 396132 493280 396138 493292
rect 522022 493280 522028 493292
rect 522080 493280 522086 493332
rect 500218 493008 500224 493060
rect 500276 493048 500282 493060
rect 505094 493048 505100 493060
rect 500276 493020 505100 493048
rect 500276 493008 500282 493020
rect 505094 493008 505100 493020
rect 505152 493008 505158 493060
rect 479242 492056 479248 492108
rect 479300 492096 479306 492108
rect 516134 492096 516140 492108
rect 479300 492068 516140 492096
rect 479300 492056 479306 492068
rect 516134 492056 516140 492068
rect 516192 492056 516198 492108
rect 478598 491988 478604 492040
rect 478656 492028 478662 492040
rect 558178 492028 558184 492040
rect 478656 492000 558184 492028
rect 478656 491988 478662 492000
rect 558178 491988 558184 492000
rect 558236 491988 558242 492040
rect 297358 491920 297364 491972
rect 297416 491960 297422 491972
rect 351914 491960 351920 491972
rect 297416 491932 351920 491960
rect 297416 491920 297422 491932
rect 351914 491920 351920 491932
rect 351972 491920 351978 491972
rect 353294 491920 353300 491972
rect 353352 491960 353358 491972
rect 519630 491960 519636 491972
rect 353352 491932 519636 491960
rect 353352 491920 353358 491932
rect 519630 491920 519636 491932
rect 519688 491920 519694 491972
rect 288434 491512 288440 491564
rect 288492 491552 288498 491564
rect 289354 491552 289360 491564
rect 288492 491524 289360 491552
rect 288492 491512 288498 491524
rect 289354 491512 289360 491524
rect 289412 491512 289418 491564
rect 407114 490560 407120 490612
rect 407172 490600 407178 490612
rect 519998 490600 520004 490612
rect 407172 490572 520004 490600
rect 407172 490560 407178 490572
rect 519998 490560 520004 490572
rect 520056 490560 520062 490612
rect 254578 488520 254584 488572
rect 254636 488560 254642 488572
rect 279510 488560 279516 488572
rect 254636 488532 279516 488560
rect 254636 488520 254642 488532
rect 279510 488520 279516 488532
rect 279568 488520 279574 488572
rect 49602 487840 49608 487892
rect 49660 487880 49666 487892
rect 50338 487880 50344 487892
rect 49660 487852 50344 487880
rect 49660 487840 49666 487852
rect 50338 487840 50344 487852
rect 50396 487840 50402 487892
rect 307846 487840 307852 487892
rect 307904 487880 307910 487892
rect 349706 487880 349712 487892
rect 307904 487852 349712 487880
rect 307904 487840 307910 487852
rect 349706 487840 349712 487852
rect 349764 487840 349770 487892
rect 478690 487840 478696 487892
rect 478748 487880 478754 487892
rect 582374 487880 582380 487892
rect 478748 487852 582380 487880
rect 478748 487840 478754 487852
rect 582374 487840 582380 487852
rect 582432 487840 582438 487892
rect 267734 487772 267740 487824
rect 267792 487812 267798 487824
rect 318978 487812 318984 487824
rect 267792 487784 318984 487812
rect 267792 487772 267798 487784
rect 318978 487772 318984 487784
rect 319036 487772 319042 487824
rect 355502 487772 355508 487824
rect 355560 487812 355566 487824
rect 494146 487812 494152 487824
rect 355560 487784 494152 487812
rect 355560 487772 355566 487784
rect 494146 487772 494152 487784
rect 494204 487772 494210 487824
rect 276014 486412 276020 486464
rect 276072 486452 276078 486464
rect 320266 486452 320272 486464
rect 276072 486424 320272 486452
rect 276072 486412 276078 486424
rect 320266 486412 320272 486424
rect 320324 486412 320330 486464
rect 479334 486412 479340 486464
rect 479392 486452 479398 486464
rect 534074 486452 534080 486464
rect 479392 486424 534080 486452
rect 479392 486412 479398 486424
rect 534074 486412 534080 486424
rect 534132 486412 534138 486464
rect 525150 485732 525156 485784
rect 525208 485772 525214 485784
rect 580166 485772 580172 485784
rect 525208 485744 580172 485772
rect 525208 485732 525214 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 479150 483624 479156 483676
rect 479208 483664 479214 483676
rect 569954 483664 569960 483676
rect 479208 483636 569960 483664
rect 479208 483624 479214 483636
rect 569954 483624 569960 483636
rect 570012 483624 570018 483676
rect 289906 482264 289912 482316
rect 289964 482304 289970 482316
rect 332594 482304 332600 482316
rect 289964 482276 332600 482304
rect 289964 482264 289970 482276
rect 332594 482264 332600 482276
rect 332652 482264 332658 482316
rect 254578 481652 254584 481704
rect 254636 481692 254642 481704
rect 268470 481692 268476 481704
rect 254636 481664 268476 481692
rect 254636 481652 254642 481664
rect 268470 481652 268476 481664
rect 268528 481652 268534 481704
rect 49418 481584 49424 481636
rect 49476 481624 49482 481636
rect 50430 481624 50436 481636
rect 49476 481596 50436 481624
rect 49476 481584 49482 481596
rect 50430 481584 50436 481596
rect 50488 481584 50494 481636
rect 364334 480904 364340 480956
rect 364392 480944 364398 480956
rect 460198 480944 460204 480956
rect 364392 480916 460204 480944
rect 364392 480904 364398 480916
rect 460198 480904 460204 480916
rect 460256 480904 460262 480956
rect 389174 479476 389180 479528
rect 389232 479516 389238 479528
rect 515398 479516 515404 479528
rect 389232 479488 515404 479516
rect 389232 479476 389238 479488
rect 515398 479476 515404 479488
rect 515456 479476 515462 479528
rect 371234 478116 371240 478168
rect 371292 478156 371298 478168
rect 503898 478156 503904 478168
rect 371292 478128 503904 478156
rect 371292 478116 371298 478128
rect 503898 478116 503904 478128
rect 503956 478116 503962 478168
rect 254210 476076 254216 476128
rect 254268 476116 254274 476128
rect 265710 476116 265716 476128
rect 254268 476088 265716 476116
rect 254268 476076 254274 476088
rect 265710 476076 265716 476088
rect 265768 476076 265774 476128
rect 363598 475328 363604 475380
rect 363656 475368 363662 475380
rect 481910 475368 481916 475380
rect 363656 475340 481916 475368
rect 363656 475328 363662 475340
rect 481910 475328 481916 475340
rect 481968 475328 481974 475380
rect 46382 473288 46388 473340
rect 46440 473328 46446 473340
rect 48958 473328 48964 473340
rect 46440 473300 48964 473328
rect 46440 473288 46446 473300
rect 48958 473288 48964 473300
rect 49016 473288 49022 473340
rect 338758 471928 338764 471980
rect 338816 471968 338822 471980
rect 580166 471968 580172 471980
rect 338816 471940 580172 471968
rect 338816 471928 338822 471940
rect 580166 471928 580172 471940
rect 580224 471928 580230 471980
rect 254578 470568 254584 470620
rect 254636 470608 254642 470620
rect 264330 470608 264336 470620
rect 254636 470580 264336 470608
rect 254636 470568 254642 470580
rect 264330 470568 264336 470580
rect 264388 470568 264394 470620
rect 45462 467780 45468 467832
rect 45520 467820 45526 467832
rect 48774 467820 48780 467832
rect 45520 467792 48780 467820
rect 45520 467780 45526 467792
rect 48774 467780 48780 467792
rect 48832 467820 48838 467832
rect 49050 467820 49056 467832
rect 48832 467792 49056 467820
rect 48832 467780 48838 467792
rect 49050 467780 49056 467792
rect 49108 467780 49114 467832
rect 254578 465060 254584 465112
rect 254636 465100 254642 465112
rect 271322 465100 271328 465112
rect 254636 465072 271328 465100
rect 254636 465060 254642 465072
rect 271322 465060 271328 465072
rect 271380 465060 271386 465112
rect 46474 462272 46480 462324
rect 46532 462312 46538 462324
rect 50798 462312 50804 462324
rect 46532 462284 50804 462312
rect 46532 462272 46538 462284
rect 50798 462272 50804 462284
rect 50856 462272 50862 462324
rect 254578 458192 254584 458244
rect 254636 458232 254642 458244
rect 278222 458232 278228 458244
rect 254636 458204 278228 458232
rect 254636 458192 254642 458204
rect 278222 458192 278228 458204
rect 278280 458192 278286 458244
rect 359826 458124 359832 458176
rect 359884 458164 359890 458176
rect 580166 458164 580172 458176
rect 359884 458136 580172 458164
rect 359884 458124 359890 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 46566 456356 46572 456408
rect 46624 456396 46630 456408
rect 49786 456396 49792 456408
rect 46624 456368 49792 456396
rect 46624 456356 46630 456368
rect 49786 456356 49792 456368
rect 49844 456356 49850 456408
rect 299566 453976 299572 454028
rect 299624 454016 299630 454028
rect 300946 454016 300952 454028
rect 299624 453988 300952 454016
rect 299624 453976 299630 453988
rect 300946 453976 300952 453988
rect 301004 453976 301010 454028
rect 254302 452616 254308 452668
rect 254360 452656 254366 452668
rect 289078 452656 289084 452668
rect 254360 452628 289084 452656
rect 254360 452616 254366 452628
rect 289078 452616 289084 452628
rect 289136 452616 289142 452668
rect 254670 447108 254676 447160
rect 254728 447148 254734 447160
rect 275462 447148 275468 447160
rect 254728 447120 275468 447148
rect 254728 447108 254734 447120
rect 275462 447108 275468 447120
rect 275520 447108 275526 447160
rect 46658 445680 46664 445732
rect 46716 445720 46722 445732
rect 48314 445720 48320 445732
rect 46716 445692 48320 445720
rect 46716 445680 46722 445692
rect 48314 445680 48320 445692
rect 48372 445680 48378 445732
rect 254394 441736 254400 441788
rect 254452 441776 254458 441788
rect 257522 441776 257528 441788
rect 254452 441748 257528 441776
rect 254452 441736 254458 441748
rect 257522 441736 257528 441748
rect 257580 441736 257586 441788
rect 46750 438812 46756 438864
rect 46808 438852 46814 438864
rect 48314 438852 48320 438864
rect 46808 438824 48320 438852
rect 46808 438812 46814 438824
rect 48314 438812 48320 438824
rect 48372 438812 48378 438864
rect 254394 434732 254400 434784
rect 254452 434772 254458 434784
rect 291838 434772 291844 434784
rect 254452 434744 291844 434772
rect 254452 434732 254458 434744
rect 291838 434732 291844 434744
rect 291896 434732 291902 434784
rect 46842 433236 46848 433288
rect 46900 433276 46906 433288
rect 49142 433276 49148 433288
rect 46900 433248 49148 433276
rect 46900 433236 46906 433248
rect 49142 433236 49148 433248
rect 49200 433236 49206 433288
rect 477862 431876 477868 431928
rect 477920 431916 477926 431928
rect 579798 431916 579804 431928
rect 477920 431888 579804 431916
rect 477920 431876 477926 431888
rect 579798 431876 579804 431888
rect 579856 431876 579862 431928
rect 254578 429156 254584 429208
rect 254636 429196 254642 429208
rect 350902 429196 350908 429208
rect 254636 429168 350908 429196
rect 254636 429156 254642 429168
rect 350902 429156 350908 429168
rect 350960 429156 350966 429208
rect 254578 423648 254584 423700
rect 254636 423688 254642 423700
rect 323578 423688 323584 423700
rect 254636 423660 323584 423688
rect 254636 423648 254642 423660
rect 323578 423648 323584 423660
rect 323636 423648 323642 423700
rect 324958 419432 324964 419484
rect 325016 419472 325022 419484
rect 580166 419472 580172 419484
rect 325016 419444 580172 419472
rect 325016 419432 325022 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 254578 418140 254584 418192
rect 254636 418180 254642 418192
rect 282178 418180 282184 418192
rect 254636 418152 282184 418180
rect 254636 418140 254642 418152
rect 282178 418140 282184 418152
rect 282236 418140 282242 418192
rect 254578 411272 254584 411324
rect 254636 411312 254642 411324
rect 349982 411312 349988 411324
rect 254636 411284 349988 411312
rect 254636 411272 254642 411284
rect 349982 411272 349988 411284
rect 350040 411272 350046 411324
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 50522 409884 50528 409896
rect 3200 409856 50528 409884
rect 3200 409844 3206 409856
rect 50522 409844 50528 409856
rect 50580 409844 50586 409896
rect 376018 405628 376024 405680
rect 376076 405668 376082 405680
rect 580166 405668 580172 405680
rect 376076 405640 580172 405668
rect 376076 405628 376082 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 254026 400188 254032 400240
rect 254084 400228 254090 400240
rect 350810 400228 350816 400240
rect 254084 400200 350816 400228
rect 254084 400188 254090 400200
rect 350810 400188 350816 400200
rect 350868 400188 350874 400240
rect 46842 397468 46848 397520
rect 46900 397508 46906 397520
rect 49418 397508 49424 397520
rect 46900 397480 49424 397508
rect 46900 397468 46906 397480
rect 49418 397468 49424 397480
rect 49476 397468 49482 397520
rect 254670 394748 254676 394800
rect 254728 394788 254734 394800
rect 260282 394788 260288 394800
rect 254728 394760 260288 394788
rect 254728 394748 254734 394760
rect 260282 394748 260288 394760
rect 260340 394748 260346 394800
rect 46750 391960 46756 392012
rect 46808 392000 46814 392012
rect 48314 392000 48320 392012
rect 46808 391972 48320 392000
rect 46808 391960 46814 391972
rect 48314 391960 48320 391972
rect 48372 391960 48378 392012
rect 254670 389172 254676 389224
rect 254728 389212 254734 389224
rect 317414 389212 317420 389224
rect 254728 389184 317420 389212
rect 254728 389172 254734 389184
rect 317414 389172 317420 389184
rect 317472 389172 317478 389224
rect 46658 385024 46664 385076
rect 46716 385064 46722 385076
rect 48314 385064 48320 385076
rect 46716 385036 48320 385064
rect 46716 385024 46722 385036
rect 48314 385024 48320 385036
rect 48372 385024 48378 385076
rect 254394 382236 254400 382288
rect 254452 382276 254458 382288
rect 289170 382276 289176 382288
rect 254452 382248 289176 382276
rect 254452 382236 254458 382248
rect 289170 382236 289176 382248
rect 289228 382236 289234 382288
rect 46566 379516 46572 379568
rect 46624 379556 46630 379568
rect 49418 379556 49424 379568
rect 46624 379528 49424 379556
rect 46624 379516 46630 379528
rect 49418 379516 49424 379528
rect 49476 379516 49482 379568
rect 544378 379448 544384 379500
rect 544436 379488 544442 379500
rect 580166 379488 580172 379500
rect 544436 379460 580172 379488
rect 544436 379448 544442 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 254118 376728 254124 376780
rect 254176 376768 254182 376780
rect 351086 376768 351092 376780
rect 254176 376740 351092 376768
rect 254176 376728 254182 376740
rect 351086 376728 351092 376740
rect 351144 376728 351150 376780
rect 254670 371220 254676 371272
rect 254728 371260 254734 371272
rect 301498 371260 301504 371272
rect 254728 371232 301504 371260
rect 254728 371220 254734 371232
rect 301498 371220 301504 371232
rect 301556 371220 301562 371272
rect 281534 369112 281540 369164
rect 281592 369152 281598 369164
rect 283558 369152 283564 369164
rect 281592 369124 283564 369152
rect 281592 369112 281598 369124
rect 283558 369112 283564 369124
rect 283616 369112 283622 369164
rect 254670 365712 254676 365764
rect 254728 365752 254734 365764
rect 282270 365752 282276 365764
rect 254728 365724 282276 365752
rect 254728 365712 254734 365724
rect 282270 365712 282276 365724
rect 282328 365712 282334 365764
rect 320818 365644 320824 365696
rect 320876 365684 320882 365696
rect 580166 365684 580172 365696
rect 320876 365656 580172 365684
rect 320876 365644 320882 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 253934 358844 253940 358896
rect 253992 358884 253998 358896
rect 256234 358884 256240 358896
rect 253992 358856 256240 358884
rect 253992 358844 253998 358856
rect 256234 358844 256240 358856
rect 256292 358844 256298 358896
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 50614 357456 50620 357468
rect 3200 357428 50620 357456
rect 3200 357416 3206 357428
rect 50614 357416 50620 357428
rect 50672 357416 50678 357468
rect 288526 353948 288532 354000
rect 288584 353988 288590 354000
rect 352190 353988 352196 354000
rect 288584 353960 352196 353988
rect 288584 353948 288590 353960
rect 352190 353948 352196 353960
rect 352248 353948 352254 354000
rect 498746 353948 498752 354000
rect 498804 353988 498810 354000
rect 540974 353988 540980 354000
rect 498804 353960 540980 353988
rect 498804 353948 498810 353960
rect 540974 353948 540980 353960
rect 541032 353948 541038 354000
rect 254210 353268 254216 353320
rect 254268 353308 254274 353320
rect 289262 353308 289268 353320
rect 254268 353280 289268 353308
rect 254268 353268 254274 353280
rect 289262 353268 289268 353280
rect 289320 353268 289326 353320
rect 362218 353200 362224 353252
rect 362276 353240 362282 353252
rect 580166 353240 580172 353252
rect 362276 353212 580172 353240
rect 362276 353200 362282 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 385034 352520 385040 352572
rect 385092 352560 385098 352572
rect 521930 352560 521936 352572
rect 385092 352532 521936 352560
rect 385092 352520 385098 352532
rect 521930 352520 521936 352532
rect 521988 352520 521994 352572
rect 297634 351228 297640 351280
rect 297692 351268 297698 351280
rect 313366 351268 313372 351280
rect 297692 351240 313372 351268
rect 297692 351228 297698 351240
rect 313366 351228 313372 351240
rect 313424 351228 313430 351280
rect 298002 351160 298008 351212
rect 298060 351200 298066 351212
rect 320174 351200 320180 351212
rect 298060 351172 320180 351200
rect 298060 351160 298066 351172
rect 320174 351160 320180 351172
rect 320232 351160 320238 351212
rect 287146 349800 287152 349852
rect 287204 349840 287210 349852
rect 350074 349840 350080 349852
rect 287204 349812 350080 349840
rect 287204 349800 287210 349812
rect 350074 349800 350080 349812
rect 350132 349800 350138 349852
rect 254486 347760 254492 347812
rect 254544 347800 254550 347812
rect 346486 347800 346492 347812
rect 254544 347772 346492 347800
rect 254544 347760 254550 347772
rect 346486 347760 346492 347772
rect 346544 347760 346550 347812
rect 299658 345652 299664 345704
rect 299716 345692 299722 345704
rect 314654 345692 314660 345704
rect 299716 345664 314660 345692
rect 299716 345652 299722 345664
rect 314654 345652 314660 345664
rect 314712 345652 314718 345704
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 50246 345080 50252 345092
rect 3384 345052 50252 345080
rect 3384 345040 3390 345052
rect 50246 345040 50252 345052
rect 50304 345040 50310 345092
rect 284386 344292 284392 344344
rect 284444 344332 284450 344344
rect 352006 344332 352012 344344
rect 284444 344304 352012 344332
rect 284444 344292 284450 344304
rect 352006 344292 352012 344304
rect 352064 344292 352070 344344
rect 254578 342864 254584 342916
rect 254636 342904 254642 342916
rect 351362 342904 351368 342916
rect 254636 342876 351368 342904
rect 254636 342864 254642 342876
rect 351362 342864 351368 342876
rect 351420 342864 351426 342916
rect 254578 342252 254584 342304
rect 254636 342292 254642 342304
rect 287698 342292 287704 342304
rect 254636 342264 287704 342292
rect 254636 342252 254642 342264
rect 287698 342252 287704 342264
rect 287756 342252 287762 342304
rect 296990 341572 296996 341624
rect 297048 341612 297054 341624
rect 311986 341612 311992 341624
rect 297048 341584 311992 341612
rect 297048 341572 297054 341584
rect 311986 341572 311992 341584
rect 312044 341572 312050 341624
rect 289814 341504 289820 341556
rect 289872 341544 289878 341556
rect 349798 341544 349804 341556
rect 289872 341516 349804 341544
rect 289872 341504 289878 341516
rect 349798 341504 349804 341516
rect 349856 341504 349862 341556
rect 271874 340212 271880 340264
rect 271932 340252 271938 340264
rect 318886 340252 318892 340264
rect 271932 340224 318892 340252
rect 271932 340212 271938 340224
rect 318886 340212 318892 340224
rect 318944 340212 318950 340264
rect 285766 340144 285772 340196
rect 285824 340184 285830 340196
rect 352282 340184 352288 340196
rect 285824 340156 352288 340184
rect 285824 340144 285830 340156
rect 352282 340144 352288 340156
rect 352340 340144 352346 340196
rect 282914 338784 282920 338836
rect 282972 338824 282978 338836
rect 318794 338824 318800 338836
rect 282972 338796 318800 338824
rect 282972 338784 282978 338796
rect 318794 338784 318800 338796
rect 318852 338784 318858 338836
rect 310606 338716 310612 338768
rect 310664 338756 310670 338768
rect 350258 338756 350264 338768
rect 310664 338728 350264 338756
rect 310664 338716 310670 338728
rect 350258 338716 350264 338728
rect 350316 338716 350322 338768
rect 289814 337424 289820 337476
rect 289872 337464 289878 337476
rect 322290 337464 322296 337476
rect 289872 337436 322296 337464
rect 289872 337424 289878 337436
rect 322290 337424 322296 337436
rect 322348 337424 322354 337476
rect 288434 337356 288440 337408
rect 288492 337396 288498 337408
rect 352098 337396 352104 337408
rect 288492 337368 352104 337396
rect 288492 337356 288498 337368
rect 352098 337356 352104 337368
rect 352156 337356 352162 337408
rect 299474 335996 299480 336048
rect 299532 336036 299538 336048
rect 319346 336036 319352 336048
rect 299532 336008 319352 336036
rect 299532 335996 299538 336008
rect 319346 335996 319352 336008
rect 319404 335996 319410 336048
rect 254394 335316 254400 335368
rect 254452 335356 254458 335368
rect 332226 335356 332232 335368
rect 254452 335328 332232 335356
rect 254452 335316 254458 335328
rect 332226 335316 332232 335328
rect 332284 335316 332290 335368
rect 310514 334704 310520 334756
rect 310572 334744 310578 334756
rect 352558 334744 352564 334756
rect 310572 334716 352564 334744
rect 310572 334704 310578 334716
rect 352558 334704 352564 334716
rect 352616 334704 352622 334756
rect 291286 334636 291292 334688
rect 291344 334676 291350 334688
rect 351270 334676 351276 334688
rect 291344 334648 351276 334676
rect 291344 334636 291350 334648
rect 351270 334636 351276 334648
rect 351328 334636 351334 334688
rect 260834 334568 260840 334620
rect 260892 334608 260898 334620
rect 321554 334608 321560 334620
rect 260892 334580 321560 334608
rect 260892 334568 260898 334580
rect 321554 334568 321560 334580
rect 321612 334568 321618 334620
rect 298646 333344 298652 333396
rect 298704 333384 298710 333396
rect 307754 333384 307760 333396
rect 298704 333356 307760 333384
rect 298704 333344 298710 333356
rect 307754 333344 307760 333356
rect 307812 333344 307818 333396
rect 306466 333276 306472 333328
rect 306524 333316 306530 333328
rect 352466 333316 352472 333328
rect 306524 333288 352472 333316
rect 306524 333276 306530 333288
rect 352466 333276 352472 333288
rect 352524 333276 352530 333328
rect 283098 333208 283104 333260
rect 283156 333248 283162 333260
rect 350166 333248 350172 333260
rect 283156 333220 350172 333248
rect 283156 333208 283162 333220
rect 350166 333208 350172 333220
rect 350224 333208 350230 333260
rect 301498 332936 301504 332988
rect 301556 332976 301562 332988
rect 306466 332976 306472 332988
rect 301556 332948 306472 332976
rect 301556 332936 301562 332948
rect 306466 332936 306472 332948
rect 306524 332936 306530 332988
rect 297910 332596 297916 332648
rect 297968 332636 297974 332648
rect 298094 332636 298100 332648
rect 297968 332608 298100 332636
rect 297968 332596 297974 332608
rect 298094 332596 298100 332608
rect 298152 332596 298158 332648
rect 299750 332528 299756 332580
rect 299808 332568 299814 332580
rect 306374 332568 306380 332580
rect 299808 332540 306380 332568
rect 299808 332528 299814 332540
rect 306374 332528 306380 332540
rect 306432 332528 306438 332580
rect 323578 332324 323584 332376
rect 323636 332364 323642 332376
rect 325142 332364 325148 332376
rect 323636 332336 325148 332364
rect 323636 332324 323642 332336
rect 325142 332324 325148 332336
rect 325200 332324 325206 332376
rect 298830 332256 298836 332308
rect 298888 332296 298894 332308
rect 347682 332296 347688 332308
rect 298888 332268 347688 332296
rect 298888 332256 298894 332268
rect 347682 332256 347688 332268
rect 347740 332256 347746 332308
rect 294598 332188 294604 332240
rect 294656 332228 294662 332240
rect 310330 332228 310336 332240
rect 294656 332200 310336 332228
rect 294656 332188 294662 332200
rect 310330 332188 310336 332200
rect 310388 332188 310394 332240
rect 296254 332052 296260 332104
rect 296312 332092 296318 332104
rect 309226 332092 309232 332104
rect 296312 332064 309232 332092
rect 296312 332052 296318 332064
rect 309226 332052 309232 332064
rect 309284 332052 309290 332104
rect 303798 331984 303804 332036
rect 303856 332024 303862 332036
rect 320634 332024 320640 332036
rect 303856 331996 320640 332024
rect 303856 331984 303862 331996
rect 320634 331984 320640 331996
rect 320692 331984 320698 332036
rect 294966 331916 294972 331968
rect 295024 331956 295030 331968
rect 305086 331956 305092 331968
rect 295024 331928 305092 331956
rect 295024 331916 295030 331928
rect 305086 331916 305092 331928
rect 305144 331916 305150 331968
rect 309134 331916 309140 331968
rect 309192 331956 309198 331968
rect 353754 331956 353760 331968
rect 309192 331928 353760 331956
rect 309192 331916 309198 331928
rect 353754 331916 353760 331928
rect 353812 331916 353818 331968
rect 295058 331848 295064 331900
rect 295116 331888 295122 331900
rect 302418 331888 302424 331900
rect 295116 331860 302424 331888
rect 295116 331848 295122 331860
rect 302418 331848 302424 331860
rect 302476 331848 302482 331900
rect 303614 331848 303620 331900
rect 303672 331888 303678 331900
rect 353846 331888 353852 331900
rect 303672 331860 353852 331888
rect 303672 331848 303678 331860
rect 353846 331848 353852 331860
rect 353904 331848 353910 331900
rect 285030 331780 285036 331832
rect 285088 331820 285094 331832
rect 321922 331820 321928 331832
rect 285088 331792 321928 331820
rect 285088 331780 285094 331792
rect 321922 331780 321928 331792
rect 321980 331780 321986 331832
rect 296346 331712 296352 331764
rect 296404 331752 296410 331764
rect 309042 331752 309048 331764
rect 296404 331724 309048 331752
rect 296404 331712 296410 331724
rect 309042 331712 309048 331724
rect 309100 331712 309106 331764
rect 253290 331644 253296 331696
rect 253348 331684 253354 331696
rect 341886 331684 341892 331696
rect 253348 331656 341892 331684
rect 253348 331644 253354 331656
rect 341886 331644 341892 331656
rect 341944 331644 341950 331696
rect 294874 331576 294880 331628
rect 294932 331616 294938 331628
rect 313550 331616 313556 331628
rect 294932 331588 313556 331616
rect 294932 331576 294938 331588
rect 313550 331576 313556 331588
rect 313608 331576 313614 331628
rect 296438 331508 296444 331560
rect 296496 331548 296502 331560
rect 330938 331548 330944 331560
rect 296496 331520 330944 331548
rect 296496 331508 296502 331520
rect 330938 331508 330944 331520
rect 330996 331508 331002 331560
rect 339310 331508 339316 331560
rect 339368 331548 339374 331560
rect 354122 331548 354128 331560
rect 339368 331520 354128 331548
rect 339368 331508 339374 331520
rect 354122 331508 354128 331520
rect 354180 331508 354186 331560
rect 287790 331440 287796 331492
rect 287848 331480 287854 331492
rect 323210 331480 323216 331492
rect 287848 331452 323216 331480
rect 287848 331440 287854 331452
rect 323210 331440 323216 331452
rect 323268 331440 323274 331492
rect 336090 331440 336096 331492
rect 336148 331480 336154 331492
rect 352650 331480 352656 331492
rect 336148 331452 352656 331480
rect 336148 331440 336154 331452
rect 352650 331440 352656 331452
rect 352708 331440 352714 331492
rect 298554 331372 298560 331424
rect 298612 331412 298618 331424
rect 307754 331412 307760 331424
rect 298612 331384 307760 331412
rect 298612 331372 298618 331384
rect 307754 331372 307760 331384
rect 307812 331372 307818 331424
rect 327718 331372 327724 331424
rect 327776 331412 327782 331424
rect 352742 331412 352748 331424
rect 327776 331384 352748 331412
rect 327776 331372 327782 331384
rect 352742 331372 352748 331384
rect 352800 331372 352806 331424
rect 253198 331304 253204 331356
rect 253256 331344 253262 331356
rect 300670 331344 300676 331356
rect 253256 331316 300676 331344
rect 253256 331304 253262 331316
rect 300670 331304 300676 331316
rect 300728 331304 300734 331356
rect 338022 331304 338028 331356
rect 338080 331344 338086 331356
rect 353662 331344 353668 331356
rect 338080 331316 353668 331344
rect 338080 331304 338086 331316
rect 353662 331304 353668 331316
rect 353720 331304 353726 331356
rect 295150 331236 295156 331288
rect 295208 331276 295214 331288
rect 301958 331276 301964 331288
rect 295208 331248 301964 331276
rect 295208 331236 295214 331248
rect 301958 331236 301964 331248
rect 302016 331236 302022 331288
rect 345106 331236 345112 331288
rect 345164 331276 345170 331288
rect 349890 331276 349896 331288
rect 345164 331248 349896 331276
rect 345164 331236 345170 331248
rect 349890 331236 349896 331248
rect 349948 331236 349954 331288
rect 299014 330148 299020 330200
rect 299072 330188 299078 330200
rect 326430 330188 326436 330200
rect 299072 330160 326436 330188
rect 299072 330148 299078 330160
rect 326430 330148 326436 330160
rect 326488 330148 326494 330200
rect 299106 330080 299112 330132
rect 299164 330120 299170 330132
rect 329006 330120 329012 330132
rect 299164 330092 329012 330120
rect 299164 330080 299170 330092
rect 329006 330080 329012 330092
rect 329064 330080 329070 330132
rect 299198 330012 299204 330064
rect 299256 330052 299262 330064
rect 334526 330052 334532 330064
rect 299256 330024 334532 330052
rect 299256 330012 299262 330024
rect 334526 330012 334532 330024
rect 334584 330012 334590 330064
rect 298922 329944 298928 329996
rect 298980 329984 298986 329996
rect 340230 329984 340236 329996
rect 298980 329956 340236 329984
rect 298980 329944 298986 329956
rect 340230 329944 340236 329956
rect 340288 329944 340294 329996
rect 254210 329876 254216 329928
rect 254268 329916 254274 329928
rect 284938 329916 284944 329928
rect 254268 329888 284944 329916
rect 254268 329876 254274 329888
rect 284938 329876 284944 329888
rect 284996 329876 285002 329928
rect 299290 329876 299296 329928
rect 299348 329916 299354 329928
rect 343634 329916 343640 329928
rect 299348 329888 343640 329916
rect 299348 329876 299354 329888
rect 343634 329876 343640 329888
rect 343692 329876 343698 329928
rect 254670 329808 254676 329860
rect 254728 329848 254734 329860
rect 351454 329848 351460 329860
rect 254728 329820 351460 329848
rect 254728 329808 254734 329820
rect 351454 329808 351460 329820
rect 351512 329808 351518 329860
rect 254486 325592 254492 325644
rect 254544 325632 254550 325644
rect 285030 325632 285036 325644
rect 254544 325604 285036 325632
rect 254544 325592 254550 325604
rect 285030 325592 285036 325604
rect 285088 325592 285094 325644
rect 490558 325592 490564 325644
rect 490616 325632 490622 325644
rect 580166 325632 580172 325644
rect 490616 325604 580172 325632
rect 490616 325592 490622 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 283558 324232 283564 324284
rect 283616 324272 283622 324284
rect 297818 324272 297824 324284
rect 283616 324244 297824 324272
rect 283616 324232 283622 324244
rect 297818 324232 297824 324244
rect 297876 324232 297882 324284
rect 254302 320084 254308 320136
rect 254360 320124 254366 320136
rect 287790 320124 287796 320136
rect 254360 320096 287796 320124
rect 254360 320084 254366 320096
rect 287790 320084 287796 320096
rect 287848 320084 287854 320136
rect 282270 318724 282276 318776
rect 282328 318764 282334 318776
rect 297726 318764 297732 318776
rect 282328 318736 297732 318764
rect 282328 318724 282334 318736
rect 297726 318724 297732 318736
rect 297784 318724 297790 318776
rect 349798 318724 349804 318776
rect 349856 318764 349862 318776
rect 349856 318736 350028 318764
rect 349856 318724 349862 318736
rect 350000 318708 350028 318736
rect 349982 318656 349988 318708
rect 350040 318656 350046 318708
rect 284938 317364 284944 317416
rect 284996 317404 285002 317416
rect 297726 317404 297732 317416
rect 284996 317376 297732 317404
rect 284996 317364 285002 317376
rect 297726 317364 297732 317376
rect 297784 317364 297790 317416
rect 292758 313216 292764 313268
rect 292816 313256 292822 313268
rect 297910 313256 297916 313268
rect 292816 313228 297916 313256
rect 292816 313216 292822 313228
rect 297910 313216 297916 313228
rect 297968 313216 297974 313268
rect 356974 313216 356980 313268
rect 357032 313256 357038 313268
rect 580166 313256 580172 313268
rect 357032 313228 580172 313256
rect 357032 313216 357038 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 349982 312168 349988 312180
rect 349816 312140 349988 312168
rect 349816 312112 349844 312140
rect 349982 312128 349988 312140
rect 350040 312128 350046 312180
rect 349798 312060 349804 312112
rect 349856 312060 349862 312112
rect 297910 311040 297916 311092
rect 297968 311080 297974 311092
rect 298738 311080 298744 311092
rect 297968 311052 298744 311080
rect 297968 311040 297974 311052
rect 298738 311040 298744 311052
rect 298796 311040 298802 311092
rect 351178 310564 351184 310616
rect 351236 310604 351242 310616
rect 351914 310604 351920 310616
rect 351236 310576 351920 310604
rect 351236 310564 351242 310576
rect 351914 310564 351920 310576
rect 351972 310564 351978 310616
rect 350258 309068 350264 309120
rect 350316 309108 350322 309120
rect 351914 309108 351920 309120
rect 350316 309080 351920 309108
rect 350316 309068 350322 309080
rect 351914 309068 351920 309080
rect 351972 309068 351978 309120
rect 260282 307708 260288 307760
rect 260340 307748 260346 307760
rect 297266 307748 297272 307760
rect 260340 307720 297272 307748
rect 260340 307708 260346 307720
rect 297266 307708 297272 307720
rect 297324 307708 297330 307760
rect 254210 306348 254216 306400
rect 254268 306388 254274 306400
rect 293310 306388 293316 306400
rect 254268 306360 293316 306388
rect 254268 306348 254274 306360
rect 293310 306348 293316 306360
rect 293368 306348 293374 306400
rect 256234 306280 256240 306332
rect 256292 306320 256298 306332
rect 298002 306320 298008 306332
rect 256292 306292 298008 306320
rect 256292 306280 256298 306292
rect 298002 306280 298008 306292
rect 298060 306280 298066 306332
rect 293954 303560 293960 303612
rect 294012 303600 294018 303612
rect 298002 303600 298008 303612
rect 294012 303572 298008 303600
rect 294012 303560 294018 303572
rect 298002 303560 298008 303572
rect 298060 303560 298066 303612
rect 254670 300840 254676 300892
rect 254728 300880 254734 300892
rect 294690 300880 294696 300892
rect 254728 300852 294696 300880
rect 254728 300840 254734 300852
rect 294690 300840 294696 300852
rect 294748 300840 294754 300892
rect 383194 299412 383200 299464
rect 383252 299452 383258 299464
rect 580166 299452 580172 299464
rect 383252 299424 580172 299452
rect 383252 299412 383258 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 254670 295332 254676 295384
rect 254728 295372 254734 295384
rect 284938 295372 284944 295384
rect 254728 295344 284944 295372
rect 254728 295332 254734 295344
rect 284938 295332 284944 295344
rect 284996 295332 285002 295384
rect 297818 295128 297824 295180
rect 297876 295168 297882 295180
rect 299842 295168 299848 295180
rect 297876 295140 299848 295168
rect 297876 295128 297882 295140
rect 299842 295128 299848 295140
rect 299900 295128 299906 295180
rect 284294 292476 284300 292528
rect 284352 292516 284358 292528
rect 298002 292516 298008 292528
rect 284352 292488 298008 292516
rect 284352 292476 284358 292488
rect 298002 292476 298008 292488
rect 298060 292476 298066 292528
rect 351362 291660 351368 291712
rect 351420 291700 351426 291712
rect 353570 291700 353576 291712
rect 351420 291672 353576 291700
rect 351420 291660 351426 291672
rect 353570 291660 353576 291672
rect 353628 291660 353634 291712
rect 295426 289416 295432 289468
rect 295484 289456 295490 289468
rect 298002 289456 298008 289468
rect 295484 289428 298008 289456
rect 295484 289416 295490 289428
rect 298002 289416 298008 289428
rect 298060 289416 298066 289468
rect 254394 288396 254400 288448
rect 254452 288436 254458 288448
rect 296162 288436 296168 288448
rect 254452 288408 296168 288436
rect 254452 288396 254458 288408
rect 296162 288396 296168 288408
rect 296220 288396 296226 288448
rect 292022 288328 292028 288380
rect 292080 288368 292086 288380
rect 298002 288368 298008 288380
rect 292080 288340 298008 288368
rect 292080 288328 292086 288340
rect 298002 288328 298008 288340
rect 298060 288328 298066 288380
rect 297818 287376 297824 287428
rect 297876 287376 297882 287428
rect 297836 287088 297864 287376
rect 297818 287036 297824 287088
rect 297876 287036 297882 287088
rect 297818 285880 297824 285932
rect 297876 285880 297882 285932
rect 297836 285728 297864 285880
rect 297818 285676 297824 285728
rect 297876 285676 297882 285728
rect 289170 285608 289176 285660
rect 289228 285648 289234 285660
rect 297910 285648 297916 285660
rect 289228 285620 297916 285648
rect 289228 285608 289234 285620
rect 297910 285608 297916 285620
rect 297968 285608 297974 285660
rect 254302 282888 254308 282940
rect 254360 282928 254366 282940
rect 264422 282928 264428 282940
rect 254360 282900 264428 282928
rect 254360 282888 254366 282900
rect 264422 282888 264428 282900
rect 264480 282888 264486 282940
rect 50614 282004 50620 282056
rect 50672 282044 50678 282056
rect 298094 282044 298100 282056
rect 50672 282016 298100 282044
rect 50672 282004 50678 282016
rect 298094 282004 298100 282016
rect 298152 282004 298158 282056
rect 46658 281936 46664 281988
rect 46716 281976 46722 281988
rect 279786 281976 279792 281988
rect 46716 281948 279792 281976
rect 46716 281936 46722 281948
rect 279786 281936 279792 281948
rect 279844 281936 279850 281988
rect 49142 281868 49148 281920
rect 49200 281908 49206 281920
rect 278314 281908 278320 281920
rect 49200 281880 278320 281908
rect 49200 281868 49206 281880
rect 278314 281868 278320 281880
rect 278372 281868 278378 281920
rect 3510 281460 3516 281512
rect 3568 281500 3574 281512
rect 519538 281500 519544 281512
rect 3568 281472 519544 281500
rect 3568 281460 3574 281472
rect 519538 281460 519544 281472
rect 519596 281460 519602 281512
rect 3418 281392 3424 281444
rect 3476 281432 3482 281444
rect 485774 281432 485780 281444
rect 3476 281404 485780 281432
rect 3476 281392 3482 281404
rect 485774 281392 485780 281404
rect 485832 281392 485838 281444
rect 50522 281324 50528 281376
rect 50580 281364 50586 281376
rect 521838 281364 521844 281376
rect 50580 281336 521844 281364
rect 50580 281324 50586 281336
rect 521838 281324 521844 281336
rect 521896 281324 521902 281376
rect 48958 281256 48964 281308
rect 49016 281296 49022 281308
rect 53098 281296 53104 281308
rect 49016 281268 53104 281296
rect 49016 281256 49022 281268
rect 53098 281256 53104 281268
rect 53156 281256 53162 281308
rect 284938 281256 284944 281308
rect 284996 281296 285002 281308
rect 352006 281296 352012 281308
rect 284996 281268 352012 281296
rect 284996 281256 285002 281268
rect 352006 281256 352012 281268
rect 352064 281256 352070 281308
rect 49050 281188 49056 281240
rect 49108 281228 49114 281240
rect 54478 281228 54484 281240
rect 49108 281200 54484 281228
rect 49108 281188 49114 281200
rect 54478 281188 54484 281200
rect 54536 281188 54542 281240
rect 54570 281188 54576 281240
rect 54628 281228 54634 281240
rect 279694 281228 279700 281240
rect 54628 281200 279700 281228
rect 54628 281188 54634 281200
rect 279694 281188 279700 281200
rect 279752 281188 279758 281240
rect 52086 281120 52092 281172
rect 52144 281160 52150 281172
rect 280982 281160 280988 281172
rect 52144 281132 280988 281160
rect 52144 281120 52150 281132
rect 280982 281120 280988 281132
rect 281040 281120 281046 281172
rect 48682 281052 48688 281104
rect 48740 281092 48746 281104
rect 280798 281092 280804 281104
rect 48740 281064 280804 281092
rect 48740 281052 48746 281064
rect 280798 281052 280804 281064
rect 280856 281052 280862 281104
rect 49234 280984 49240 281036
rect 49292 281024 49298 281036
rect 276658 281024 276664 281036
rect 49292 280996 276664 281024
rect 49292 280984 49298 280996
rect 276658 280984 276664 280996
rect 276716 280984 276722 281036
rect 48038 280916 48044 280968
rect 48096 280956 48102 280968
rect 54570 280956 54576 280968
rect 48096 280928 54576 280956
rect 48096 280916 48102 280928
rect 54570 280916 54576 280928
rect 54628 280916 54634 280968
rect 272518 280956 272524 280968
rect 55186 280928 272524 280956
rect 48774 280848 48780 280900
rect 48832 280888 48838 280900
rect 55186 280888 55214 280928
rect 272518 280916 272524 280928
rect 272576 280916 272582 280968
rect 48832 280860 55214 280888
rect 48832 280848 48838 280860
rect 49326 280712 49332 280764
rect 49384 280752 49390 280764
rect 287330 280752 287336 280764
rect 49384 280724 287336 280752
rect 49384 280712 49390 280724
rect 287330 280712 287336 280724
rect 287388 280712 287394 280764
rect 297726 280576 297732 280628
rect 297784 280616 297790 280628
rect 300118 280616 300124 280628
rect 297784 280588 300124 280616
rect 297784 280576 297790 280588
rect 300118 280576 300124 280588
rect 300176 280576 300182 280628
rect 3602 280100 3608 280152
rect 3660 280140 3666 280152
rect 468570 280140 468576 280152
rect 3660 280112 468576 280140
rect 3660 280100 3666 280112
rect 468570 280100 468576 280112
rect 468628 280100 468634 280152
rect 50246 280032 50252 280084
rect 50304 280072 50310 280084
rect 507670 280072 507676 280084
rect 50304 280044 507676 280072
rect 50304 280032 50310 280044
rect 507670 280032 507676 280044
rect 507728 280032 507734 280084
rect 48222 279964 48228 280016
rect 48280 280004 48286 280016
rect 279602 280004 279608 280016
rect 48280 279976 279608 280004
rect 48280 279964 48286 279976
rect 279602 279964 279608 279976
rect 279660 279964 279666 280016
rect 296162 279964 296168 280016
rect 296220 280004 296226 280016
rect 351914 280004 351920 280016
rect 296220 279976 351920 280004
rect 296220 279964 296226 279976
rect 351914 279964 351920 279976
rect 351972 279964 351978 280016
rect 298554 279896 298560 279948
rect 298612 279936 298618 279948
rect 303798 279936 303804 279948
rect 298612 279908 303804 279936
rect 298612 279896 298618 279908
rect 303798 279896 303804 279908
rect 303856 279896 303862 279948
rect 294874 279420 294880 279472
rect 294932 279460 294938 279472
rect 310514 279460 310520 279472
rect 294932 279432 310520 279460
rect 294932 279420 294938 279432
rect 310514 279420 310520 279432
rect 310572 279420 310578 279472
rect 321646 279420 321652 279472
rect 321704 279460 321710 279472
rect 354122 279460 354128 279472
rect 321704 279432 354128 279460
rect 321704 279420 321710 279432
rect 354122 279420 354128 279432
rect 354180 279420 354186 279472
rect 289262 279012 289268 279064
rect 289320 279052 289326 279064
rect 315482 279052 315488 279064
rect 289320 279024 315488 279052
rect 289320 279012 289326 279024
rect 315482 279012 315488 279024
rect 315540 279012 315546 279064
rect 282270 278944 282276 278996
rect 282328 278984 282334 278996
rect 321278 278984 321284 278996
rect 282328 278956 321284 278984
rect 282328 278944 282334 278956
rect 321278 278944 321284 278956
rect 321336 278944 321342 278996
rect 287698 278876 287704 278928
rect 287756 278916 287762 278928
rect 330938 278916 330944 278928
rect 287756 278888 330944 278916
rect 287756 278876 287762 278888
rect 330938 278876 330944 278888
rect 330996 278876 331002 278928
rect 294690 278808 294696 278860
rect 294748 278848 294754 278860
rect 342530 278848 342536 278860
rect 294748 278820 342536 278848
rect 294748 278808 294754 278820
rect 342530 278808 342536 278820
rect 342588 278808 342594 278860
rect 293310 278740 293316 278792
rect 293368 278780 293374 278792
rect 349614 278780 349620 278792
rect 293368 278752 349620 278780
rect 293368 278740 293374 278752
rect 349614 278740 349620 278752
rect 349672 278740 349678 278792
rect 295978 278672 295984 278724
rect 296036 278712 296042 278724
rect 301314 278712 301320 278724
rect 296036 278684 301320 278712
rect 296036 278672 296042 278684
rect 301314 278672 301320 278684
rect 301372 278672 301378 278724
rect 308398 278672 308404 278724
rect 308456 278712 308462 278724
rect 313366 278712 313372 278724
rect 308456 278684 313372 278712
rect 308456 278672 308462 278684
rect 313366 278672 313372 278684
rect 313424 278672 313430 278724
rect 316770 278672 316776 278724
rect 316828 278712 316834 278724
rect 323118 278712 323124 278724
rect 316828 278684 323124 278712
rect 316828 278672 316834 278684
rect 323118 278672 323124 278684
rect 323176 278672 323182 278724
rect 347038 278672 347044 278724
rect 347096 278712 347102 278724
rect 353846 278712 353852 278724
rect 347096 278684 353852 278712
rect 347096 278672 347102 278684
rect 353846 278672 353852 278684
rect 353904 278672 353910 278724
rect 296530 278604 296536 278656
rect 296588 278644 296594 278656
rect 305178 278644 305184 278656
rect 296588 278616 305184 278644
rect 296588 278604 296594 278616
rect 305178 278604 305184 278616
rect 305236 278604 305242 278656
rect 339954 278604 339960 278656
rect 340012 278644 340018 278656
rect 353754 278644 353760 278656
rect 340012 278616 353760 278644
rect 340012 278604 340018 278616
rect 353754 278604 353760 278616
rect 353812 278604 353818 278656
rect 295334 278536 295340 278588
rect 295392 278576 295398 278588
rect 335446 278576 335452 278588
rect 295392 278548 335452 278576
rect 295392 278536 295398 278548
rect 335446 278536 335452 278548
rect 335504 278536 335510 278588
rect 292666 278468 292672 278520
rect 292724 278508 292730 278520
rect 319990 278508 319996 278520
rect 292724 278480 319996 278508
rect 292724 278468 292730 278480
rect 319990 278468 319996 278480
rect 320048 278468 320054 278520
rect 296254 278400 296260 278452
rect 296312 278440 296318 278452
rect 322566 278440 322572 278452
rect 296312 278412 322572 278440
rect 296312 278400 296318 278412
rect 322566 278400 322572 278412
rect 322624 278400 322630 278452
rect 299750 278332 299756 278384
rect 299808 278372 299814 278384
rect 318058 278372 318064 278384
rect 299808 278344 318064 278372
rect 299808 278332 299814 278344
rect 318058 278332 318064 278344
rect 318116 278332 318122 278384
rect 337378 278332 337384 278384
rect 337436 278372 337442 278384
rect 341242 278372 341248 278384
rect 337436 278344 341248 278372
rect 337436 278332 337442 278344
rect 341242 278332 341248 278344
rect 341300 278332 341306 278384
rect 287054 278264 287060 278316
rect 287112 278304 287118 278316
rect 303890 278304 303896 278316
rect 287112 278276 303896 278304
rect 287112 278264 287118 278276
rect 303890 278264 303896 278276
rect 303948 278264 303954 278316
rect 294966 278196 294972 278248
rect 295024 278236 295030 278248
rect 338022 278236 338028 278248
rect 295024 278208 338028 278236
rect 295024 278196 295030 278208
rect 338022 278196 338028 278208
rect 338080 278196 338086 278248
rect 298738 278128 298744 278180
rect 298796 278168 298802 278180
rect 303706 278168 303712 278180
rect 298796 278140 303712 278168
rect 298796 278128 298802 278140
rect 303706 278128 303712 278140
rect 303764 278128 303770 278180
rect 334158 278060 334164 278112
rect 334216 278100 334222 278112
rect 338206 278100 338212 278112
rect 334216 278072 338212 278100
rect 334216 278060 334222 278072
rect 338206 278060 338212 278072
rect 338264 278060 338270 278112
rect 59446 277992 59452 278044
rect 59504 278032 59510 278044
rect 297358 278032 297364 278044
rect 59504 278004 297364 278032
rect 59504 277992 59510 278004
rect 297358 277992 297364 278004
rect 297416 277992 297422 278044
rect 317414 277992 317420 278044
rect 317472 278032 317478 278044
rect 343818 278032 343824 278044
rect 317472 278004 343824 278032
rect 317472 277992 317478 278004
rect 343818 277992 343824 278004
rect 343876 277992 343882 278044
rect 295058 277924 295064 277976
rect 295116 277964 295122 277976
rect 345750 277964 345756 277976
rect 295116 277936 345756 277964
rect 295116 277924 295122 277936
rect 345750 277924 345756 277936
rect 345808 277924 345814 277976
rect 300026 277584 300032 277636
rect 300084 277624 300090 277636
rect 305638 277624 305644 277636
rect 300084 277596 305644 277624
rect 300084 277584 300090 277596
rect 305638 277584 305644 277596
rect 305696 277584 305702 277636
rect 323854 277516 323860 277568
rect 323912 277556 323918 277568
rect 326338 277556 326344 277568
rect 323912 277528 326344 277556
rect 323912 277516 323918 277528
rect 326338 277516 326344 277528
rect 326396 277516 326402 277568
rect 324314 277380 324320 277432
rect 324372 277420 324378 277432
rect 327074 277420 327080 277432
rect 324372 277392 327080 277420
rect 324372 277380 324378 277392
rect 327074 277380 327080 277392
rect 327132 277380 327138 277432
rect 297450 276768 297456 276820
rect 297508 276808 297514 276820
rect 309134 276808 309140 276820
rect 297508 276780 309140 276808
rect 297508 276768 297514 276780
rect 309134 276768 309140 276780
rect 309192 276768 309198 276820
rect 314746 276768 314752 276820
rect 314804 276808 314810 276820
rect 351086 276808 351092 276820
rect 314804 276780 351092 276808
rect 314804 276768 314810 276780
rect 351086 276768 351092 276780
rect 351144 276768 351150 276820
rect 59262 276700 59268 276752
rect 59320 276740 59326 276752
rect 352098 276740 352104 276752
rect 59320 276712 352104 276740
rect 59320 276700 59326 276712
rect 352098 276700 352104 276712
rect 352156 276700 352162 276752
rect 3418 276632 3424 276684
rect 3476 276672 3482 276684
rect 519446 276672 519452 276684
rect 3476 276644 519452 276672
rect 3476 276632 3482 276644
rect 519446 276632 519452 276644
rect 519504 276632 519510 276684
rect 299658 276088 299664 276140
rect 299716 276128 299722 276140
rect 304994 276128 305000 276140
rect 299716 276100 305000 276128
rect 299716 276088 299722 276100
rect 304994 276088 305000 276100
rect 305052 276088 305058 276140
rect 297634 276020 297640 276072
rect 297692 276060 297698 276072
rect 298830 276060 298836 276072
rect 297692 276032 298836 276060
rect 297692 276020 297698 276032
rect 298830 276020 298836 276032
rect 298888 276020 298894 276072
rect 297174 275340 297180 275392
rect 297232 275380 297238 275392
rect 311158 275380 311164 275392
rect 297232 275352 311164 275380
rect 297232 275340 297238 275352
rect 311158 275340 311164 275352
rect 311216 275340 311222 275392
rect 7558 275272 7564 275324
rect 7616 275312 7622 275324
rect 501874 275312 501880 275324
rect 7616 275284 501880 275312
rect 7616 275272 7622 275284
rect 501874 275272 501880 275284
rect 501932 275272 501938 275324
rect 297542 273980 297548 274032
rect 297600 274020 297606 274032
rect 335354 274020 335360 274032
rect 297600 273992 335360 274020
rect 297600 273980 297606 273992
rect 335354 273980 335360 273992
rect 335412 273980 335418 274032
rect 3694 273912 3700 273964
rect 3752 273952 3758 273964
rect 520734 273952 520740 273964
rect 3752 273924 520740 273952
rect 3752 273912 3758 273924
rect 520734 273912 520740 273924
rect 520792 273912 520798 273964
rect 499942 273164 499948 273216
rect 500000 273204 500006 273216
rect 580166 273204 580172 273216
rect 500000 273176 580172 273204
rect 500000 273164 500006 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 333974 272620 333980 272672
rect 334032 272660 334038 272672
rect 349798 272660 349804 272672
rect 334032 272632 349804 272660
rect 334032 272620 334038 272632
rect 349798 272620 349804 272632
rect 349856 272620 349862 272672
rect 58894 272552 58900 272604
rect 58952 272592 58958 272604
rect 352374 272592 352380 272604
rect 58952 272564 352380 272592
rect 58952 272552 58958 272564
rect 352374 272552 352380 272564
rect 352432 272552 352438 272604
rect 4798 272484 4804 272536
rect 4856 272524 4862 272536
rect 496722 272524 496728 272536
rect 4856 272496 496728 272524
rect 4856 272484 4862 272496
rect 496722 272484 496728 272496
rect 496780 272484 496786 272536
rect 299566 271124 299572 271176
rect 299624 271164 299630 271176
rect 318794 271164 318800 271176
rect 299624 271136 318800 271164
rect 299624 271124 299630 271136
rect 318794 271124 318800 271136
rect 318852 271124 318858 271176
rect 9674 268336 9680 268388
rect 9732 268376 9738 268388
rect 478230 268376 478236 268388
rect 9732 268348 478236 268376
rect 9732 268336 9738 268348
rect 478230 268336 478236 268348
rect 478288 268336 478294 268388
rect 13814 266976 13820 267028
rect 13872 267016 13878 267028
rect 457438 267016 457444 267028
rect 13872 266988 457444 267016
rect 13872 266976 13878 266988
rect 457438 266976 457444 266988
rect 457496 266976 457502 267028
rect 318886 260108 318892 260160
rect 318944 260148 318950 260160
rect 350994 260148 351000 260160
rect 318944 260120 351000 260148
rect 318944 260108 318950 260120
rect 350994 260108 351000 260120
rect 351052 260108 351058 260160
rect 301498 258680 301504 258732
rect 301556 258720 301562 258732
rect 350902 258720 350908 258732
rect 301556 258692 350908 258720
rect 301556 258680 301562 258692
rect 350902 258680 350908 258692
rect 350960 258680 350966 258732
rect 302326 257320 302332 257372
rect 302384 257360 302390 257372
rect 384482 257360 384488 257372
rect 302384 257332 384488 257360
rect 302384 257320 302390 257332
rect 384482 257320 384488 257332
rect 384540 257320 384546 257372
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 436830 255252 436836 255264
rect 3200 255224 436836 255252
rect 3200 255212 3206 255224
rect 436830 255212 436836 255224
rect 436888 255212 436894 255264
rect 59078 253172 59084 253224
rect 59136 253212 59142 253224
rect 347774 253212 347780 253224
rect 59136 253184 347780 253212
rect 59136 253172 59142 253184
rect 347774 253172 347780 253184
rect 347832 253172 347838 253224
rect 359642 245556 359648 245608
rect 359700 245596 359706 245608
rect 580166 245596 580172 245608
rect 359700 245568 580172 245596
rect 359700 245556 359706 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 423030 241448 423036 241460
rect 3568 241420 423036 241448
rect 3568 241408 3574 241420
rect 423030 241408 423036 241420
rect 423088 241408 423094 241460
rect 58986 236648 58992 236700
rect 59044 236688 59050 236700
rect 352282 236688 352288 236700
rect 59044 236660 352288 236688
rect 59044 236648 59050 236660
rect 352282 236648 352288 236660
rect 352340 236648 352346 236700
rect 59630 235220 59636 235272
rect 59688 235260 59694 235272
rect 311894 235260 311900 235272
rect 59688 235232 311900 235260
rect 59688 235220 59694 235232
rect 311894 235220 311900 235232
rect 311952 235220 311958 235272
rect 58802 233860 58808 233912
rect 58860 233900 58866 233912
rect 310606 233900 310612 233912
rect 58860 233872 310612 233900
rect 58860 233860 58866 233872
rect 310606 233860 310612 233872
rect 310664 233860 310670 233912
rect 534718 233180 534724 233232
rect 534776 233220 534782 233232
rect 579982 233220 579988 233232
rect 534776 233192 579988 233220
rect 534776 233180 534782 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 8938 231072 8944 231124
rect 8996 231112 9002 231124
rect 487062 231112 487068 231124
rect 8996 231084 487068 231112
rect 8996 231072 9002 231084
rect 487062 231072 487068 231084
rect 487120 231072 487126 231124
rect 59998 229712 60004 229764
rect 60056 229752 60062 229764
rect 507118 229752 507124 229764
rect 60056 229724 507124 229752
rect 60056 229712 60062 229724
rect 507118 229712 507124 229724
rect 507176 229712 507182 229764
rect 57330 228420 57336 228472
rect 57388 228460 57394 228472
rect 256142 228460 256148 228472
rect 57388 228432 256148 228460
rect 57388 228420 57394 228432
rect 256142 228420 256148 228432
rect 256200 228420 256206 228472
rect 59538 228352 59544 228404
rect 59596 228392 59602 228404
rect 324406 228392 324412 228404
rect 59596 228364 324412 228392
rect 59596 228352 59602 228364
rect 324406 228352 324412 228364
rect 324464 228352 324470 228404
rect 326062 228352 326068 228404
rect 326120 228392 326126 228404
rect 349706 228392 349712 228404
rect 326120 228364 349712 228392
rect 326120 228352 326126 228364
rect 349706 228352 349712 228364
rect 349764 228352 349770 228404
rect 31018 226992 31024 227044
rect 31076 227032 31082 227044
rect 478138 227032 478144 227044
rect 31076 227004 478144 227032
rect 31076 226992 31082 227004
rect 478138 226992 478144 227004
rect 478196 226992 478202 227044
rect 59170 225632 59176 225684
rect 59228 225672 59234 225684
rect 283190 225672 283196 225684
rect 59228 225644 283196 225672
rect 59228 225632 59234 225644
rect 283190 225632 283196 225644
rect 283248 225632 283254 225684
rect 57790 225564 57796 225616
rect 57848 225604 57854 225616
rect 296070 225604 296076 225616
rect 57848 225576 296076 225604
rect 57848 225564 57854 225576
rect 296070 225564 296076 225576
rect 296128 225564 296134 225616
rect 308858 225564 308864 225616
rect 308916 225604 308922 225616
rect 332594 225604 332600 225616
rect 308916 225576 332600 225604
rect 308916 225564 308922 225576
rect 332594 225564 332600 225576
rect 332652 225564 332658 225616
rect 318794 224272 318800 224324
rect 318852 224312 318858 224324
rect 319622 224312 319628 224324
rect 318852 224284 319628 224312
rect 318852 224272 318858 224284
rect 319622 224272 319628 224284
rect 319680 224272 319686 224324
rect 3786 224204 3792 224256
rect 3844 224244 3850 224256
rect 454770 224244 454776 224256
rect 3844 224216 454776 224244
rect 3844 224204 3850 224216
rect 454770 224204 454776 224216
rect 454828 224204 454834 224256
rect 305638 223524 305644 223576
rect 305696 223564 305702 223576
rect 307846 223564 307852 223576
rect 305696 223536 307852 223564
rect 305696 223524 305702 223536
rect 307846 223524 307852 223536
rect 307904 223524 307910 223576
rect 299934 223456 299940 223508
rect 299992 223496 299998 223508
rect 306834 223496 306840 223508
rect 299992 223468 306840 223496
rect 299992 223456 299998 223468
rect 306834 223456 306840 223468
rect 306892 223456 306898 223508
rect 302234 223184 302240 223236
rect 302292 223224 302298 223236
rect 314930 223224 314936 223236
rect 302292 223196 314936 223224
rect 302292 223184 302298 223196
rect 314930 223184 314936 223196
rect 314988 223184 314994 223236
rect 329098 223184 329104 223236
rect 329156 223224 329162 223236
rect 329156 223196 335354 223224
rect 329156 223184 329162 223196
rect 309226 223116 309232 223168
rect 309284 223156 309290 223168
rect 323026 223156 323032 223168
rect 309284 223128 323032 223156
rect 309284 223116 309290 223128
rect 323026 223116 323032 223128
rect 323084 223116 323090 223168
rect 328086 223116 328092 223168
rect 328144 223156 328150 223168
rect 335326 223156 335354 223196
rect 337194 223184 337200 223236
rect 337252 223224 337258 223236
rect 350074 223224 350080 223236
rect 337252 223196 350080 223224
rect 337252 223184 337258 223196
rect 350074 223184 350080 223196
rect 350132 223184 350138 223236
rect 352650 223156 352656 223168
rect 328144 223128 333284 223156
rect 335326 223128 352656 223156
rect 328144 223116 328150 223128
rect 296346 223048 296352 223100
rect 296404 223088 296410 223100
rect 296404 223060 325694 223088
rect 296404 223048 296410 223060
rect 299842 222980 299848 223032
rect 299900 223020 299906 223032
rect 321002 223020 321008 223032
rect 299900 222992 321008 223020
rect 299900 222980 299906 222992
rect 321002 222980 321008 222992
rect 321060 222980 321066 223032
rect 325666 223020 325694 223060
rect 326338 223048 326344 223100
rect 326396 223088 326402 223100
rect 333146 223088 333152 223100
rect 326396 223060 333152 223088
rect 326396 223048 326402 223060
rect 333146 223048 333152 223060
rect 333204 223048 333210 223100
rect 331122 223020 331128 223032
rect 325666 222992 331128 223020
rect 331122 222980 331128 222992
rect 331180 222980 331186 223032
rect 333256 223020 333284 223128
rect 352650 223116 352656 223128
rect 352708 223116 352714 223168
rect 334158 223048 334164 223100
rect 334216 223088 334222 223100
rect 349890 223088 349896 223100
rect 334216 223060 349896 223088
rect 334216 223048 334222 223060
rect 349890 223048 349896 223060
rect 349948 223048 349954 223100
rect 353662 223020 353668 223032
rect 333256 222992 353668 223020
rect 353662 222980 353668 222992
rect 353720 222980 353726 223032
rect 57514 222912 57520 222964
rect 57572 222952 57578 222964
rect 253290 222952 253296 222964
rect 57572 222924 253296 222952
rect 57572 222912 57578 222924
rect 253290 222912 253296 222924
rect 253348 222912 253354 222964
rect 295150 222912 295156 222964
rect 295208 222952 295214 222964
rect 330110 222952 330116 222964
rect 295208 222924 330116 222952
rect 295208 222912 295214 222924
rect 330110 222912 330116 222924
rect 330168 222912 330174 222964
rect 332134 222912 332140 222964
rect 332192 222952 332198 222964
rect 352742 222952 352748 222964
rect 332192 222924 352748 222952
rect 332192 222912 332198 222924
rect 352742 222912 352748 222924
rect 352800 222912 352806 222964
rect 57054 222844 57060 222896
rect 57112 222884 57118 222896
rect 267090 222884 267096 222896
rect 57112 222856 267096 222884
rect 57112 222844 57118 222856
rect 267090 222844 267096 222856
rect 267148 222844 267154 222896
rect 296438 222844 296444 222896
rect 296496 222884 296502 222896
rect 296496 222856 296714 222884
rect 296496 222844 296502 222856
rect 296686 222816 296714 222856
rect 311158 222844 311164 222896
rect 311216 222884 311222 222896
rect 312906 222884 312912 222896
rect 311216 222856 312912 222884
rect 311216 222844 311222 222856
rect 312906 222844 312912 222856
rect 312964 222844 312970 222896
rect 316954 222844 316960 222896
rect 317012 222884 317018 222896
rect 351178 222884 351184 222896
rect 317012 222856 351184 222884
rect 317012 222844 317018 222856
rect 351178 222844 351184 222856
rect 351236 222844 351242 222896
rect 311894 222816 311900 222828
rect 296686 222788 311900 222816
rect 311894 222776 311900 222788
rect 311952 222776 311958 222828
rect 222838 222232 222844 222284
rect 222896 222272 222902 222284
rect 301498 222272 301504 222284
rect 222896 222244 301504 222272
rect 222896 222232 222902 222244
rect 301498 222232 301504 222244
rect 301556 222232 301562 222284
rect 224402 222164 224408 222216
rect 224460 222204 224466 222216
rect 339218 222204 339224 222216
rect 224460 222176 339224 222204
rect 224460 222164 224466 222176
rect 339218 222164 339224 222176
rect 339276 222164 339282 222216
rect 299474 222096 299480 222148
rect 299532 222136 299538 222148
rect 300762 222136 300768 222148
rect 299532 222108 300768 222136
rect 299532 222096 299538 222108
rect 300762 222096 300768 222108
rect 300820 222096 300826 222148
rect 297358 221552 297364 221604
rect 297416 221592 297422 221604
rect 336918 221592 336924 221604
rect 297416 221564 336924 221592
rect 297416 221552 297422 221564
rect 336918 221552 336924 221564
rect 336976 221552 336982 221604
rect 57238 221484 57244 221536
rect 57296 221524 57302 221536
rect 254578 221524 254584 221536
rect 57296 221496 254584 221524
rect 57296 221484 57302 221496
rect 254578 221484 254584 221496
rect 254636 221484 254642 221536
rect 297450 221484 297456 221536
rect 297508 221524 297514 221536
rect 337378 221524 337384 221536
rect 297508 221496 337384 221524
rect 297508 221484 297514 221496
rect 337378 221484 337384 221496
rect 337436 221484 337442 221536
rect 58710 221416 58716 221468
rect 58768 221456 58774 221468
rect 352834 221456 352840 221468
rect 58768 221428 352840 221456
rect 58768 221416 58774 221428
rect 352834 221416 352840 221428
rect 352892 221416 352898 221468
rect 226058 220804 226064 220856
rect 226116 220844 226122 220856
rect 300762 220844 300768 220856
rect 226116 220816 300768 220844
rect 226116 220804 226122 220816
rect 300762 220804 300768 220816
rect 300820 220844 300826 220856
rect 578878 220844 578884 220856
rect 300820 220816 578884 220844
rect 300820 220804 300826 220816
rect 578878 220804 578884 220816
rect 578936 220804 578942 220856
rect 299382 220260 299388 220312
rect 299440 220300 299446 220312
rect 306374 220300 306380 220312
rect 299440 220272 306380 220300
rect 299440 220260 299446 220272
rect 306374 220260 306380 220272
rect 306432 220260 306438 220312
rect 57146 220192 57152 220244
rect 57204 220232 57210 220244
rect 291930 220232 291936 220244
rect 57204 220204 291936 220232
rect 57204 220192 57210 220204
rect 291930 220192 291936 220204
rect 291988 220192 291994 220244
rect 298830 220192 298836 220244
rect 298888 220232 298894 220244
rect 313274 220232 313280 220244
rect 298888 220204 313280 220232
rect 298888 220192 298894 220204
rect 313274 220192 313280 220204
rect 313332 220192 313338 220244
rect 60550 220124 60556 220176
rect 60608 220164 60614 220176
rect 293218 220164 293224 220176
rect 60608 220136 293224 220164
rect 60608 220124 60614 220136
rect 293218 220124 293224 220136
rect 293276 220124 293282 220176
rect 298738 220124 298744 220176
rect 298796 220164 298802 220176
rect 328454 220164 328460 220176
rect 298796 220136 328460 220164
rect 298796 220124 298802 220136
rect 328454 220124 328460 220136
rect 328512 220124 328518 220176
rect 3602 220056 3608 220108
rect 3660 220096 3666 220108
rect 520642 220096 520648 220108
rect 3660 220068 520648 220096
rect 3660 220056 3666 220068
rect 520642 220056 520648 220068
rect 520700 220056 520706 220108
rect 57882 218832 57888 218884
rect 57940 218872 57946 218884
rect 253198 218872 253204 218884
rect 57940 218844 253204 218872
rect 57940 218832 57946 218844
rect 253198 218832 253204 218844
rect 253256 218832 253262 218884
rect 57422 218764 57428 218816
rect 57480 218804 57486 218816
rect 258810 218804 258816 218816
rect 57480 218776 258816 218804
rect 57480 218764 57486 218776
rect 258810 218764 258816 218776
rect 258868 218764 258874 218816
rect 57606 218696 57612 218748
rect 57664 218736 57670 218748
rect 294598 218736 294604 218748
rect 57664 218708 294604 218736
rect 57664 218696 57670 218708
rect 294598 218696 294604 218708
rect 294656 218696 294662 218748
rect 222930 216656 222936 216708
rect 222988 216696 222994 216708
rect 297910 216696 297916 216708
rect 222988 216668 297916 216696
rect 222988 216656 222994 216668
rect 297910 216656 297916 216668
rect 297968 216656 297974 216708
rect 247678 215296 247684 215348
rect 247736 215336 247742 215348
rect 297910 215336 297916 215348
rect 247736 215308 297916 215336
rect 247736 215296 247742 215308
rect 297910 215296 297916 215308
rect 297968 215296 297974 215348
rect 57238 214548 57244 214600
rect 57296 214588 57302 214600
rect 57698 214588 57704 214600
rect 57296 214560 57704 214588
rect 57296 214548 57302 214560
rect 57698 214548 57704 214560
rect 57756 214548 57762 214600
rect 246298 213936 246304 213988
rect 246356 213976 246362 213988
rect 297910 213976 297916 213988
rect 246356 213948 297916 213976
rect 246356 213936 246362 213948
rect 297910 213936 297916 213948
rect 297968 213936 297974 213988
rect 222286 212984 222292 213036
rect 222344 213024 222350 213036
rect 226058 213024 226064 213036
rect 222344 212996 226064 213024
rect 222344 212984 222350 212996
rect 226058 212984 226064 212996
rect 226116 212984 226122 213036
rect 242158 212508 242164 212560
rect 242216 212548 242222 212560
rect 297910 212548 297916 212560
rect 242216 212520 297916 212548
rect 242216 212508 242222 212520
rect 297910 212508 297916 212520
rect 297968 212508 297974 212560
rect 239398 211148 239404 211200
rect 239456 211188 239462 211200
rect 297910 211188 297916 211200
rect 239456 211160 297916 211188
rect 239456 211148 239462 211160
rect 297910 211148 297916 211160
rect 297968 211148 297974 211200
rect 238018 209788 238024 209840
rect 238076 209828 238082 209840
rect 297910 209828 297916 209840
rect 238076 209800 297916 209828
rect 238076 209788 238082 209800
rect 297910 209788 297916 209800
rect 297968 209788 297974 209840
rect 235258 208360 235264 208412
rect 235316 208400 235322 208412
rect 296806 208400 296812 208412
rect 235316 208372 296812 208400
rect 235316 208360 235322 208372
rect 296806 208360 296812 208372
rect 296864 208360 296870 208412
rect 287698 207000 287704 207052
rect 287756 207040 287762 207052
rect 297910 207040 297916 207052
rect 287756 207012 297916 207040
rect 287756 207000 287762 207012
rect 297910 207000 297916 207012
rect 297968 207000 297974 207052
rect 409138 206932 409144 206984
rect 409196 206972 409202 206984
rect 579798 206972 579804 206984
rect 409196 206944 579804 206972
rect 409196 206932 409202 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 284938 205640 284944 205692
rect 284996 205680 285002 205692
rect 296806 205680 296812 205692
rect 284996 205652 296812 205680
rect 284996 205640 285002 205652
rect 296806 205640 296812 205652
rect 296864 205640 296870 205692
rect 223206 205572 223212 205624
rect 223264 205612 223270 205624
rect 229738 205612 229744 205624
rect 223264 205584 229744 205612
rect 223264 205572 223270 205584
rect 229738 205572 229744 205584
rect 229796 205572 229802 205624
rect 282178 202852 282184 202904
rect 282236 202892 282242 202904
rect 297910 202892 297916 202904
rect 282236 202864 297916 202892
rect 282236 202852 282242 202864
rect 297910 202852 297916 202864
rect 297968 202852 297974 202904
rect 253198 201492 253204 201544
rect 253256 201532 253262 201544
rect 297910 201532 297916 201544
rect 253256 201504 297916 201532
rect 253256 201492 253262 201504
rect 297910 201492 297916 201504
rect 297968 201492 297974 201544
rect 51074 201424 51080 201476
rect 51132 201464 51138 201476
rect 57330 201464 57336 201476
rect 51132 201436 57336 201464
rect 51132 201424 51138 201436
rect 57330 201424 57336 201436
rect 57388 201424 57394 201476
rect 228358 200132 228364 200184
rect 228416 200172 228422 200184
rect 297910 200172 297916 200184
rect 228416 200144 297916 200172
rect 228416 200132 228422 200144
rect 297910 200132 297916 200144
rect 297968 200132 297974 200184
rect 225598 198704 225604 198756
rect 225656 198744 225662 198756
rect 297910 198744 297916 198756
rect 225656 198716 297916 198744
rect 225656 198704 225662 198716
rect 297910 198704 297916 198716
rect 297968 198704 297974 198756
rect 224310 197344 224316 197396
rect 224368 197384 224374 197396
rect 297910 197384 297916 197396
rect 224368 197356 297916 197384
rect 224368 197344 224374 197356
rect 297910 197344 297916 197356
rect 297968 197344 297974 197396
rect 50430 197276 50436 197328
rect 50488 197316 50494 197328
rect 57330 197316 57336 197328
rect 50488 197288 57336 197316
rect 50488 197276 50494 197288
rect 57330 197276 57336 197288
rect 57388 197276 57394 197328
rect 224218 195984 224224 196036
rect 224276 196024 224282 196036
rect 297910 196024 297916 196036
rect 224276 195996 297916 196024
rect 224276 195984 224282 195996
rect 297910 195984 297916 195996
rect 297968 195984 297974 196036
rect 223482 194556 223488 194608
rect 223540 194596 223546 194608
rect 233970 194596 233976 194608
rect 223540 194568 233976 194596
rect 223540 194556 223546 194568
rect 233970 194556 233976 194568
rect 234028 194556 234034 194608
rect 250438 194556 250444 194608
rect 250496 194596 250502 194608
rect 297910 194596 297916 194608
rect 250496 194568 297916 194596
rect 250496 194556 250502 194568
rect 297910 194556 297916 194568
rect 297968 194556 297974 194608
rect 243538 193196 243544 193248
rect 243596 193236 243602 193248
rect 297910 193236 297916 193248
rect 243596 193208 297916 193236
rect 243596 193196 243602 193208
rect 297910 193196 297916 193208
rect 297968 193196 297974 193248
rect 229738 193128 229744 193180
rect 229796 193168 229802 193180
rect 297726 193168 297732 193180
rect 229796 193140 297732 193168
rect 229796 193128 229802 193140
rect 297726 193128 297732 193140
rect 297784 193128 297790 193180
rect 516870 193128 516876 193180
rect 516928 193168 516934 193180
rect 580166 193168 580172 193180
rect 516928 193140 580172 193168
rect 516928 193128 516934 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 50982 192924 50988 192976
rect 51040 192964 51046 192976
rect 57330 192964 57336 192976
rect 51040 192936 57336 192964
rect 51040 192924 51046 192936
rect 57330 192924 57336 192936
rect 57388 192924 57394 192976
rect 223482 191836 223488 191888
rect 223540 191876 223546 191888
rect 232498 191876 232504 191888
rect 223540 191848 232504 191876
rect 223540 191836 223546 191848
rect 232498 191836 232504 191848
rect 232556 191836 232562 191888
rect 233878 190476 233884 190528
rect 233936 190516 233942 190528
rect 297910 190516 297916 190528
rect 233936 190488 297916 190516
rect 233936 190476 233942 190488
rect 297910 190476 297916 190488
rect 297968 190476 297974 190528
rect 222838 190408 222844 190460
rect 222896 190448 222902 190460
rect 297726 190448 297732 190460
rect 222896 190420 297732 190448
rect 222896 190408 222902 190420
rect 297726 190408 297732 190420
rect 297784 190408 297790 190460
rect 223482 189048 223488 189100
rect 223540 189088 223546 189100
rect 230382 189088 230388 189100
rect 223540 189060 230388 189088
rect 223540 189048 223546 189060
rect 230382 189048 230388 189060
rect 230440 189048 230446 189100
rect 50890 188980 50896 189032
rect 50948 189020 50954 189032
rect 57330 189020 57336 189032
rect 50948 188992 57336 189020
rect 50948 188980 50954 188992
rect 57330 188980 57336 188992
rect 57388 188980 57394 189032
rect 223022 188980 223028 189032
rect 223080 189020 223086 189032
rect 297910 189020 297916 189032
rect 223080 188992 297916 189020
rect 223080 188980 223086 188992
rect 297910 188980 297916 188992
rect 297968 188980 297974 189032
rect 223482 186328 223488 186380
rect 223540 186368 223546 186380
rect 295978 186368 295984 186380
rect 223540 186340 295984 186368
rect 223540 186328 223546 186340
rect 295978 186328 295984 186340
rect 296036 186328 296042 186380
rect 222930 186260 222936 186312
rect 222988 186300 222994 186312
rect 296806 186300 296812 186312
rect 222988 186272 296812 186300
rect 222988 186260 222994 186272
rect 296806 186260 296812 186272
rect 296864 186260 296870 186312
rect 51166 184832 51172 184884
rect 51224 184872 51230 184884
rect 56686 184872 56692 184884
rect 51224 184844 56692 184872
rect 51224 184832 51230 184844
rect 56686 184832 56692 184844
rect 56744 184832 56750 184884
rect 233970 184832 233976 184884
rect 234028 184872 234034 184884
rect 297910 184872 297916 184884
rect 234028 184844 297916 184872
rect 234028 184832 234034 184844
rect 297910 184832 297916 184844
rect 297968 184832 297974 184884
rect 222286 184152 222292 184204
rect 222344 184192 222350 184204
rect 225690 184192 225696 184204
rect 222344 184164 225696 184192
rect 222344 184152 222350 184164
rect 225690 184152 225696 184164
rect 225748 184152 225754 184204
rect 232498 183472 232504 183524
rect 232556 183512 232562 183524
rect 297910 183512 297916 183524
rect 232556 183484 297916 183512
rect 232556 183472 232562 183484
rect 297910 183472 297916 183484
rect 297968 183472 297974 183524
rect 230382 182112 230388 182164
rect 230440 182152 230446 182164
rect 297910 182152 297916 182164
rect 230440 182124 297916 182152
rect 230440 182112 230446 182124
rect 297910 182112 297916 182124
rect 297968 182112 297974 182164
rect 51258 180752 51264 180804
rect 51316 180792 51322 180804
rect 56686 180792 56692 180804
rect 51316 180764 56692 180792
rect 51316 180752 51322 180764
rect 56686 180752 56692 180764
rect 56744 180752 56750 180804
rect 225690 179324 225696 179376
rect 225748 179364 225754 179376
rect 297910 179364 297916 179376
rect 225748 179336 297916 179364
rect 225748 179324 225754 179336
rect 297910 179324 297916 179336
rect 297968 179324 297974 179376
rect 356882 179324 356888 179376
rect 356940 179364 356946 179376
rect 580166 179364 580172 179376
rect 356940 179336 580172 179364
rect 356940 179324 356946 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 223482 177964 223488 178016
rect 223540 178004 223546 178016
rect 297910 178004 297916 178016
rect 223540 177976 297916 178004
rect 223540 177964 223546 177976
rect 297910 177964 297916 177976
rect 297968 177964 297974 178016
rect 357618 177352 357624 177404
rect 357676 177392 357682 177404
rect 473446 177392 473452 177404
rect 357676 177364 473452 177392
rect 357676 177352 357682 177364
rect 473446 177352 473452 177364
rect 473504 177352 473510 177404
rect 382274 177284 382280 177336
rect 382332 177324 382338 177336
rect 521746 177324 521752 177336
rect 382332 177296 521752 177324
rect 382332 177284 382338 177296
rect 521746 177284 521752 177296
rect 521804 177284 521810 177336
rect 50338 176604 50344 176656
rect 50396 176644 50402 176656
rect 57330 176644 57336 176656
rect 50396 176616 57336 176644
rect 50396 176604 50402 176616
rect 57330 176604 57336 176616
rect 57388 176604 57394 176656
rect 222654 176604 222660 176656
rect 222712 176644 222718 176656
rect 297910 176644 297916 176656
rect 222712 176616 297916 176644
rect 222712 176604 222718 176616
rect 297910 176604 297916 176616
rect 297968 176604 297974 176656
rect 358538 175924 358544 175976
rect 358596 175964 358602 175976
rect 426434 175964 426440 175976
rect 358596 175936 426440 175964
rect 358596 175924 358602 175936
rect 426434 175924 426440 175936
rect 426492 175924 426498 175976
rect 222654 175176 222660 175228
rect 222712 175216 222718 175228
rect 297910 175216 297916 175228
rect 222712 175188 297916 175216
rect 222712 175176 222718 175188
rect 297910 175176 297916 175188
rect 297968 175176 297974 175228
rect 48866 173340 48872 173392
rect 48924 173380 48930 173392
rect 57238 173380 57244 173392
rect 48924 173352 57244 173380
rect 48924 173340 48930 173352
rect 57238 173340 57244 173352
rect 57296 173340 57302 173392
rect 222378 173136 222384 173188
rect 222436 173176 222442 173188
rect 297910 173176 297916 173188
rect 222436 173148 297916 173176
rect 222436 173136 222442 173148
rect 297910 173136 297916 173148
rect 297968 173136 297974 173188
rect 222470 171096 222476 171148
rect 222528 171136 222534 171148
rect 297910 171136 297916 171148
rect 222528 171108 297916 171136
rect 222528 171096 222534 171108
rect 297910 171096 297916 171108
rect 297968 171096 297974 171148
rect 222930 169736 222936 169788
rect 222988 169776 222994 169788
rect 296806 169776 296812 169788
rect 222988 169748 296812 169776
rect 222988 169736 222994 169748
rect 296806 169736 296812 169748
rect 296864 169736 296870 169788
rect 49510 169668 49516 169720
rect 49568 169708 49574 169720
rect 57330 169708 57336 169720
rect 49568 169680 57336 169708
rect 49568 169668 49574 169680
rect 57330 169668 57336 169680
rect 57388 169668 57394 169720
rect 223482 167016 223488 167068
rect 223540 167056 223546 167068
rect 297910 167056 297916 167068
rect 223540 167028 297916 167056
rect 223540 167016 223546 167028
rect 297910 167016 297916 167028
rect 297968 167016 297974 167068
rect 405090 166948 405096 167000
rect 405148 166988 405154 167000
rect 580166 166988 580172 167000
rect 405148 166960 580172 166988
rect 405148 166948 405154 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 223022 165588 223028 165640
rect 223080 165628 223086 165640
rect 297910 165628 297916 165640
rect 223080 165600 297916 165628
rect 223080 165588 223086 165600
rect 297910 165588 297916 165600
rect 297968 165588 297974 165640
rect 222930 164228 222936 164280
rect 222988 164268 222994 164280
rect 297910 164268 297916 164280
rect 222988 164240 297916 164268
rect 222988 164228 222994 164240
rect 297910 164228 297916 164240
rect 297968 164228 297974 164280
rect 223482 162868 223488 162920
rect 223540 162908 223546 162920
rect 297910 162908 297916 162920
rect 223540 162880 297916 162908
rect 223540 162868 223546 162880
rect 297910 162868 297916 162880
rect 297968 162868 297974 162920
rect 229094 161440 229100 161492
rect 229152 161480 229158 161492
rect 297910 161480 297916 161492
rect 229152 161452 297916 161480
rect 229152 161440 229158 161452
rect 297910 161440 297916 161452
rect 297968 161440 297974 161492
rect 54570 161372 54576 161424
rect 54628 161412 54634 161424
rect 57054 161412 57060 161424
rect 54628 161384 57060 161412
rect 54628 161372 54634 161384
rect 57054 161372 57060 161384
rect 57112 161372 57118 161424
rect 225782 158720 225788 158772
rect 225840 158760 225846 158772
rect 297910 158760 297916 158772
rect 225840 158732 297916 158760
rect 225840 158720 225846 158732
rect 297910 158720 297916 158732
rect 297968 158720 297974 158772
rect 232590 157360 232596 157412
rect 232648 157400 232654 157412
rect 297910 157400 297916 157412
rect 232648 157372 297916 157400
rect 232648 157360 232654 157372
rect 297910 157360 297916 157372
rect 297968 157360 297974 157412
rect 53098 157292 53104 157344
rect 53156 157332 53162 157344
rect 57054 157332 57060 157344
rect 53156 157304 57060 157332
rect 53156 157292 53162 157304
rect 57054 157292 57060 157304
rect 57112 157292 57118 157344
rect 222654 157292 222660 157344
rect 222712 157332 222718 157344
rect 229094 157332 229100 157344
rect 222712 157304 229100 157332
rect 222712 157292 222718 157304
rect 229094 157292 229100 157304
rect 229152 157292 229158 157344
rect 229830 155932 229836 155984
rect 229888 155972 229894 155984
rect 297910 155972 297916 155984
rect 229888 155944 297916 155972
rect 229888 155932 229894 155944
rect 297910 155932 297916 155944
rect 297968 155932 297974 155984
rect 222930 154572 222936 154624
rect 222988 154612 222994 154624
rect 297910 154612 297916 154624
rect 222988 154584 297916 154612
rect 222988 154572 222994 154584
rect 297910 154572 297916 154584
rect 297968 154572 297974 154624
rect 222838 153212 222844 153264
rect 222896 153252 222902 153264
rect 297910 153252 297916 153264
rect 222896 153224 297916 153252
rect 222896 153212 222902 153224
rect 297910 153212 297916 153224
rect 297968 153212 297974 153264
rect 54478 153144 54484 153196
rect 54536 153184 54542 153196
rect 57330 153184 57336 153196
rect 54536 153156 57336 153184
rect 54536 153144 54542 153156
rect 57330 153144 57336 153156
rect 57388 153144 57394 153196
rect 518618 153144 518624 153196
rect 518676 153184 518682 153196
rect 580166 153184 580172 153196
rect 518676 153156 580172 153184
rect 518676 153144 518682 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 231118 151784 231124 151836
rect 231176 151824 231182 151836
rect 296806 151824 296812 151836
rect 231176 151796 296812 151824
rect 231176 151784 231182 151796
rect 296806 151784 296812 151796
rect 296864 151784 296870 151836
rect 223206 151036 223212 151088
rect 223264 151076 223270 151088
rect 295978 151076 295984 151088
rect 223264 151048 295984 151076
rect 223264 151036 223270 151048
rect 295978 151036 295984 151048
rect 296036 151036 296042 151088
rect 2774 150288 2780 150340
rect 2832 150328 2838 150340
rect 4798 150328 4804 150340
rect 2832 150300 4804 150328
rect 2832 150288 2838 150300
rect 4798 150288 4804 150300
rect 4856 150288 4862 150340
rect 228450 149064 228456 149116
rect 228508 149104 228514 149116
rect 297910 149104 297916 149116
rect 228508 149076 297916 149104
rect 228508 149064 228514 149076
rect 297910 149064 297916 149076
rect 297968 149064 297974 149116
rect 50798 148996 50804 149048
rect 50856 149036 50862 149048
rect 57330 149036 57336 149048
rect 50856 149008 57336 149036
rect 50856 148996 50862 149008
rect 57330 148996 57336 149008
rect 57388 148996 57394 149048
rect 222562 147092 222568 147144
rect 222620 147132 222626 147144
rect 225782 147132 225788 147144
rect 222620 147104 225788 147132
rect 222620 147092 222626 147104
rect 225782 147092 225788 147104
rect 225840 147092 225846 147144
rect 225690 146276 225696 146328
rect 225748 146316 225754 146328
rect 297910 146316 297916 146328
rect 225748 146288 297916 146316
rect 225748 146276 225754 146288
rect 297910 146276 297916 146288
rect 297968 146276 297974 146328
rect 229738 144916 229744 144968
rect 229796 144956 229802 144968
rect 297910 144956 297916 144968
rect 229796 144928 297916 144956
rect 229796 144916 229802 144928
rect 297910 144916 297916 144928
rect 297968 144916 297974 144968
rect 223482 144848 223488 144900
rect 223540 144888 223546 144900
rect 232590 144888 232596 144900
rect 223540 144860 232596 144888
rect 223540 144848 223546 144860
rect 232590 144848 232596 144860
rect 232648 144848 232654 144900
rect 50706 144508 50712 144560
rect 50764 144548 50770 144560
rect 57330 144548 57336 144560
rect 50764 144520 57336 144548
rect 50764 144508 50770 144520
rect 57330 144508 57336 144520
rect 57388 144508 57394 144560
rect 232498 143556 232504 143608
rect 232556 143596 232562 143608
rect 297910 143596 297916 143608
rect 232556 143568 297916 143596
rect 232556 143556 232562 143568
rect 297910 143556 297916 143568
rect 297968 143556 297974 143608
rect 257338 142060 257344 142112
rect 257396 142100 257402 142112
rect 297910 142100 297916 142112
rect 257396 142072 297916 142100
rect 257396 142060 257402 142072
rect 297910 142060 297916 142072
rect 297968 142060 297974 142112
rect 223482 141448 223488 141500
rect 223540 141488 223546 141500
rect 229830 141488 229836 141500
rect 223540 141460 229836 141488
rect 223540 141448 223546 141460
rect 229830 141448 229836 141460
rect 229888 141448 229894 141500
rect 51350 140700 51356 140752
rect 51408 140740 51414 140752
rect 57422 140740 57428 140752
rect 51408 140712 57428 140740
rect 51408 140700 51414 140712
rect 57422 140700 57428 140712
rect 57480 140700 57486 140752
rect 257430 140700 257436 140752
rect 257488 140740 257494 140752
rect 297910 140740 297916 140752
rect 257488 140712 297916 140740
rect 257488 140700 257494 140712
rect 297910 140700 297916 140712
rect 297968 140700 297974 140752
rect 269850 139340 269856 139392
rect 269908 139380 269914 139392
rect 297910 139380 297916 139392
rect 269908 139352 297916 139380
rect 269908 139340 269914 139352
rect 297910 139340 297916 139352
rect 297968 139340 297974 139392
rect 354030 139340 354036 139392
rect 354088 139380 354094 139392
rect 580166 139380 580172 139392
rect 354088 139352 580172 139380
rect 354088 139340 354094 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 222654 137912 222660 137964
rect 222712 137952 222718 137964
rect 231118 137952 231124 137964
rect 222712 137924 231124 137952
rect 222712 137912 222718 137924
rect 231118 137912 231124 137924
rect 231176 137912 231182 137964
rect 275370 137912 275376 137964
rect 275428 137952 275434 137964
rect 297910 137952 297916 137964
rect 275428 137924 297916 137952
rect 275428 137912 275434 137924
rect 297910 137912 297916 137924
rect 297968 137912 297974 137964
rect 273990 136552 273996 136604
rect 274048 136592 274054 136604
rect 297910 136592 297916 136604
rect 274048 136564 297916 136592
rect 274048 136552 274054 136564
rect 297910 136552 297916 136564
rect 297968 136552 297974 136604
rect 274082 135192 274088 135244
rect 274140 135232 274146 135244
rect 297910 135232 297916 135244
rect 274140 135204 297916 135232
rect 274140 135192 274146 135204
rect 297910 135192 297916 135204
rect 297968 135192 297974 135244
rect 222838 133152 222844 133204
rect 222896 133192 222902 133204
rect 296070 133192 296076 133204
rect 222896 133164 296076 133192
rect 222896 133152 222902 133164
rect 296070 133152 296076 133164
rect 296128 133152 296134 133204
rect 258718 132404 258724 132456
rect 258776 132444 258782 132456
rect 296806 132444 296812 132456
rect 258776 132416 296812 132444
rect 258776 132404 258782 132416
rect 296806 132404 296812 132416
rect 296864 132404 296870 132456
rect 271230 131044 271236 131096
rect 271288 131084 271294 131096
rect 297910 131084 297916 131096
rect 271288 131056 297916 131084
rect 271288 131044 271294 131056
rect 297910 131044 297916 131056
rect 297968 131044 297974 131096
rect 223022 130024 223028 130076
rect 223080 130064 223086 130076
rect 228450 130064 228456 130076
rect 223080 130036 228456 130064
rect 223080 130024 223086 130036
rect 228450 130024 228456 130036
rect 228508 130024 228514 130076
rect 269942 129684 269948 129736
rect 270000 129724 270006 129736
rect 296806 129724 296812 129736
rect 270000 129696 296812 129724
rect 270000 129684 270006 129696
rect 296806 129684 296812 129696
rect 296864 129684 296870 129736
rect 222286 128256 222292 128308
rect 222344 128296 222350 128308
rect 225690 128296 225696 128308
rect 222344 128268 225696 128296
rect 222344 128256 222350 128268
rect 225690 128256 225696 128268
rect 225748 128256 225754 128308
rect 262858 128256 262864 128308
rect 262916 128296 262922 128308
rect 297910 128296 297916 128308
rect 262916 128268 297916 128296
rect 262916 128256 262922 128268
rect 297910 128256 297916 128268
rect 297968 128256 297974 128308
rect 261570 126896 261576 126948
rect 261628 126936 261634 126948
rect 297910 126936 297916 126948
rect 261628 126908 297916 126936
rect 261628 126896 261634 126908
rect 297910 126896 297916 126908
rect 297968 126896 297974 126948
rect 372890 126896 372896 126948
rect 372948 126936 372954 126948
rect 580166 126936 580172 126948
rect 372948 126908 580172 126936
rect 372948 126896 372954 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 279510 125536 279516 125588
rect 279568 125576 279574 125588
rect 297910 125576 297916 125588
rect 279568 125548 297916 125576
rect 279568 125536 279574 125548
rect 297910 125536 297916 125548
rect 297968 125536 297974 125588
rect 268470 124108 268476 124160
rect 268528 124148 268534 124160
rect 297910 124148 297916 124160
rect 268528 124120 297916 124148
rect 268528 124108 268534 124120
rect 297910 124108 297916 124120
rect 297968 124108 297974 124160
rect 265710 122748 265716 122800
rect 265768 122788 265774 122800
rect 297910 122788 297916 122800
rect 265768 122760 297916 122788
rect 265768 122748 265774 122760
rect 297910 122748 297916 122760
rect 297968 122748 297974 122800
rect 264330 121388 264336 121440
rect 264388 121428 264394 121440
rect 297910 121428 297916 121440
rect 264388 121400 297916 121428
rect 264388 121388 264394 121400
rect 297910 121388 297916 121400
rect 297968 121388 297974 121440
rect 223482 120640 223488 120692
rect 223540 120680 223546 120692
rect 229738 120680 229744 120692
rect 223540 120652 229744 120680
rect 223540 120640 223546 120652
rect 229738 120640 229744 120652
rect 229796 120640 229802 120692
rect 271322 120028 271328 120080
rect 271380 120068 271386 120080
rect 297910 120068 297916 120080
rect 271380 120040 297916 120068
rect 271380 120028 271386 120040
rect 297910 120028 297916 120040
rect 297968 120028 297974 120080
rect 223482 118600 223488 118652
rect 223540 118640 223546 118652
rect 232498 118640 232504 118652
rect 223540 118612 232504 118640
rect 223540 118600 223546 118612
rect 232498 118600 232504 118612
rect 232556 118600 232562 118652
rect 278222 118600 278228 118652
rect 278280 118640 278286 118652
rect 297910 118640 297916 118652
rect 278280 118612 297916 118640
rect 278280 118600 278286 118612
rect 297910 118600 297916 118612
rect 297968 118600 297974 118652
rect 289078 117240 289084 117292
rect 289136 117280 289142 117292
rect 297910 117280 297916 117292
rect 289136 117252 297916 117280
rect 289136 117240 289142 117252
rect 297910 117240 297916 117252
rect 297968 117240 297974 117292
rect 342346 117240 342352 117292
rect 342404 117280 342410 117292
rect 363598 117280 363604 117292
rect 342404 117252 363604 117280
rect 342404 117240 342410 117252
rect 363598 117240 363604 117252
rect 363656 117240 363662 117292
rect 223482 115880 223488 115932
rect 223540 115920 223546 115932
rect 295978 115920 295984 115932
rect 223540 115892 295984 115920
rect 223540 115880 223546 115892
rect 295978 115880 295984 115892
rect 296036 115880 296042 115932
rect 275462 114452 275468 114504
rect 275520 114492 275526 114504
rect 296806 114492 296812 114504
rect 275520 114464 296812 114492
rect 275520 114452 275526 114464
rect 296806 114452 296812 114464
rect 296864 114452 296870 114504
rect 257522 113092 257528 113144
rect 257580 113132 257586 113144
rect 297910 113132 297916 113144
rect 257580 113104 297916 113132
rect 257580 113092 257586 113104
rect 297910 113092 297916 113104
rect 297968 113092 297974 113144
rect 530578 113092 530584 113144
rect 530636 113132 530642 113144
rect 579798 113132 579804 113144
rect 530636 113104 579804 113132
rect 530636 113092 530642 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 222194 112956 222200 113008
rect 222252 112996 222258 113008
rect 224402 112996 224408 113008
rect 222252 112968 224408 112996
rect 222252 112956 222258 112968
rect 224402 112956 224408 112968
rect 224460 112956 224466 113008
rect 223482 110372 223488 110424
rect 223540 110412 223546 110424
rect 247678 110412 247684 110424
rect 223540 110384 247684 110412
rect 223540 110372 223546 110384
rect 247678 110372 247684 110384
rect 247736 110372 247742 110424
rect 357710 109692 357716 109744
rect 357768 109732 357774 109744
rect 580258 109732 580264 109744
rect 357768 109704 580264 109732
rect 357768 109692 357774 109704
rect 580258 109692 580264 109704
rect 580316 109692 580322 109744
rect 342346 108944 342352 108996
rect 342404 108984 342410 108996
rect 440878 108984 440884 108996
rect 342404 108956 440884 108984
rect 342404 108944 342410 108956
rect 440878 108944 440884 108956
rect 440936 108944 440942 108996
rect 222654 107584 222660 107636
rect 222712 107624 222718 107636
rect 246298 107624 246304 107636
rect 222712 107596 246304 107624
rect 222712 107584 222718 107596
rect 246298 107584 246304 107596
rect 246356 107584 246362 107636
rect 342346 106224 342352 106276
rect 342404 106264 342410 106276
rect 518250 106264 518256 106276
rect 342404 106236 518256 106264
rect 342404 106224 342410 106236
rect 518250 106224 518256 106236
rect 518308 106224 518314 106276
rect 222838 104796 222844 104848
rect 222896 104836 222902 104848
rect 242158 104836 242164 104848
rect 222896 104808 242164 104836
rect 222896 104796 222902 104808
rect 242158 104796 242164 104808
rect 242216 104796 242222 104848
rect 223482 102076 223488 102128
rect 223540 102116 223546 102128
rect 239398 102116 239404 102128
rect 223540 102088 239404 102116
rect 223540 102076 223546 102088
rect 239398 102076 239404 102088
rect 239456 102076 239462 102128
rect 223022 99288 223028 99340
rect 223080 99328 223086 99340
rect 238018 99328 238024 99340
rect 223080 99300 238024 99328
rect 223080 99288 223086 99300
rect 238018 99288 238024 99300
rect 238076 99288 238082 99340
rect 223114 96568 223120 96620
rect 223172 96608 223178 96620
rect 235258 96608 235264 96620
rect 223172 96580 235264 96608
rect 223172 96568 223178 96580
rect 235258 96568 235264 96580
rect 235316 96568 235322 96620
rect 223482 93780 223488 93832
rect 223540 93820 223546 93832
rect 287698 93820 287704 93832
rect 223540 93792 287704 93820
rect 223540 93780 223546 93792
rect 287698 93780 287704 93792
rect 287756 93780 287762 93832
rect 223482 91740 223488 91792
rect 223540 91780 223546 91792
rect 284938 91780 284944 91792
rect 223540 91752 284944 91780
rect 223540 91740 223546 91752
rect 284938 91740 284944 91752
rect 284996 91740 285002 91792
rect 266998 90312 267004 90364
rect 267056 90352 267062 90364
rect 297358 90352 297364 90364
rect 267056 90324 297364 90352
rect 267056 90312 267062 90324
rect 297358 90312 297364 90324
rect 297416 90312 297422 90364
rect 264238 88952 264244 89004
rect 264296 88992 264302 89004
rect 296806 88992 296812 89004
rect 264296 88964 296812 88992
rect 264296 88952 264302 88964
rect 296806 88952 296812 88964
rect 296864 88952 296870 89004
rect 357802 88952 357808 89004
rect 357860 88992 357866 89004
rect 415394 88992 415400 89004
rect 357860 88964 415400 88992
rect 357860 88952 357866 88964
rect 415394 88952 415400 88964
rect 415452 88952 415458 89004
rect 223206 88272 223212 88324
rect 223264 88312 223270 88324
rect 282178 88312 282184 88324
rect 223264 88284 282184 88312
rect 223264 88272 223270 88284
rect 282178 88272 282184 88284
rect 282236 88272 282242 88324
rect 291838 88272 291844 88324
rect 291896 88312 291902 88324
rect 298002 88312 298008 88324
rect 291896 88284 298008 88312
rect 291896 88272 291902 88284
rect 298002 88272 298008 88284
rect 298060 88272 298066 88324
rect 260190 86912 260196 86964
rect 260248 86952 260254 86964
rect 297174 86952 297180 86964
rect 260248 86924 297180 86952
rect 260248 86912 260254 86924
rect 297174 86912 297180 86924
rect 297232 86912 297238 86964
rect 223206 85484 223212 85536
rect 223264 85524 223270 85536
rect 253198 85524 253204 85536
rect 223264 85496 253204 85524
rect 223264 85484 223270 85496
rect 253198 85484 253204 85496
rect 253256 85484 253262 85536
rect 3418 85008 3424 85060
rect 3476 85048 3482 85060
rect 8938 85048 8944 85060
rect 3476 85020 8944 85048
rect 3476 85008 3482 85020
rect 8938 85008 8944 85020
rect 8996 85008 9002 85060
rect 273898 84124 273904 84176
rect 273956 84164 273962 84176
rect 297910 84164 297916 84176
rect 273956 84136 297916 84164
rect 273956 84124 273962 84136
rect 297910 84124 297916 84136
rect 297968 84124 297974 84176
rect 271138 82764 271144 82816
rect 271196 82804 271202 82816
rect 297910 82804 297916 82816
rect 271196 82776 297916 82804
rect 271196 82764 271202 82776
rect 297910 82764 297916 82776
rect 297968 82764 297974 82816
rect 223482 81336 223488 81388
rect 223540 81376 223546 81388
rect 228358 81376 228364 81388
rect 223540 81348 228364 81376
rect 223540 81336 223546 81348
rect 228358 81336 228364 81348
rect 228416 81336 228422 81388
rect 269758 79976 269764 80028
rect 269816 80016 269822 80028
rect 298002 80016 298008 80028
rect 269816 79988 298008 80016
rect 269816 79976 269822 79988
rect 298002 79976 298008 79988
rect 298060 79976 298066 80028
rect 275278 78616 275284 78668
rect 275336 78656 275342 78668
rect 297542 78656 297548 78668
rect 275336 78628 297548 78656
rect 275336 78616 275342 78628
rect 297542 78616 297548 78628
rect 297600 78616 297606 78668
rect 222470 78548 222476 78600
rect 222528 78588 222534 78600
rect 225598 78588 225604 78600
rect 222528 78560 225604 78588
rect 222528 78548 222534 78560
rect 225598 78548 225604 78560
rect 225656 78548 225662 78600
rect 260098 77188 260104 77240
rect 260156 77228 260162 77240
rect 297174 77228 297180 77240
rect 260156 77200 297180 77228
rect 260156 77188 260162 77200
rect 297174 77188 297180 77200
rect 297232 77188 297238 77240
rect 255958 75828 255964 75880
rect 256016 75868 256022 75880
rect 298002 75868 298008 75880
rect 256016 75840 298008 75868
rect 256016 75828 256022 75840
rect 298002 75828 298008 75840
rect 298060 75828 298066 75880
rect 222194 75692 222200 75744
rect 222252 75732 222258 75744
rect 224310 75732 224316 75744
rect 222252 75704 224316 75732
rect 222252 75692 222258 75704
rect 224310 75692 224316 75704
rect 224368 75692 224374 75744
rect 278038 74468 278044 74520
rect 278096 74508 278102 74520
rect 298002 74508 298008 74520
rect 278096 74480 298008 74508
rect 278096 74468 278102 74480
rect 298002 74468 298008 74480
rect 298060 74468 298066 74520
rect 256050 73108 256056 73160
rect 256108 73148 256114 73160
rect 296806 73148 296812 73160
rect 256108 73120 296812 73148
rect 256108 73108 256114 73120
rect 296806 73108 296812 73120
rect 296864 73108 296870 73160
rect 542998 73108 543004 73160
rect 543056 73148 543062 73160
rect 580166 73148 580172 73160
rect 543056 73120 580172 73148
rect 543056 73108 543062 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 222194 73040 222200 73092
rect 222252 73080 222258 73092
rect 224218 73080 224224 73092
rect 222252 73052 224224 73080
rect 222252 73040 222258 73052
rect 224218 73040 224224 73052
rect 224276 73040 224282 73092
rect 279418 71680 279424 71732
rect 279476 71720 279482 71732
rect 297726 71720 297732 71732
rect 279476 71692 297732 71720
rect 279476 71680 279482 71692
rect 297726 71680 297732 71692
rect 297784 71680 297790 71732
rect 223482 70320 223488 70372
rect 223540 70360 223546 70372
rect 250438 70360 250444 70372
rect 223540 70332 250444 70360
rect 223540 70320 223546 70332
rect 250438 70320 250444 70332
rect 250496 70320 250502 70372
rect 265618 70320 265624 70372
rect 265676 70360 265682 70372
rect 298002 70360 298008 70372
rect 265676 70332 298008 70360
rect 265676 70320 265682 70332
rect 298002 70320 298008 70332
rect 298060 70320 298066 70372
rect 342990 69028 342996 69080
rect 343048 69068 343054 69080
rect 489914 69068 489920 69080
rect 343048 69040 489920 69068
rect 343048 69028 343054 69040
rect 489914 69028 489920 69040
rect 489972 69028 489978 69080
rect 268378 68960 268384 69012
rect 268436 69000 268442 69012
rect 297174 69000 297180 69012
rect 268436 68972 297180 69000
rect 268436 68960 268442 68972
rect 297174 68960 297180 68972
rect 297232 68960 297238 69012
rect 223482 67532 223488 67584
rect 223540 67572 223546 67584
rect 243538 67572 243544 67584
rect 223540 67544 243544 67572
rect 223540 67532 223546 67544
rect 243538 67532 243544 67544
rect 243596 67532 243602 67584
rect 261478 67532 261484 67584
rect 261536 67572 261542 67584
rect 297542 67572 297548 67584
rect 261536 67544 297548 67572
rect 261536 67532 261542 67544
rect 297542 67532 297548 67544
rect 297600 67532 297606 67584
rect 342990 66240 342996 66292
rect 343048 66280 343054 66292
rect 418890 66280 418896 66292
rect 343048 66252 418896 66280
rect 343048 66240 343054 66252
rect 418890 66240 418896 66252
rect 418948 66240 418954 66292
rect 222838 64812 222844 64864
rect 222896 64852 222902 64864
rect 233878 64852 233884 64864
rect 222896 64824 233884 64852
rect 222896 64812 222902 64824
rect 233878 64812 233884 64824
rect 233936 64812 233942 64864
rect 278130 64812 278136 64864
rect 278188 64852 278194 64864
rect 297910 64852 297916 64864
rect 278188 64824 297916 64852
rect 278188 64812 278194 64824
rect 297910 64812 297916 64824
rect 297968 64812 297974 64864
rect 342990 63520 342996 63572
rect 343048 63560 343054 63572
rect 483014 63560 483020 63572
rect 343048 63532 483020 63560
rect 343048 63520 343054 63532
rect 483014 63520 483020 63532
rect 483072 63520 483078 63572
rect 342438 62840 342444 62892
rect 342496 62880 342502 62892
rect 342990 62880 342996 62892
rect 342496 62852 342996 62880
rect 342496 62840 342502 62852
rect 342990 62840 342996 62852
rect 343048 62840 343054 62892
rect 342346 62092 342352 62144
rect 342404 62132 342410 62144
rect 480254 62132 480260 62144
rect 342404 62104 480260 62132
rect 342404 62092 342410 62104
rect 480254 62092 480260 62104
rect 480312 62092 480318 62144
rect 264422 62024 264428 62076
rect 264480 62064 264486 62076
rect 298002 62064 298008 62076
rect 264480 62036 298008 62064
rect 264480 62024 264486 62036
rect 298002 62024 298008 62036
rect 298060 62024 298066 62076
rect 215294 61480 215300 61532
rect 215352 61520 215358 61532
rect 342622 61520 342628 61532
rect 215352 61492 342628 61520
rect 215352 61480 215358 61492
rect 342622 61480 342628 61492
rect 342680 61480 342686 61532
rect 158714 61412 158720 61464
rect 158772 61452 158778 61464
rect 342806 61452 342812 61464
rect 158772 61424 342812 61452
rect 158772 61412 158778 61424
rect 342806 61412 342812 61424
rect 342864 61412 342870 61464
rect 154574 61344 154580 61396
rect 154632 61384 154638 61396
rect 342898 61384 342904 61396
rect 154632 61356 342904 61384
rect 154632 61344 154638 61356
rect 342898 61344 342904 61356
rect 342956 61344 342962 61396
rect 353938 60664 353944 60716
rect 353996 60704 354002 60716
rect 580166 60704 580172 60716
rect 353996 60676 580172 60704
rect 353996 60664 354002 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 296622 60324 296628 60376
rect 296680 60364 296686 60376
rect 303614 60364 303620 60376
rect 296680 60336 303620 60364
rect 296680 60324 296686 60336
rect 303614 60324 303620 60336
rect 303672 60324 303678 60376
rect 295242 60256 295248 60308
rect 295300 60296 295306 60308
rect 310514 60296 310520 60308
rect 295300 60268 310520 60296
rect 295300 60256 295306 60268
rect 310514 60256 310520 60268
rect 310572 60256 310578 60308
rect 314654 60256 314660 60308
rect 314712 60296 314718 60308
rect 355594 60296 355600 60308
rect 314712 60268 355600 60296
rect 314712 60256 314718 60268
rect 355594 60256 355600 60268
rect 355652 60256 355658 60308
rect 211154 60188 211160 60240
rect 211212 60228 211218 60240
rect 342714 60228 342720 60240
rect 211212 60200 342720 60228
rect 211212 60188 211218 60200
rect 342714 60188 342720 60200
rect 342772 60188 342778 60240
rect 197354 60120 197360 60172
rect 197412 60160 197418 60172
rect 341334 60160 341340 60172
rect 197412 60132 341340 60160
rect 197412 60120 197418 60132
rect 341334 60120 341340 60132
rect 341392 60120 341398 60172
rect 168374 60052 168380 60104
rect 168432 60092 168438 60104
rect 341702 60092 341708 60104
rect 168432 60064 341708 60092
rect 168432 60052 168438 60064
rect 341702 60052 341708 60064
rect 341760 60052 341766 60104
rect 133874 59984 133880 60036
rect 133932 60024 133938 60036
rect 340506 60024 340512 60036
rect 133932 59996 340512 60024
rect 133932 59984 133938 59996
rect 340506 59984 340512 59996
rect 340564 59984 340570 60036
rect 247034 58828 247040 58880
rect 247092 58868 247098 58880
rect 340138 58868 340144 58880
rect 247092 58840 340144 58868
rect 247092 58828 247098 58840
rect 340138 58828 340144 58840
rect 340196 58828 340202 58880
rect 172514 58760 172520 58812
rect 172572 58800 172578 58812
rect 341610 58800 341616 58812
rect 172572 58772 341616 58800
rect 172572 58760 172578 58772
rect 341610 58760 341616 58772
rect 341668 58760 341674 58812
rect 151814 58692 151820 58744
rect 151872 58732 151878 58744
rect 343174 58732 343180 58744
rect 151872 58704 343180 58732
rect 151872 58692 151878 58704
rect 343174 58692 343180 58704
rect 343232 58692 343238 58744
rect 140774 58624 140780 58676
rect 140832 58664 140838 58676
rect 342438 58664 342444 58676
rect 140832 58636 342444 58664
rect 140832 58624 140838 58636
rect 342438 58624 342444 58636
rect 342496 58624 342502 58676
rect 233234 57332 233240 57384
rect 233292 57372 233298 57384
rect 342990 57372 342996 57384
rect 233292 57344 342996 57372
rect 233292 57332 233298 57344
rect 342990 57332 342996 57344
rect 343048 57332 343054 57384
rect 179414 57264 179420 57316
rect 179472 57304 179478 57316
rect 341426 57304 341432 57316
rect 179472 57276 341432 57304
rect 179472 57264 179478 57276
rect 341426 57264 341432 57276
rect 341484 57264 341490 57316
rect 176654 57196 176660 57248
rect 176712 57236 176718 57248
rect 341518 57236 341524 57248
rect 176712 57208 341524 57236
rect 176712 57196 176718 57208
rect 341518 57196 341524 57208
rect 341576 57196 341582 57248
rect 235994 55904 236000 55956
rect 236052 55944 236058 55956
rect 340230 55944 340236 55956
rect 236052 55916 340236 55944
rect 236052 55904 236058 55916
rect 340230 55904 340236 55916
rect 340288 55904 340294 55956
rect 190454 55836 190460 55888
rect 190512 55876 190518 55888
rect 340414 55876 340420 55888
rect 190512 55848 340420 55876
rect 190512 55836 190518 55848
rect 340414 55836 340420 55848
rect 340472 55836 340478 55888
rect 218054 54476 218060 54528
rect 218112 54516 218118 54528
rect 342530 54516 342536 54528
rect 218112 54488 342536 54516
rect 218112 54476 218118 54488
rect 342530 54476 342536 54488
rect 342588 54476 342594 54528
rect 226334 53048 226340 53100
rect 226392 53088 226398 53100
rect 341150 53088 341156 53100
rect 226392 53060 341156 53088
rect 226392 53048 226398 53060
rect 341150 53048 341156 53060
rect 341208 53048 341214 53100
rect 251174 51688 251180 51740
rect 251232 51728 251238 51740
rect 341058 51728 341064 51740
rect 251232 51700 341064 51728
rect 251232 51688 251238 51700
rect 341058 51688 341064 51700
rect 341116 51688 341122 51740
rect 201494 47540 201500 47592
rect 201552 47580 201558 47592
rect 498838 47580 498844 47592
rect 201552 47552 498844 47580
rect 201552 47540 201558 47552
rect 498838 47540 498844 47552
rect 498896 47540 498902 47592
rect 359550 46860 359556 46912
rect 359608 46900 359614 46912
rect 580166 46900 580172 46912
rect 359608 46872 580172 46900
rect 359608 46860 359614 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 242894 46180 242900 46232
rect 242952 46220 242958 46232
rect 343082 46220 343088 46232
rect 242952 46192 343088 46220
rect 242952 46180 242958 46192
rect 343082 46180 343088 46192
rect 343140 46180 343146 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 355502 45540 355508 45552
rect 3476 45512 355508 45540
rect 3476 45500 3482 45512
rect 355502 45500 355508 45512
rect 355560 45500 355566 45552
rect 204254 44820 204260 44872
rect 204312 44860 204318 44872
rect 340322 44860 340328 44872
rect 204312 44832 340328 44860
rect 204312 44820 204318 44832
rect 340322 44820 340328 44832
rect 340380 44820 340386 44872
rect 222194 42168 222200 42220
rect 222252 42208 222258 42220
rect 340046 42208 340052 42220
rect 222252 42180 340052 42208
rect 222252 42168 222258 42180
rect 340046 42168 340052 42180
rect 340104 42168 340110 42220
rect 193214 42100 193220 42152
rect 193272 42140 193278 42152
rect 341242 42140 341248 42152
rect 193272 42112 341248 42140
rect 193272 42100 193278 42112
rect 341242 42100 341248 42112
rect 341300 42100 341306 42152
rect 99374 42032 99380 42084
rect 99432 42072 99438 42084
rect 520550 42072 520556 42084
rect 99432 42044 520556 42072
rect 99432 42032 99438 42044
rect 520550 42032 520556 42044
rect 520608 42032 520614 42084
rect 120074 40672 120080 40724
rect 120132 40712 120138 40724
rect 509694 40712 509700 40724
rect 120132 40684 509700 40712
rect 120132 40672 120138 40684
rect 509694 40672 509700 40684
rect 509752 40672 509758 40724
rect 85574 35164 85580 35216
rect 85632 35204 85638 35216
rect 486418 35204 486424 35216
rect 85632 35176 486424 35204
rect 85632 35164 85638 35176
rect 486418 35164 486424 35176
rect 486476 35164 486482 35216
rect 510890 33056 510896 33108
rect 510948 33096 510954 33108
rect 580166 33096 580172 33108
rect 510948 33068 580172 33096
rect 510948 33056 510954 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 77294 32376 77300 32428
rect 77352 32416 77358 32428
rect 436738 32416 436744 32428
rect 77352 32388 436744 32416
rect 77352 32376 77358 32388
rect 436738 32376 436744 32388
rect 436796 32376 436802 32428
rect 74534 31016 74540 31068
rect 74592 31056 74598 31068
rect 493318 31056 493324 31068
rect 74592 31028 493324 31056
rect 74592 31016 74598 31028
rect 493318 31016 493324 31028
rect 493376 31016 493382 31068
rect 349154 28296 349160 28348
rect 349212 28336 349218 28348
rect 476850 28336 476856 28348
rect 349212 28308 476856 28336
rect 349212 28296 349218 28308
rect 476850 28296 476856 28308
rect 476908 28296 476914 28348
rect 113174 28228 113180 28280
rect 113232 28268 113238 28280
rect 454678 28268 454684 28280
rect 113232 28240 454684 28268
rect 113232 28228 113238 28240
rect 454678 28228 454684 28240
rect 454736 28228 454742 28280
rect 63494 26868 63500 26920
rect 63552 26908 63558 26920
rect 472618 26908 472624 26920
rect 63552 26880 472624 26908
rect 63552 26868 63558 26880
rect 472618 26868 472624 26880
rect 472676 26868 472682 26920
rect 60734 25508 60740 25560
rect 60792 25548 60798 25560
rect 475470 25548 475476 25560
rect 60792 25520 475476 25548
rect 60792 25508 60798 25520
rect 475470 25508 475476 25520
rect 475528 25508 475534 25560
rect 391934 24080 391940 24132
rect 391992 24120 391998 24132
rect 468478 24120 468484 24132
rect 391992 24092 468484 24120
rect 391992 24080 391998 24092
rect 468478 24080 468484 24092
rect 468536 24080 468542 24132
rect 346394 22720 346400 22772
rect 346452 22760 346458 22772
rect 413278 22760 413284 22772
rect 346452 22732 413284 22760
rect 346452 22720 346458 22732
rect 413278 22720 413284 22732
rect 413336 22720 413342 22772
rect 392210 21428 392216 21480
rect 392268 21468 392274 21480
rect 412634 21468 412640 21480
rect 392268 21440 412640 21468
rect 392268 21428 392274 21440
rect 412634 21428 412640 21440
rect 412692 21428 412698 21480
rect 2774 21360 2780 21412
rect 2832 21400 2838 21412
rect 422938 21400 422944 21412
rect 2832 21372 422944 21400
rect 2832 21360 2838 21372
rect 422938 21360 422944 21372
rect 422996 21360 423002 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 450538 20652 450544 20664
rect 3476 20624 450544 20652
rect 3476 20612 3482 20624
rect 450538 20612 450544 20624
rect 450596 20612 450602 20664
rect 356790 20544 356796 20596
rect 356848 20584 356854 20596
rect 580166 20584 580172 20596
rect 356848 20556 580172 20584
rect 356848 20544 356854 20556
rect 580166 20544 580172 20556
rect 580224 20544 580230 20596
rect 1394 18572 1400 18624
rect 1452 18612 1458 18624
rect 476758 18612 476764 18624
rect 1452 18584 476764 18612
rect 1452 18572 1458 18584
rect 476758 18572 476764 18584
rect 476816 18572 476822 18624
rect 378134 17212 378140 17264
rect 378192 17252 378198 17264
rect 462958 17252 462964 17264
rect 378192 17224 462964 17252
rect 378192 17212 378198 17224
rect 462958 17212 462964 17224
rect 463016 17212 463022 17264
rect 390922 15920 390928 15972
rect 390980 15960 390986 15972
rect 440234 15960 440240 15972
rect 390980 15932 440240 15960
rect 390980 15920 390986 15932
rect 440234 15920 440240 15932
rect 440292 15920 440298 15972
rect 95786 15852 95792 15904
rect 95844 15892 95850 15904
rect 400858 15892 400864 15904
rect 95844 15864 400864 15892
rect 95844 15852 95850 15864
rect 400858 15852 400864 15864
rect 400916 15852 400922 15904
rect 367738 14492 367744 14544
rect 367796 14532 367802 14544
rect 418798 14532 418804 14544
rect 367796 14504 418804 14532
rect 367796 14492 367802 14504
rect 418798 14492 418804 14504
rect 418856 14492 418862 14544
rect 102134 14424 102140 14476
rect 102192 14464 102198 14476
rect 519906 14464 519912 14476
rect 102192 14436 519912 14464
rect 102192 14424 102198 14436
rect 519906 14424 519912 14436
rect 519964 14424 519970 14476
rect 258258 13064 258264 13116
rect 258316 13104 258322 13116
rect 494698 13104 494704 13116
rect 258316 13076 494704 13104
rect 258316 13064 258322 13076
rect 494698 13064 494704 13076
rect 494756 13064 494762 13116
rect 240134 10276 240140 10328
rect 240192 10316 240198 10328
rect 340874 10316 340880 10328
rect 240192 10288 340880 10316
rect 240192 10276 240198 10288
rect 340874 10276 340880 10288
rect 340932 10276 340938 10328
rect 427722 9052 427728 9104
rect 427780 9092 427786 9104
rect 494698 9092 494704 9104
rect 427780 9064 494704 9092
rect 427780 9052 427786 9064
rect 494698 9052 494704 9064
rect 494756 9052 494762 9104
rect 110506 8984 110512 9036
rect 110564 9024 110570 9036
rect 521102 9024 521108 9036
rect 110564 8996 521108 9024
rect 110564 8984 110570 8996
rect 521102 8984 521108 8996
rect 521160 8984 521166 9036
rect 82078 8916 82084 8968
rect 82136 8956 82142 8968
rect 521010 8956 521016 8968
rect 82136 8928 521016 8956
rect 82136 8916 82142 8928
rect 521010 8916 521016 8928
rect 521068 8916 521074 8968
rect 396166 8236 396172 8288
rect 396224 8276 396230 8288
rect 402514 8276 402520 8288
rect 396224 8248 402520 8276
rect 396224 8236 396230 8248
rect 402514 8236 402520 8248
rect 402572 8236 402578 8288
rect 229830 7624 229836 7676
rect 229888 7664 229894 7676
rect 342254 7664 342260 7676
rect 229888 7636 342260 7664
rect 229888 7624 229894 7636
rect 342254 7624 342260 7636
rect 342312 7624 342318 7676
rect 418890 7624 418896 7676
rect 418948 7664 418954 7676
rect 487614 7664 487620 7676
rect 418948 7636 487620 7664
rect 418948 7624 418954 7636
rect 487614 7624 487620 7636
rect 487672 7624 487678 7676
rect 39574 7556 39580 7608
rect 39632 7596 39638 7608
rect 522574 7596 522580 7608
rect 39632 7568 522580 7596
rect 39632 7556 39638 7568
rect 522574 7556 522580 7568
rect 522632 7556 522638 7608
rect 359458 6808 359464 6860
rect 359516 6848 359522 6860
rect 580166 6848 580172 6860
rect 359516 6820 580172 6848
rect 359516 6808 359522 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 7558 6644 7564 6656
rect 3476 6616 7564 6644
rect 3476 6604 3482 6616
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 32398 6128 32404 6180
rect 32456 6168 32462 6180
rect 491570 6168 491576 6180
rect 32456 6140 491576 6168
rect 32456 6128 32462 6140
rect 491570 6128 491576 6140
rect 491628 6128 491634 6180
rect 208578 4836 208584 4888
rect 208636 4876 208642 4888
rect 340966 4876 340972 4888
rect 208636 4848 340972 4876
rect 208636 4836 208642 4848
rect 340966 4836 340972 4848
rect 341024 4836 341030 4888
rect 357526 4836 357532 4888
rect 357584 4876 357590 4888
rect 517974 4876 517980 4888
rect 357584 4848 517980 4876
rect 357584 4836 357590 4848
rect 517974 4836 517980 4848
rect 518032 4836 518038 4888
rect 50154 4768 50160 4820
rect 50212 4808 50218 4820
rect 508314 4808 508320 4820
rect 50212 4780 508320 4808
rect 50212 4768 50218 4780
rect 508314 4768 508320 4780
rect 508372 4768 508378 4820
rect 332686 4088 332692 4140
rect 332744 4128 332750 4140
rect 350626 4128 350632 4140
rect 332744 4100 350632 4128
rect 332744 4088 332750 4100
rect 350626 4088 350632 4100
rect 350684 4088 350690 4140
rect 499390 4088 499396 4140
rect 499448 4128 499454 4140
rect 500218 4128 500224 4140
rect 499448 4100 500224 4128
rect 499448 4088 499454 4100
rect 500218 4088 500224 4100
rect 500276 4088 500282 4140
rect 336274 4020 336280 4072
rect 336332 4060 336338 4072
rect 355410 4060 355416 4072
rect 336332 4032 355416 4060
rect 336332 4020 336338 4032
rect 355410 4020 355416 4032
rect 355468 4020 355474 4072
rect 325602 3952 325608 4004
rect 325660 3992 325666 4004
rect 350534 3992 350540 4004
rect 325660 3964 350540 3992
rect 325660 3952 325666 3964
rect 350534 3952 350540 3964
rect 350592 3952 350598 4004
rect 322106 3884 322112 3936
rect 322164 3924 322170 3936
rect 350718 3924 350724 3936
rect 322164 3896 350724 3924
rect 322164 3884 322170 3896
rect 350718 3884 350724 3896
rect 350776 3884 350782 3936
rect 307938 3816 307944 3868
rect 307996 3856 308002 3868
rect 355318 3856 355324 3868
rect 307996 3828 355324 3856
rect 307996 3816 308002 3828
rect 355318 3816 355324 3828
rect 355376 3816 355382 3868
rect 361114 3816 361120 3868
rect 361172 3856 361178 3868
rect 404998 3856 405004 3868
rect 361172 3828 405004 3856
rect 361172 3816 361178 3828
rect 404998 3816 405004 3828
rect 405056 3816 405062 3868
rect 117590 3748 117596 3800
rect 117648 3788 117654 3800
rect 406378 3788 406384 3800
rect 117648 3760 406384 3788
rect 117648 3748 117654 3760
rect 406378 3748 406384 3760
rect 406436 3748 406442 3800
rect 124674 3680 124680 3732
rect 124732 3720 124738 3732
rect 475378 3720 475384 3732
rect 124732 3692 475384 3720
rect 124732 3680 124738 3692
rect 475378 3680 475384 3692
rect 475436 3680 475442 3732
rect 491294 3680 491300 3732
rect 491352 3720 491358 3732
rect 491938 3720 491944 3732
rect 491352 3692 491944 3720
rect 491352 3680 491358 3692
rect 491938 3680 491944 3692
rect 491996 3680 492002 3732
rect 46658 3612 46664 3664
rect 46716 3652 46722 3664
rect 403710 3652 403716 3664
rect 46716 3624 403716 3652
rect 46716 3612 46722 3624
rect 403710 3612 403716 3624
rect 403768 3612 403774 3664
rect 478138 3612 478144 3664
rect 478196 3652 478202 3664
rect 518158 3652 518164 3664
rect 478196 3624 518164 3652
rect 478196 3612 478202 3624
rect 518158 3612 518164 3624
rect 518216 3612 518222 3664
rect 540238 3612 540244 3664
rect 540296 3652 540302 3664
rect 582190 3652 582196 3664
rect 540296 3624 582196 3652
rect 540296 3612 540302 3624
rect 582190 3612 582196 3624
rect 582248 3612 582254 3664
rect 28902 3544 28908 3596
rect 28960 3584 28966 3596
rect 410518 3584 410524 3596
rect 28960 3556 410524 3584
rect 28960 3544 28966 3556
rect 410518 3544 410524 3556
rect 410576 3544 410582 3596
rect 415394 3544 415400 3596
rect 415452 3584 415458 3596
rect 416682 3584 416688 3596
rect 415452 3556 416688 3584
rect 415452 3544 415458 3556
rect 416682 3544 416688 3556
rect 416740 3544 416746 3596
rect 423674 3544 423680 3596
rect 423732 3584 423738 3596
rect 424962 3584 424968 3596
rect 423732 3556 424968 3584
rect 423732 3544 423738 3556
rect 424962 3544 424968 3556
rect 425020 3544 425026 3596
rect 440234 3544 440240 3596
rect 440292 3584 440298 3596
rect 441522 3584 441528 3596
rect 440292 3556 441528 3584
rect 440292 3544 440298 3556
rect 441522 3544 441528 3556
rect 441580 3544 441586 3596
rect 449802 3544 449808 3596
rect 449860 3584 449866 3596
rect 516778 3584 516784 3596
rect 449860 3556 516784 3584
rect 449860 3544 449866 3556
rect 516778 3544 516784 3556
rect 516836 3544 516842 3596
rect 525058 3544 525064 3596
rect 525116 3584 525122 3596
rect 531314 3584 531320 3596
rect 525116 3556 531320 3584
rect 525116 3544 525122 3556
rect 531314 3544 531320 3556
rect 531372 3544 531378 3596
rect 536098 3544 536104 3596
rect 536156 3584 536162 3596
rect 573910 3584 573916 3596
rect 536156 3556 573916 3584
rect 536156 3544 536162 3556
rect 573910 3544 573916 3556
rect 573968 3544 573974 3596
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 59998 3516 60004 3528
rect 57296 3488 60004 3516
rect 57296 3476 57302 3488
rect 59998 3476 60004 3488
rect 60056 3476 60062 3528
rect 102134 3476 102140 3528
rect 102192 3516 102198 3528
rect 103330 3516 103336 3528
rect 102192 3488 103336 3516
rect 102192 3476 102198 3488
rect 103330 3476 103336 3488
rect 103388 3476 103394 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 491294 3516 491300 3528
rect 106976 3488 491300 3516
rect 106976 3476 106982 3488
rect 491294 3476 491300 3488
rect 491352 3476 491358 3528
rect 526438 3476 526444 3528
rect 526496 3516 526502 3528
rect 527818 3516 527824 3528
rect 526496 3488 527824 3516
rect 526496 3476 526502 3488
rect 527818 3476 527824 3488
rect 527876 3476 527882 3528
rect 527910 3476 527916 3528
rect 527968 3516 527974 3528
rect 538398 3516 538404 3528
rect 527968 3488 538404 3516
rect 527968 3476 527974 3488
rect 538398 3476 538404 3488
rect 538456 3476 538462 3528
rect 538858 3476 538864 3528
rect 538916 3516 538922 3528
rect 538916 3488 578832 3516
rect 538916 3476 538922 3488
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 31018 3448 31024 3460
rect 19484 3420 31024 3448
rect 19484 3408 19490 3420
rect 31018 3408 31024 3420
rect 31076 3408 31082 3460
rect 35986 3408 35992 3460
rect 36044 3448 36050 3460
rect 48958 3448 48964 3460
rect 36044 3420 48964 3448
rect 36044 3408 36050 3420
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 89162 3408 89168 3460
rect 89220 3448 89226 3460
rect 489178 3448 489184 3460
rect 89220 3420 489184 3448
rect 89220 3408 89226 3420
rect 489178 3408 489184 3420
rect 489236 3408 489242 3460
rect 504450 3408 504456 3460
rect 504508 3448 504514 3460
rect 577406 3448 577412 3460
rect 504508 3420 577412 3448
rect 504508 3408 504514 3420
rect 577406 3408 577412 3420
rect 577464 3408 577470 3460
rect 578804 3448 578832 3488
rect 578878 3476 578884 3528
rect 578936 3516 578942 3528
rect 579798 3516 579804 3528
rect 578936 3488 579804 3516
rect 578936 3476 578942 3488
rect 579798 3476 579804 3488
rect 579856 3476 579862 3528
rect 580994 3448 581000 3460
rect 578804 3420 581000 3448
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 168374 3340 168380 3392
rect 168432 3380 168438 3392
rect 169570 3380 169576 3392
rect 168432 3352 169576 3380
rect 168432 3340 168438 3352
rect 169570 3340 169576 3352
rect 169628 3340 169634 3392
rect 193214 3340 193220 3392
rect 193272 3380 193278 3392
rect 194410 3380 194416 3392
rect 193272 3352 194416 3380
rect 193272 3340 193278 3352
rect 194410 3340 194416 3352
rect 194468 3340 194474 3392
rect 218054 3340 218060 3392
rect 218112 3380 218118 3392
rect 219250 3380 219256 3392
rect 218112 3352 219256 3380
rect 218112 3340 218118 3352
rect 219250 3340 219256 3352
rect 219308 3340 219314 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 339862 3340 339868 3392
rect 339920 3380 339926 3392
rect 339920 3352 349108 3380
rect 339920 3340 339926 3352
rect 349080 3312 349108 3352
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474182 3380 474188 3392
rect 473412 3352 474188 3380
rect 473412 3340 473418 3352
rect 474182 3340 474188 3352
rect 474240 3340 474246 3392
rect 558178 3340 558184 3392
rect 558236 3380 558242 3392
rect 559742 3380 559748 3392
rect 558236 3352 559748 3380
rect 558236 3340 558242 3352
rect 559742 3340 559748 3352
rect 559800 3340 559806 3392
rect 353478 3312 353484 3324
rect 349080 3284 353484 3312
rect 353478 3272 353484 3284
rect 353536 3272 353542 3324
rect 343358 3204 343364 3256
rect 343416 3244 343422 3256
rect 353386 3244 353392 3256
rect 343416 3216 353392 3244
rect 343416 3204 343422 3216
rect 353386 3204 353392 3216
rect 353444 3204 353450 3256
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 235172 700612 235224 700664
rect 253204 700612 253256 700664
rect 202788 700544 202840 700596
rect 253296 700544 253348 700596
rect 348792 700544 348844 700596
rect 409236 700544 409288 700596
rect 154120 700476 154172 700528
rect 260104 700476 260156 700528
rect 405004 700476 405056 700528
rect 559656 700476 559708 700528
rect 137836 700408 137888 700460
rect 253388 700408 253440 700460
rect 317420 700408 317472 700460
rect 543464 700408 543516 700460
rect 89168 700340 89220 700392
rect 406476 700340 406528 700392
rect 24308 700272 24360 700324
rect 472716 700272 472768 700324
rect 526444 699660 526496 699712
rect 527180 699660 527232 699712
rect 397460 698912 397512 698964
rect 458824 698912 458876 698964
rect 105452 697552 105504 697604
rect 337384 697552 337436 697604
rect 525064 696940 525116 696992
rect 580172 696940 580224 696992
rect 267648 694764 267700 694816
rect 427084 694764 427136 694816
rect 316132 683136 316184 683188
rect 580172 683136 580224 683188
rect 403716 670692 403768 670744
rect 580172 670692 580224 670744
rect 3240 667156 3292 667208
rect 479524 667156 479576 667208
rect 40040 665796 40092 665848
rect 476948 665796 477000 665848
rect 46572 663756 46624 663808
rect 352840 663756 352892 663808
rect 52000 663144 52052 663196
rect 276664 663144 276716 663196
rect 51908 663076 51960 663128
rect 276756 663076 276808 663128
rect 46664 663008 46716 663060
rect 276848 663008 276900 663060
rect 52184 662940 52236 662992
rect 353024 662940 353076 662992
rect 51172 662872 51224 662924
rect 352656 662872 352708 662924
rect 47860 662804 47912 662856
rect 349804 662804 349856 662856
rect 51080 662736 51132 662788
rect 355416 662736 355468 662788
rect 50988 662668 51040 662720
rect 355324 662668 355376 662720
rect 46480 662600 46532 662652
rect 352748 662600 352800 662652
rect 45468 662532 45520 662584
rect 352564 662532 352616 662584
rect 51816 662464 51868 662516
rect 403256 662464 403308 662516
rect 46388 662396 46440 662448
rect 405280 662396 405332 662448
rect 52092 661784 52144 661836
rect 279516 661784 279568 661836
rect 218060 661716 218112 661768
rect 521844 661716 521896 661768
rect 6920 661648 6972 661700
rect 520740 661648 520792 661700
rect 48872 661580 48924 661632
rect 279608 661580 279660 661632
rect 48504 661512 48556 661564
rect 310520 661512 310572 661564
rect 50896 661444 50948 661496
rect 356704 661444 356756 661496
rect 50804 661376 50856 661428
rect 358820 661376 358872 661428
rect 50620 661308 50672 661360
rect 401600 661308 401652 661360
rect 51724 661240 51776 661292
rect 407120 661240 407172 661292
rect 50344 661172 50396 661224
rect 478328 661172 478380 661224
rect 50528 661104 50580 661156
rect 478420 661104 478472 661156
rect 3516 661036 3568 661088
rect 522028 661036 522080 661088
rect 49608 660560 49660 660612
rect 278136 660560 278188 660612
rect 50712 660492 50764 660544
rect 279700 660492 279752 660544
rect 50436 660424 50488 660476
rect 502340 660424 502392 660476
rect 49424 660356 49476 660408
rect 279148 660356 279200 660408
rect 331220 660356 331272 660408
rect 520464 660356 520516 660408
rect 49884 660288 49936 660340
rect 507860 660288 507912 660340
rect 49516 660220 49568 660272
rect 280068 660220 280120 660272
rect 48136 660152 48188 660204
rect 279332 660152 279384 660204
rect 48044 660084 48096 660136
rect 279240 660084 279292 660136
rect 48228 660016 48280 660068
rect 279884 660016 279936 660068
rect 50252 659948 50304 660000
rect 521660 659948 521712 660000
rect 3424 659880 3476 659932
rect 478972 659880 479024 659932
rect 3332 659812 3384 659864
rect 520372 659812 520424 659864
rect 49976 657976 50028 658028
rect 50252 657976 50304 658028
rect 50528 657500 50580 657552
rect 50896 657500 50948 657552
rect 49332 655052 49384 655104
rect 49608 655052 49660 655104
rect 48688 652740 48740 652792
rect 50160 652740 50212 652792
rect 50988 651380 51040 651432
rect 52184 651380 52236 651432
rect 49424 648524 49476 648576
rect 50068 648524 50120 648576
rect 254308 645872 254360 645924
rect 257344 645872 257396 645924
rect 282920 643696 282972 643748
rect 477040 643696 477092 643748
rect 534724 643084 534776 643136
rect 580172 643084 580224 643136
rect 360936 642676 360988 642728
rect 379428 642676 379480 642728
rect 370044 642608 370096 642660
rect 403808 642608 403860 642660
rect 359556 642540 359608 642592
rect 376116 642540 376168 642592
rect 392676 642540 392728 642592
rect 400772 642540 400824 642592
rect 327724 642472 327776 642524
rect 377772 642472 377824 642524
rect 389916 642472 389968 642524
rect 399484 642472 399536 642524
rect 371148 642404 371200 642456
rect 405372 642404 405424 642456
rect 287612 642336 287664 642388
rect 349896 642336 349948 642388
rect 360844 642336 360896 642388
rect 396540 642336 396592 642388
rect 293776 642268 293828 642320
rect 321192 642268 321244 642320
rect 359464 642268 359516 642320
rect 373356 642268 373408 642320
rect 373908 642268 373960 642320
rect 400864 642268 400916 642320
rect 300768 642200 300820 642252
rect 331864 642200 331916 642252
rect 358820 642200 358872 642252
rect 388260 642200 388312 642252
rect 394332 642200 394384 642252
rect 405188 642200 405240 642252
rect 295248 642132 295300 642184
rect 329104 642132 329156 642184
rect 359740 642132 359792 642184
rect 390468 642132 390520 642184
rect 393228 642132 393280 642184
rect 400680 642132 400732 642184
rect 286508 642064 286560 642116
rect 322296 642064 322348 642116
rect 357348 642064 357400 642116
rect 388812 642064 388864 642116
rect 392124 642064 392176 642116
rect 400404 642064 400456 642116
rect 282092 641996 282144 642048
rect 319536 641996 319588 642048
rect 353116 641996 353168 642048
rect 386604 641996 386656 642048
rect 387708 641996 387760 642048
rect 399576 641996 399628 642048
rect 282736 641928 282788 641980
rect 321008 641928 321060 641980
rect 355968 641928 356020 641980
rect 391020 641928 391072 641980
rect 284208 641860 284260 641912
rect 327816 641860 327868 641912
rect 360016 641860 360068 641912
rect 371700 641860 371752 641912
rect 375288 641860 375340 641912
rect 389364 641860 389416 641912
rect 394884 641860 394936 641912
rect 400588 641860 400640 641912
rect 297548 641792 297600 641844
rect 352932 641792 352984 641844
rect 358912 641792 358964 641844
rect 366732 641792 366784 641844
rect 379520 641792 379572 641844
rect 386052 641792 386104 641844
rect 393780 641792 393832 641844
rect 399300 641792 399352 641844
rect 475384 641792 475436 641844
rect 493232 641792 493284 641844
rect 49148 641724 49200 641776
rect 50252 641724 50304 641776
rect 299296 641724 299348 641776
rect 321100 641724 321152 641776
rect 349988 641724 350040 641776
rect 363420 641724 363472 641776
rect 367008 641724 367060 641776
rect 372252 641724 372304 641776
rect 378048 641724 378100 641776
rect 384396 641724 384448 641776
rect 395436 641724 395488 641776
rect 399668 641724 399720 641776
rect 406384 641724 406436 641776
rect 510620 641724 510672 641776
rect 278688 640976 278740 641028
rect 310060 640976 310112 641028
rect 315856 640976 315908 641028
rect 523684 640976 523736 641028
rect 314108 640908 314160 640960
rect 527824 640908 527876 640960
rect 359832 640840 359884 640892
rect 381636 640840 381688 640892
rect 355508 640772 355560 640824
rect 378324 640772 378376 640824
rect 357072 640704 357124 640756
rect 384948 640704 385000 640756
rect 313004 640636 313056 640688
rect 338764 640636 338816 640688
rect 372804 640636 372856 640688
rect 400312 640636 400364 640688
rect 309692 640568 309744 640620
rect 356980 640568 357032 640620
rect 357164 640568 357216 640620
rect 385500 640568 385552 640620
rect 304816 640500 304868 640552
rect 354036 640500 354088 640552
rect 354128 640500 354180 640552
rect 383844 640500 383896 640552
rect 387156 640500 387208 640552
rect 402336 640500 402388 640552
rect 254308 640432 254360 640484
rect 257436 640432 257488 640484
rect 301964 640432 302016 640484
rect 356796 640432 356848 640484
rect 364524 640432 364576 640484
rect 400220 640432 400272 640484
rect 315212 640364 315264 640416
rect 322388 640364 322440 640416
rect 361212 640364 361264 640416
rect 379980 640364 380032 640416
rect 310336 640296 310388 640348
rect 320824 640296 320876 640348
rect 361120 640296 361172 640348
rect 382740 640296 382792 640348
rect 364984 639888 365036 639940
rect 365260 639888 365312 639940
rect 358636 639752 358688 639804
rect 367008 639820 367060 639872
rect 358452 639684 358504 639736
rect 375288 639752 375340 639804
rect 362224 639684 362276 639736
rect 374644 639684 374696 639736
rect 367560 639616 367612 639668
rect 372528 639616 372580 639668
rect 357808 639548 357860 639600
rect 376300 639548 376352 639600
rect 361488 639480 361540 639532
rect 370228 639480 370280 639532
rect 296444 639276 296496 639328
rect 303068 639344 303120 639396
rect 306288 639276 306340 639328
rect 360108 639412 360160 639464
rect 368204 639412 368256 639464
rect 358544 639344 358596 639396
rect 362224 639344 362276 639396
rect 364984 639344 365036 639396
rect 365352 639344 365404 639396
rect 366456 639344 366508 639396
rect 311716 639276 311768 639328
rect 324964 639276 325016 639328
rect 322204 639140 322256 639192
rect 353944 639072 353996 639124
rect 356888 639004 356940 639056
rect 278780 638936 278832 638988
rect 361580 638936 361632 638988
rect 369676 639344 369728 639396
rect 374736 639412 374788 639464
rect 372528 639344 372580 639396
rect 375840 639344 375892 639396
rect 377496 639412 377548 639464
rect 399116 639616 399168 639668
rect 396172 639548 396224 639600
rect 399024 639548 399076 639600
rect 391204 639480 391256 639532
rect 404636 639480 404688 639532
rect 391204 639344 391256 639396
rect 397920 639412 397972 639464
rect 398932 639412 398984 639464
rect 403164 639276 403216 639328
rect 399944 639208 399996 639260
rect 400496 639140 400548 639192
rect 403900 639072 403952 639124
rect 402152 639004 402204 639056
rect 401784 638936 401836 638988
rect 403624 634788 403676 634840
rect 477684 634788 477736 634840
rect 254676 633428 254728 633480
rect 269856 633428 269908 633480
rect 523684 632000 523736 632052
rect 580172 632000 580224 632052
rect 49332 629688 49384 629740
rect 52092 629688 52144 629740
rect 254676 627920 254728 627972
rect 275376 627920 275428 627972
rect 48872 618944 48924 618996
rect 52000 618944 52052 618996
rect 254400 616836 254452 616888
rect 264244 616836 264296 616888
rect 538864 616836 538916 616888
rect 580172 616836 580224 616888
rect 48780 612756 48832 612808
rect 51908 612756 51960 612808
rect 254492 611328 254544 611380
rect 273904 611328 273956 611380
rect 254216 604460 254268 604512
rect 271144 604460 271196 604512
rect 398380 600244 398432 600296
rect 403624 600244 403676 600296
rect 391940 599972 391992 600024
rect 392308 599972 392360 600024
rect 301964 599904 302016 599956
rect 302194 599904 302246 599956
rect 296720 599836 296772 599888
rect 297778 599836 297830 599888
rect 298100 599836 298152 599888
rect 299434 599836 299486 599888
rect 392308 599836 392360 599888
rect 399208 599836 399260 599888
rect 382280 599768 382332 599820
rect 400588 599768 400640 599820
rect 378508 599700 378560 599752
rect 400772 599700 400824 599752
rect 372620 599632 372672 599684
rect 399300 599632 399352 599684
rect 254584 599564 254636 599616
rect 320180 599564 320232 599616
rect 365720 599564 365772 599616
rect 400680 599564 400732 599616
rect 297824 599224 297876 599276
rect 327724 599224 327776 599276
rect 300860 599156 300912 599208
rect 301964 599156 302016 599208
rect 331956 599156 332008 599208
rect 306380 599088 306432 599140
rect 306748 599088 306800 599140
rect 353116 599088 353168 599140
rect 387708 599088 387760 599140
rect 406384 599088 406436 599140
rect 299388 599020 299440 599072
rect 360936 599020 360988 599072
rect 361764 599020 361816 599072
rect 475384 599020 475436 599072
rect 283012 598952 283064 599004
rect 349988 598952 350040 599004
rect 254768 598884 254820 598936
rect 386604 598952 386656 599004
rect 387708 598952 387760 599004
rect 388260 598884 388312 598936
rect 521752 598884 521804 598936
rect 302148 598816 302200 598868
rect 303528 598748 303580 598800
rect 311256 598816 311308 598868
rect 361212 598816 361264 598868
rect 386420 598816 386472 598868
rect 387156 598816 387208 598868
rect 513840 598816 513892 598868
rect 359832 598748 359884 598800
rect 388444 598748 388496 598800
rect 478144 598748 478196 598800
rect 361120 598680 361172 598732
rect 286876 598612 286928 598664
rect 289176 598612 289228 598664
rect 292488 598612 292540 598664
rect 297456 598612 297508 598664
rect 304908 598612 304960 598664
rect 357072 598612 357124 598664
rect 361028 598612 361080 598664
rect 380532 598612 380584 598664
rect 285128 598408 285180 598460
rect 305828 598544 305880 598596
rect 306288 598544 306340 598596
rect 357164 598544 357216 598596
rect 359648 598544 359700 598596
rect 382188 598544 382240 598596
rect 388260 598544 388312 598596
rect 388536 598544 388588 598596
rect 304172 598476 304224 598528
rect 354128 598476 354180 598528
rect 360936 598476 360988 598528
rect 391572 598476 391624 598528
rect 320916 598408 320968 598460
rect 366180 598408 366232 598460
rect 397736 598408 397788 598460
rect 288992 598340 289044 598392
rect 290096 598204 290148 598256
rect 297456 598340 297508 598392
rect 303068 598340 303120 598392
rect 303528 598340 303580 598392
rect 303620 598340 303672 598392
rect 355508 598340 355560 598392
rect 363420 598340 363472 598392
rect 398104 598340 398156 598392
rect 404728 598272 404780 598324
rect 287060 598136 287112 598188
rect 287520 598136 287572 598188
rect 291108 598136 291160 598188
rect 291844 598136 291896 598188
rect 404820 598204 404872 598256
rect 472808 598204 472860 598256
rect 496452 598204 496504 598256
rect 323676 598136 323728 598188
rect 369860 598136 369912 598188
rect 370228 598136 370280 598188
rect 372712 598136 372764 598188
rect 373540 598136 373592 598188
rect 378416 598136 378468 598188
rect 379060 598136 379112 598188
rect 380992 598136 381044 598188
rect 381268 598136 381320 598188
rect 389272 598136 389324 598188
rect 389548 598136 389600 598188
rect 393320 598136 393372 598188
rect 393964 598136 394016 598188
rect 396080 598136 396132 598188
rect 396724 598136 396776 598188
rect 298652 598068 298704 598120
rect 300676 598068 300728 598120
rect 303620 598068 303672 598120
rect 304172 598068 304224 598120
rect 304816 598068 304868 598120
rect 306472 598068 306524 598120
rect 307392 598068 307444 598120
rect 309140 598068 309192 598120
rect 310152 598068 310204 598120
rect 311900 598068 311952 598120
rect 312360 598068 312412 598120
rect 313280 598068 313332 598120
rect 314016 598068 314068 598120
rect 314660 598068 314712 598120
rect 315120 598068 315172 598120
rect 389180 598068 389232 598120
rect 390100 598068 390152 598120
rect 392032 598068 392084 598120
rect 392860 598068 392912 598120
rect 300308 598000 300360 598052
rect 300584 598000 300636 598052
rect 311256 598000 311308 598052
rect 314752 598000 314804 598052
rect 315672 598000 315724 598052
rect 308312 597932 308364 597984
rect 323584 597932 323636 597984
rect 395436 597796 395488 597848
rect 400588 597796 400640 597848
rect 362868 597524 362920 597576
rect 368664 597524 368716 597576
rect 383660 597184 383712 597236
rect 384580 597184 384632 597236
rect 282920 597048 282972 597100
rect 283656 597048 283708 597100
rect 313188 596912 313240 596964
rect 337476 596912 337528 596964
rect 347688 596912 347740 596964
rect 375564 596912 375616 596964
rect 253388 596844 253440 596896
rect 502340 596844 502392 596896
rect 325608 596776 325660 596828
rect 398196 596776 398248 596828
rect 468668 596776 468720 596828
rect 479708 596776 479760 596828
rect 367284 596368 367336 596420
rect 367284 596164 367336 596216
rect 320180 596096 320232 596148
rect 325608 596096 325660 596148
rect 292580 596028 292632 596080
rect 293592 596028 293644 596080
rect 364432 596028 364484 596080
rect 365260 596028 365312 596080
rect 367100 596028 367152 596080
rect 368020 596028 368072 596080
rect 297548 595484 297600 595536
rect 341524 595484 341576 595536
rect 349988 595484 350040 595536
rect 363972 595484 364024 595536
rect 372896 595484 372948 595536
rect 383844 595484 383896 595536
rect 253296 595416 253348 595468
rect 503720 595416 503772 595468
rect 383936 595212 383988 595264
rect 392584 595212 392636 595264
rect 49516 594804 49568 594856
rect 51724 594804 51776 594856
rect 307024 594124 307076 594176
rect 327724 594124 327776 594176
rect 343548 594124 343600 594176
rect 371792 594124 371844 594176
rect 288440 594056 288492 594108
rect 345664 594056 345716 594108
rect 371884 594056 371936 594108
rect 391940 594056 391992 594108
rect 254492 593376 254544 593428
rect 275284 593376 275336 593428
rect 311992 592696 312044 592748
rect 322480 592696 322532 592748
rect 254860 592628 254912 592680
rect 269764 592628 269816 592680
rect 293500 592628 293552 592680
rect 347044 592628 347096 592680
rect 385684 592016 385736 592068
rect 389180 592016 389232 592068
rect 306840 591336 306892 591388
rect 334624 591336 334676 591388
rect 336096 591336 336148 591388
rect 396172 591336 396224 591388
rect 260104 591268 260156 591320
rect 480260 591268 480312 591320
rect 478788 590656 478840 590708
rect 579804 590656 579856 590708
rect 47860 590588 47912 590640
rect 48964 590588 49016 590640
rect 329748 589976 329800 590028
rect 364708 589976 364760 590028
rect 381544 589976 381596 590028
rect 386420 589976 386472 590028
rect 294604 589908 294656 589960
rect 386788 589908 386840 589960
rect 367192 589432 367244 589484
rect 367376 589432 367428 589484
rect 314844 588616 314896 588668
rect 338856 588616 338908 588668
rect 342168 588616 342220 588668
rect 367192 588616 367244 588668
rect 291384 588548 291436 588600
rect 350080 588548 350132 588600
rect 254584 587936 254636 587988
rect 260104 587936 260156 587988
rect 333888 587188 333940 587240
rect 368572 587188 368624 587240
rect 287980 587120 288032 587172
rect 342904 587120 342956 587172
rect 304724 585828 304776 585880
rect 340144 585828 340196 585880
rect 361120 585828 361172 585880
rect 392124 585828 392176 585880
rect 331956 585760 332008 585812
rect 372804 585760 372856 585812
rect 310612 584400 310664 584452
rect 345756 584400 345808 584452
rect 293960 581612 294012 581664
rect 367192 581612 367244 581664
rect 253940 581272 253992 581324
rect 255964 581272 256016 581324
rect 319444 580252 319496 580304
rect 475568 580252 475620 580304
rect 329104 578892 329156 578944
rect 382464 578892 382516 578944
rect 322388 578144 322440 578196
rect 580172 578144 580224 578196
rect 303436 577532 303488 577584
rect 336004 577532 336056 577584
rect 321192 577464 321244 577516
rect 379520 577464 379572 577516
rect 287060 576172 287112 576224
rect 354220 576172 354272 576224
rect 306472 576104 306524 576156
rect 389272 576104 389324 576156
rect 254216 575492 254268 575544
rect 278044 575492 278096 575544
rect 327816 574812 327868 574864
rect 396172 574812 396224 574864
rect 304816 574744 304868 574796
rect 394884 574744 394936 574796
rect 296720 573384 296772 573436
rect 367376 573384 367428 573436
rect 314752 573316 314804 573368
rect 390652 573316 390704 573368
rect 285680 572024 285732 572076
rect 353116 572024 353168 572076
rect 319536 571956 319588 572008
rect 522120 571956 522172 572008
rect 310520 570664 310572 570716
rect 374276 570664 374328 570716
rect 284392 570596 284444 570648
rect 386604 570596 386656 570648
rect 253940 569984 253992 570036
rect 256056 569984 256108 570036
rect 292580 569168 292632 569220
rect 357072 569168 357124 569220
rect 307760 567876 307812 567928
rect 368572 567876 368624 567928
rect 289084 567808 289136 567860
rect 386696 567808 386748 567860
rect 388536 567196 388588 567248
rect 393412 567196 393464 567248
rect 3332 567128 3384 567180
rect 50436 567128 50488 567180
rect 313372 566448 313424 566500
rect 376852 566448 376904 566500
rect 372712 565836 372764 565888
rect 404912 565836 404964 565888
rect 350448 565224 350500 565276
rect 372712 565224 372764 565276
rect 306196 565156 306248 565208
rect 365904 565156 365956 565208
rect 283012 565088 283064 565140
rect 354312 565088 354364 565140
rect 358268 565088 358320 565140
rect 396080 565088 396132 565140
rect 254584 564408 254636 564460
rect 279424 564408 279476 564460
rect 359096 563796 359148 563848
rect 386512 563796 386564 563848
rect 358360 563728 358412 563780
rect 394700 563728 394752 563780
rect 300768 563660 300820 563712
rect 362960 563660 363012 563712
rect 321100 562368 321152 562420
rect 401968 562368 402020 562420
rect 253204 562300 253256 562352
rect 381084 562300 381136 562352
rect 321008 560940 321060 560992
rect 402060 560940 402112 560992
rect 384304 560736 384356 560788
rect 390744 560736 390796 560788
rect 363236 559648 363288 559700
rect 374092 559648 374144 559700
rect 364432 559580 364484 559632
rect 376668 559580 376720 559632
rect 396080 559580 396132 559632
rect 316132 559512 316184 559564
rect 400956 559512 401008 559564
rect 359004 558220 359056 558272
rect 380992 558220 381044 558272
rect 291844 558152 291896 558204
rect 375472 558152 375524 558204
rect 376760 558152 376812 558204
rect 377128 558152 377180 558204
rect 254584 557540 254636 557592
rect 265624 557540 265676 557592
rect 357900 556860 357952 556912
rect 381176 556860 381228 556912
rect 362592 556792 362644 556844
rect 374000 556792 374052 556844
rect 378048 556792 378100 556844
rect 538864 556792 538916 556844
rect 365812 556180 365864 556232
rect 371332 556180 371384 556232
rect 359188 555500 359240 555552
rect 385132 555500 385184 555552
rect 284300 555432 284352 555484
rect 399852 555432 399904 555484
rect 369952 554820 370004 554872
rect 402980 554820 403032 554872
rect 367100 554752 367152 554804
rect 404544 554752 404596 554804
rect 2964 554684 3016 554736
rect 50344 554684 50396 554736
rect 355600 554208 355652 554260
rect 367100 554208 367152 554260
rect 355784 554140 355836 554192
rect 369952 554140 370004 554192
rect 322296 554072 322348 554124
rect 401876 554072 401928 554124
rect 314660 554004 314712 554056
rect 401232 554004 401284 554056
rect 392584 553324 392636 553376
rect 394148 553324 394200 553376
rect 385040 553256 385092 553308
rect 392216 553256 392268 553308
rect 389272 553052 389324 553104
rect 399116 553052 399168 553104
rect 360108 552916 360160 552968
rect 378692 552916 378744 552968
rect 383752 552916 383804 552968
rect 400036 552916 400088 552968
rect 347136 552780 347188 552832
rect 368664 552848 368716 552900
rect 388352 552848 388404 552900
rect 379980 552780 380032 552832
rect 400404 552780 400456 552832
rect 356704 552712 356756 552764
rect 396724 552712 396776 552764
rect 309232 552644 309284 552696
rect 360660 552644 360712 552696
rect 361488 552644 361540 552696
rect 374184 552644 374236 552696
rect 376116 552644 376168 552696
rect 399024 552644 399076 552696
rect 399484 552644 399536 552696
rect 402428 552644 402480 552696
rect 393504 552508 393556 552560
rect 400496 552508 400548 552560
rect 355232 552304 355284 552356
rect 361120 552304 361172 552356
rect 375656 552304 375708 552356
rect 403440 552304 403492 552356
rect 356612 552236 356664 552288
rect 385684 552236 385736 552288
rect 398656 552236 398708 552288
rect 409144 552236 409196 552288
rect 354404 552168 354456 552220
rect 384304 552168 384356 552220
rect 394792 552168 394844 552220
rect 430580 552168 430632 552220
rect 357164 552100 357216 552152
rect 371884 552100 371936 552152
rect 373540 552100 373592 552152
rect 498844 552100 498896 552152
rect 254584 552032 254636 552084
rect 268384 552032 268436 552084
rect 348424 552032 348476 552084
rect 381544 552032 381596 552084
rect 391204 552032 391256 552084
rect 391572 552032 391624 552084
rect 520556 552032 520608 552084
rect 398104 551964 398156 552016
rect 401600 551964 401652 552016
rect 375012 551896 375064 551948
rect 375656 551896 375708 551948
rect 358084 551692 358136 551744
rect 360936 551692 360988 551744
rect 389456 551692 389508 551744
rect 399760 551692 399812 551744
rect 355140 551624 355192 551676
rect 377128 551624 377180 551676
rect 400772 551624 400824 551676
rect 322388 551556 322440 551608
rect 376668 551556 376720 551608
rect 383660 551556 383712 551608
rect 399484 551556 399536 551608
rect 304632 551488 304684 551540
rect 403072 551488 403124 551540
rect 295524 551420 295576 551472
rect 403348 551420 403400 551472
rect 295340 551352 295392 551404
rect 403532 551352 403584 551404
rect 295432 551284 295484 551336
rect 404452 551284 404504 551336
rect 358176 551216 358228 551268
rect 361028 551216 361080 551268
rect 363144 551216 363196 551268
rect 363604 551216 363656 551268
rect 382280 551216 382332 551268
rect 382924 551216 382976 551268
rect 364340 551080 364392 551132
rect 365168 551080 365220 551132
rect 351276 550808 351328 550860
rect 388536 550808 388588 550860
rect 388996 550808 389048 550860
rect 358728 550740 358780 550792
rect 360844 550740 360896 550792
rect 367100 550740 367152 550792
rect 419540 550740 419592 550792
rect 341616 550672 341668 550724
rect 342168 550672 342220 550724
rect 404360 550672 404412 550724
rect 351184 550604 351236 550656
rect 364340 550604 364392 550656
rect 369032 550604 369084 550656
rect 448520 550604 448572 550656
rect 386604 550536 386656 550588
rect 387064 550536 387116 550588
rect 399668 550536 399720 550588
rect 401692 550536 401744 550588
rect 393320 550468 393372 550520
rect 400496 550468 400548 550520
rect 353208 549992 353260 550044
rect 375012 550060 375064 550112
rect 355876 549992 355928 550044
rect 362960 549992 363012 550044
rect 355692 549924 355744 549976
rect 380164 550060 380216 550112
rect 383936 550060 383988 550112
rect 378784 549924 378836 549976
rect 380992 549924 381044 549976
rect 397644 550060 397696 550112
rect 397552 549992 397604 550044
rect 352380 549856 352432 549908
rect 380164 549856 380216 549908
rect 359924 549788 359976 549840
rect 362316 549788 362368 549840
rect 359832 549652 359884 549704
rect 371332 549788 371384 549840
rect 378784 549788 378836 549840
rect 352472 549516 352524 549568
rect 324228 549380 324280 549432
rect 359924 549380 359976 549432
rect 327816 549312 327868 549364
rect 359832 549312 359884 549364
rect 325516 549244 325568 549296
rect 383568 549856 383620 549908
rect 383936 549856 383988 549908
rect 400680 549856 400732 549908
rect 380992 549788 381044 549840
rect 400588 549720 400640 549772
rect 401048 549720 401100 549772
rect 400588 549516 400640 549568
rect 322296 548564 322348 548616
rect 356612 548564 356664 548616
rect 302148 548496 302200 548548
rect 357072 548496 357124 548548
rect 281540 547816 281592 547868
rect 357440 547816 357492 547868
rect 254584 546456 254636 546508
rect 261484 546456 261536 546508
rect 399576 546456 399628 546508
rect 402520 546456 402572 546508
rect 322480 546388 322532 546440
rect 357440 546388 357492 546440
rect 276848 545844 276900 545896
rect 301872 545844 301924 545896
rect 279700 545776 279752 545828
rect 312912 545776 312964 545828
rect 279608 545708 279660 545760
rect 313648 545708 313700 545760
rect 317420 545708 317472 545760
rect 332600 545708 332652 545760
rect 254676 545028 254728 545080
rect 260196 545028 260248 545080
rect 306380 545028 306432 545080
rect 357440 545028 357492 545080
rect 309140 544348 309192 544400
rect 355508 544348 355560 544400
rect 482192 544348 482244 544400
rect 525064 544348 525116 544400
rect 357624 543736 357676 543788
rect 359648 543736 359700 543788
rect 279884 543668 279936 543720
rect 298192 543668 298244 543720
rect 279332 543532 279384 543584
rect 298928 543532 298980 543584
rect 401784 543532 401836 543584
rect 402060 543532 402112 543584
rect 478972 543532 479024 543584
rect 479708 543532 479760 543584
rect 279240 543464 279292 543516
rect 299664 543464 299716 543516
rect 279516 543396 279568 543448
rect 302608 543396 302660 543448
rect 401784 543396 401836 543448
rect 404544 543396 404596 543448
rect 276756 543328 276808 543380
rect 304080 543328 304132 543380
rect 279148 543260 279200 543312
rect 316316 543260 316368 543312
rect 280068 543192 280120 543244
rect 315120 543192 315172 543244
rect 278136 543124 278188 543176
rect 316592 543124 316644 543176
rect 427820 543124 427872 543176
rect 509424 543124 509476 543176
rect 276664 543056 276716 543108
rect 303620 543056 303672 543108
rect 326344 543056 326396 543108
rect 357716 543056 357768 543108
rect 420920 543056 420972 543108
rect 513380 543056 513432 543108
rect 279976 542988 280028 543040
rect 314844 542988 314896 543040
rect 316040 542988 316092 543040
rect 354128 542988 354180 543040
rect 416780 542988 416832 543040
rect 482284 542988 482336 543040
rect 498844 542988 498896 543040
rect 512000 542988 512052 543040
rect 470600 542920 470652 542972
rect 499028 542920 499080 542972
rect 476764 542852 476816 542904
rect 506112 542852 506164 542904
rect 473360 542784 473412 542836
rect 510620 542784 510672 542836
rect 472624 542716 472676 542768
rect 515772 542716 515824 542768
rect 438860 542648 438912 542700
rect 494060 542648 494112 542700
rect 279700 542580 279752 542632
rect 279608 542512 279660 542564
rect 475476 542580 475528 542632
rect 514760 542580 514812 542632
rect 279792 542444 279844 542496
rect 292764 542512 292816 542564
rect 423680 542512 423732 542564
rect 500316 542512 500368 542564
rect 503996 542512 504048 542564
rect 540244 542512 540296 542564
rect 278320 542376 278372 542428
rect 284944 542376 284996 542428
rect 293960 542444 294012 542496
rect 478236 542444 478288 542496
rect 488172 542444 488224 542496
rect 295340 542376 295392 542428
rect 466460 542376 466512 542428
rect 484860 542376 484912 542428
rect 313280 541628 313332 541680
rect 350172 541628 350224 541680
rect 406384 541356 406436 541408
rect 493232 541356 493284 541408
rect 403624 541288 403676 541340
rect 495440 541288 495492 541340
rect 475384 541220 475436 541272
rect 511264 541220 511316 541272
rect 440884 541152 440936 541204
rect 483020 541152 483072 541204
rect 484768 541152 484820 541204
rect 543004 541152 543056 541204
rect 436836 541084 436888 541136
rect 508688 541084 508740 541136
rect 492588 541016 492640 541068
rect 556160 541016 556212 541068
rect 254400 540948 254452 541000
rect 267004 540948 267056 541000
rect 401784 540948 401836 541000
rect 437480 540948 437532 541000
rect 488080 540948 488132 541000
rect 545120 540948 545172 541000
rect 306288 540268 306340 540320
rect 347228 540268 347280 540320
rect 303528 540200 303580 540252
rect 353300 540200 353352 540252
rect 402980 539996 403032 540048
rect 500960 539996 501012 540048
rect 489828 539928 489880 539980
rect 520280 539928 520332 539980
rect 486976 539860 487028 539912
rect 547880 539860 547932 539912
rect 490656 539792 490708 539844
rect 565820 539792 565872 539844
rect 410524 539724 410576 539776
rect 496452 539724 496504 539776
rect 498200 539724 498252 539776
rect 544384 539724 544436 539776
rect 493232 539656 493284 539708
rect 525064 539656 525116 539708
rect 276664 539588 276716 539640
rect 286416 539588 286468 539640
rect 405004 539588 405056 539640
rect 518348 539588 518400 539640
rect 280804 539520 280856 539572
rect 284208 539520 284260 539572
rect 332600 539520 332652 539572
rect 357440 539520 357492 539572
rect 519636 539520 519688 539572
rect 523040 539520 523092 539572
rect 322940 537548 322992 537600
rect 358268 537548 358320 537600
rect 320180 537480 320232 537532
rect 356704 537480 356756 537532
rect 358268 536868 358320 536920
rect 358912 536868 358964 536920
rect 358452 536800 358504 536852
rect 359556 536800 359608 536852
rect 523684 536800 523736 536852
rect 580172 536800 580224 536852
rect 347044 536732 347096 536784
rect 357440 536732 357492 536784
rect 355416 536664 355468 536716
rect 357900 536664 357952 536716
rect 522212 535644 522264 535696
rect 525156 535644 525208 535696
rect 357532 535508 357584 535560
rect 354220 535372 354272 535424
rect 357532 535372 357584 535424
rect 359648 535372 359700 535424
rect 322112 535304 322164 535356
rect 352380 535304 352432 535356
rect 354312 535304 354364 535356
rect 357900 535304 357952 535356
rect 337476 535236 337528 535288
rect 357440 535236 357492 535288
rect 322480 535168 322532 535220
rect 355140 535168 355192 535220
rect 322572 534692 322624 534744
rect 337936 534692 337988 534744
rect 254584 534080 254636 534132
rect 278136 534080 278188 534132
rect 400864 534080 400916 534132
rect 402060 534080 402112 534132
rect 401600 533876 401652 533928
rect 404912 533876 404964 533928
rect 322480 533400 322532 533452
rect 329564 533400 329616 533452
rect 338028 533400 338080 533452
rect 357532 533400 357584 533452
rect 322848 533332 322900 533384
rect 357164 533332 357216 533384
rect 423036 533332 423088 533384
rect 477592 533332 477644 533384
rect 454776 532720 454828 532772
rect 477592 532720 477644 532772
rect 321652 532652 321704 532704
rect 352472 532652 352524 532704
rect 353300 532652 353352 532704
rect 357532 532652 357584 532704
rect 522948 532652 523000 532704
rect 534724 532652 534776 532704
rect 345756 532584 345808 532636
rect 357440 532584 357492 532636
rect 329564 531972 329616 532024
rect 336096 531972 336148 532024
rect 342996 531972 343048 532024
rect 463700 531292 463752 531344
rect 477592 531292 477644 531344
rect 322480 531224 322532 531276
rect 338028 531224 338080 531276
rect 458824 531224 458876 531276
rect 478696 531224 478748 531276
rect 322664 530544 322716 530596
rect 350540 530544 350592 530596
rect 401600 530204 401652 530256
rect 403532 530204 403584 530256
rect 322572 529932 322624 529984
rect 357164 529932 357216 529984
rect 401784 529932 401836 529984
rect 458180 529932 458232 529984
rect 322480 529864 322532 529916
rect 351276 529864 351328 529916
rect 338856 529796 338908 529848
rect 357440 529796 357492 529848
rect 322480 529660 322532 529712
rect 322848 529660 322900 529712
rect 401600 529116 401652 529168
rect 403808 529116 403860 529168
rect 401784 528640 401836 528692
rect 405096 528640 405148 528692
rect 254584 528572 254636 528624
rect 273996 528572 274048 528624
rect 452660 528572 452712 528624
rect 477592 528572 477644 528624
rect 322112 528504 322164 528556
rect 355232 528504 355284 528556
rect 401600 528436 401652 528488
rect 404452 528436 404504 528488
rect 322572 527144 322624 527196
rect 322756 527144 322808 527196
rect 418804 527144 418856 527196
rect 477592 527144 477644 527196
rect 322204 527076 322256 527128
rect 357440 527076 357492 527128
rect 412640 527076 412692 527128
rect 477684 527076 477736 527128
rect 322480 527008 322532 527060
rect 354404 527008 354456 527060
rect 355324 527008 355376 527060
rect 357532 527008 357584 527060
rect 322572 526940 322624 526992
rect 326344 526940 326396 526992
rect 401600 526396 401652 526448
rect 403256 526396 403308 526448
rect 358268 525784 358320 525836
rect 359464 525784 359516 525836
rect 400404 525784 400456 525836
rect 432604 525784 432656 525836
rect 460204 525784 460256 525836
rect 477592 525784 477644 525836
rect 522948 525784 523000 525836
rect 536104 525784 536156 525836
rect 401600 525716 401652 525768
rect 404636 525716 404688 525768
rect 527824 525716 527876 525768
rect 579804 525716 579856 525768
rect 401600 525240 401652 525292
rect 404360 525240 404412 525292
rect 322848 525036 322900 525088
rect 348516 525036 348568 525088
rect 422944 524424 422996 524476
rect 478144 524424 478196 524476
rect 334624 524356 334676 524408
rect 357440 524356 357492 524408
rect 401600 524356 401652 524408
rect 404820 524356 404872 524408
rect 322664 523676 322716 523728
rect 355232 523676 355284 523728
rect 254308 522996 254360 523048
rect 274088 522996 274140 523048
rect 522948 522996 523000 523048
rect 534724 522996 534776 523048
rect 322572 522928 322624 522980
rect 348424 522928 348476 522980
rect 322480 522248 322532 522300
rect 352472 522248 352524 522300
rect 322112 521908 322164 521960
rect 322664 521908 322716 521960
rect 401600 521636 401652 521688
rect 423772 521636 423824 521688
rect 322480 521568 322532 521620
rect 353208 521568 353260 521620
rect 401600 521024 401652 521076
rect 403440 521024 403492 521076
rect 322204 520888 322256 520940
rect 351276 520888 351328 520940
rect 322204 520752 322256 520804
rect 322388 520752 322440 520804
rect 522948 520616 523000 520668
rect 530584 520616 530636 520668
rect 322020 520276 322072 520328
rect 347044 520276 347096 520328
rect 321652 520208 321704 520260
rect 353024 520208 353076 520260
rect 357440 520208 357492 520260
rect 347688 520140 347740 520192
rect 354220 520140 354272 520192
rect 401600 520140 401652 520192
rect 405280 520140 405332 520192
rect 322204 519256 322256 519308
rect 325056 519256 325108 519308
rect 414020 518916 414072 518968
rect 477592 518916 477644 518968
rect 350080 518848 350132 518900
rect 357440 518848 357492 518900
rect 321744 518032 321796 518084
rect 324228 518032 324280 518084
rect 254584 517760 254636 517812
rect 258724 517760 258776 517812
rect 324320 517624 324372 517676
rect 325516 517624 325568 517676
rect 350724 517624 350776 517676
rect 322296 517556 322348 517608
rect 350632 517556 350684 517608
rect 355876 517556 355928 517608
rect 468484 517556 468536 517608
rect 477592 517556 477644 517608
rect 329196 517488 329248 517540
rect 357532 517488 357584 517540
rect 450544 517488 450596 517540
rect 477684 517488 477736 517540
rect 322848 517420 322900 517472
rect 324320 517420 324372 517472
rect 340144 517420 340196 517472
rect 357440 517420 357492 517472
rect 427084 517420 427136 517472
rect 477592 517420 477644 517472
rect 401600 516128 401652 516180
rect 405740 516128 405792 516180
rect 322296 516060 322348 516112
rect 342260 516060 342312 516112
rect 401692 516060 401744 516112
rect 404728 516060 404780 516112
rect 322848 515380 322900 515432
rect 324228 515380 324280 515432
rect 331956 515380 332008 515432
rect 342260 515380 342312 515432
rect 343548 515380 343600 515432
rect 355416 515380 355468 515432
rect 457444 514836 457496 514888
rect 477592 514836 477644 514888
rect 400864 514768 400916 514820
rect 477684 514768 477736 514820
rect 342904 514700 342956 514752
rect 357440 514700 357492 514752
rect 358636 514292 358688 514344
rect 359832 514292 359884 514344
rect 322756 514020 322808 514072
rect 322940 514020 322992 514072
rect 329104 514020 329156 514072
rect 322296 513408 322348 513460
rect 355324 513408 355376 513460
rect 413284 513340 413336 513392
rect 477592 513340 477644 513392
rect 331864 513272 331916 513324
rect 357440 513272 357492 513324
rect 522856 513204 522908 513256
rect 526444 513204 526496 513256
rect 402428 513068 402480 513120
rect 405372 513068 405424 513120
rect 322204 512592 322256 512644
rect 331220 512592 331272 512644
rect 476856 512048 476908 512100
rect 478144 512048 478196 512100
rect 436744 511980 436796 512032
rect 477684 511980 477736 512032
rect 322204 511912 322256 511964
rect 355784 511912 355836 511964
rect 358084 511912 358136 511964
rect 359464 511912 359516 511964
rect 432604 511912 432656 511964
rect 477592 511912 477644 511964
rect 320088 511844 320140 511896
rect 345848 511844 345900 511896
rect 347228 511844 347280 511896
rect 357440 511844 357492 511896
rect 321560 511232 321612 511284
rect 333888 511232 333940 511284
rect 357256 511232 357308 511284
rect 522948 510688 523000 510740
rect 538864 510688 538916 510740
rect 254400 510620 254452 510672
rect 271236 510620 271288 510672
rect 319076 510620 319128 510672
rect 320088 510620 320140 510672
rect 402888 510620 402940 510672
rect 451280 510620 451332 510672
rect 526444 510620 526496 510672
rect 580172 510620 580224 510672
rect 320364 510552 320416 510604
rect 341616 510552 341668 510604
rect 342996 510552 343048 510604
rect 357440 510552 357492 510604
rect 476948 510484 477000 510536
rect 478144 510484 478196 510536
rect 324228 509872 324280 509924
rect 350080 509872 350132 509924
rect 427728 509872 427780 509924
rect 468668 509872 468720 509924
rect 402888 509260 402940 509312
rect 427728 509260 427780 509312
rect 468576 509260 468628 509312
rect 477592 509260 477644 509312
rect 322296 509192 322348 509244
rect 355600 509192 355652 509244
rect 327724 509124 327776 509176
rect 357992 509124 358044 509176
rect 345664 509056 345716 509108
rect 357440 509056 357492 509108
rect 50804 508716 50856 508768
rect 51264 508716 51316 508768
rect 321652 508580 321704 508632
rect 322296 508580 322348 508632
rect 318892 508240 318944 508292
rect 319352 508240 319404 508292
rect 320272 508104 320324 508156
rect 320640 508104 320692 508156
rect 327816 508104 327868 508156
rect 319352 507832 319404 507884
rect 356612 507832 356664 507884
rect 445760 507832 445812 507884
rect 478144 507832 478196 507884
rect 320272 507764 320324 507816
rect 320548 507764 320600 507816
rect 355692 507764 355744 507816
rect 336004 507696 336056 507748
rect 357440 507696 357492 507748
rect 318892 506472 318944 506524
rect 319352 506472 319404 506524
rect 431960 506472 432012 506524
rect 477500 506472 477552 506524
rect 522948 506472 523000 506524
rect 527824 506472 527876 506524
rect 320272 506404 320324 506456
rect 351184 506404 351236 506456
rect 353116 506404 353168 506456
rect 357440 506404 357492 506456
rect 401600 506404 401652 506456
rect 403348 506404 403400 506456
rect 318984 506336 319036 506388
rect 320088 506336 320140 506388
rect 329748 506336 329800 506388
rect 350172 506336 350224 506388
rect 357624 506336 357676 506388
rect 329748 505724 329800 505776
rect 359280 505724 359332 505776
rect 322572 505248 322624 505300
rect 322756 505248 322808 505300
rect 254308 505112 254360 505164
rect 269948 505112 270000 505164
rect 322480 505044 322532 505096
rect 329196 505044 329248 505096
rect 341524 505044 341576 505096
rect 357440 505044 357492 505096
rect 357624 504364 357676 504416
rect 357900 504364 357952 504416
rect 349068 504160 349120 504212
rect 349988 504160 350040 504212
rect 320272 503820 320324 503872
rect 320548 503820 320600 503872
rect 321560 503684 321612 503736
rect 349068 503684 349120 503736
rect 322480 503616 322532 503668
rect 347136 503616 347188 503668
rect 401600 503616 401652 503668
rect 407120 503616 407172 503668
rect 322664 502936 322716 502988
rect 359372 502936 359424 502988
rect 462964 502324 463016 502376
rect 477500 502324 477552 502376
rect 337384 502256 337436 502308
rect 357440 502256 357492 502308
rect 434720 500964 434772 501016
rect 477500 500964 477552 501016
rect 322572 500896 322624 500948
rect 399576 500896 399628 500948
rect 478788 500896 478840 500948
rect 519728 500896 519780 500948
rect 347044 500828 347096 500880
rect 401968 500828 402020 500880
rect 359280 500760 359332 500812
rect 359924 500760 359976 500812
rect 295248 500352 295300 500404
rect 322940 500352 322992 500404
rect 322480 500284 322532 500336
rect 359740 500284 359792 500336
rect 296628 500216 296680 500268
rect 321744 500216 321796 500268
rect 322756 500216 322808 500268
rect 462320 500216 462372 500268
rect 477408 500216 477460 500268
rect 360476 499944 360528 499996
rect 359740 499876 359792 499928
rect 362960 499876 363012 499928
rect 363880 499876 363932 499928
rect 254584 499536 254636 499588
rect 262864 499536 262916 499588
rect 401600 499536 401652 499588
rect 433340 499536 433392 499588
rect 454684 499536 454736 499588
rect 477500 499536 477552 499588
rect 352932 499468 352984 499520
rect 379336 499468 379388 499520
rect 394148 499468 394200 499520
rect 403716 499468 403768 499520
rect 472716 499468 472768 499520
rect 485780 499468 485832 499520
rect 358912 499400 358964 499452
rect 478420 499400 478472 499452
rect 481364 499400 481416 499452
rect 520832 499400 520884 499452
rect 323676 499332 323728 499384
rect 369676 499332 369728 499384
rect 373540 499332 373592 499384
rect 472808 499332 472860 499384
rect 477684 499332 477736 499384
rect 492220 499332 492272 499384
rect 493600 499332 493652 499384
rect 523684 499332 523736 499384
rect 323584 499264 323636 499316
rect 397368 499264 397420 499316
rect 406476 499264 406528 499316
rect 505744 499264 505796 499316
rect 352840 499196 352892 499248
rect 399484 499196 399536 499248
rect 409236 499196 409288 499248
rect 494796 499196 494848 499248
rect 357164 499128 357216 499180
rect 402336 499128 402388 499180
rect 355416 499060 355468 499112
rect 398012 499060 398064 499112
rect 357256 498992 357308 499044
rect 389640 498992 389692 499044
rect 518256 498992 518308 499044
rect 522396 498992 522448 499044
rect 359924 498924 359976 498976
rect 381912 498924 381964 498976
rect 518164 498924 518216 498976
rect 522488 498924 522540 498976
rect 357348 498856 357400 498908
rect 367100 498856 367152 498908
rect 516784 498856 516836 498908
rect 522304 498856 522356 498908
rect 278780 498788 278832 498840
rect 320640 498788 320692 498840
rect 325056 498788 325108 498840
rect 353484 498788 353536 498840
rect 367744 498788 367796 498840
rect 506480 498788 506532 498840
rect 519820 498788 519872 498840
rect 320916 498720 320968 498772
rect 370320 498720 370372 498772
rect 375472 498720 375524 498772
rect 526444 498720 526496 498772
rect 354220 498176 354272 498228
rect 355416 498176 355468 498228
rect 355600 498176 355652 498228
rect 357072 498108 357124 498160
rect 361948 498108 362000 498160
rect 399300 498108 399352 498160
rect 403900 498108 403952 498160
rect 479524 498108 479576 498160
rect 483848 498108 483900 498160
rect 355416 498040 355468 498092
rect 361304 498040 361356 498092
rect 396724 498040 396776 498092
rect 403164 498040 403216 498092
rect 475568 498040 475620 498092
rect 512184 498040 512236 498092
rect 355968 497972 356020 498024
rect 364524 497972 364576 498024
rect 477040 497972 477092 498024
rect 489644 497972 489696 498024
rect 498844 497972 498896 498024
rect 499304 497972 499356 498024
rect 513472 497972 513524 498024
rect 296536 497904 296588 497956
rect 305552 497904 305604 497956
rect 355508 497904 355560 497956
rect 383844 497904 383896 497956
rect 388352 497904 388404 497956
rect 405188 497904 405240 497956
rect 477408 497904 477460 497956
rect 516048 497904 516100 497956
rect 298744 497836 298796 497888
rect 312176 497836 312228 497888
rect 352564 497836 352616 497888
rect 379980 497836 380032 497888
rect 291936 497768 291988 497820
rect 315120 497768 315172 497820
rect 352472 497768 352524 497820
rect 376116 497768 376168 497820
rect 376392 497768 376444 497820
rect 393504 497768 393556 497820
rect 286048 497700 286100 497752
rect 292028 497700 292080 497752
rect 293224 497700 293276 497752
rect 316040 497700 316092 497752
rect 354128 497700 354180 497752
rect 378048 497700 378100 497752
rect 258816 497632 258868 497684
rect 301872 497632 301924 497684
rect 355324 497632 355376 497684
rect 371608 497632 371660 497684
rect 459560 497632 459612 497684
rect 486424 497632 486476 497684
rect 510344 497632 510396 497684
rect 526444 497632 526496 497684
rect 267096 497564 267148 497616
rect 316592 497564 316644 497616
rect 349068 497564 349120 497616
rect 401692 497564 401744 497616
rect 456800 497564 456852 497616
rect 489000 497564 489052 497616
rect 489184 497564 489236 497616
rect 512828 497564 512880 497616
rect 256148 497496 256200 497548
rect 314660 497496 314712 497548
rect 352748 497496 352800 497548
rect 366456 497496 366508 497548
rect 398840 497496 398892 497548
rect 480628 497496 480680 497548
rect 491944 497496 491996 497548
rect 517336 497496 517388 497548
rect 257620 497428 257672 497480
rect 317420 497428 317472 497480
rect 350080 497428 350132 497480
rect 402060 497428 402112 497480
rect 409880 497428 409932 497480
rect 514760 497428 514812 497480
rect 349896 497360 349948 497412
rect 394792 497360 394844 497412
rect 352656 497292 352708 497344
rect 372252 497292 372304 497344
rect 349804 497224 349856 497276
rect 363236 497224 363288 497276
rect 486424 496816 486476 496868
rect 490932 496816 490984 496868
rect 493324 496816 493376 496868
rect 497372 496816 497424 496868
rect 479064 496748 479116 496800
rect 481640 496748 481692 496800
rect 294144 496340 294196 496392
rect 295984 496340 296036 496392
rect 357532 496340 357584 496392
rect 362224 496340 362276 496392
rect 488448 496340 488500 496392
rect 490564 496340 490616 496392
rect 501328 496204 501380 496256
rect 516876 496204 516928 496256
rect 297272 496136 297324 496188
rect 311900 496136 311952 496188
rect 358176 496136 358228 496188
rect 408500 496136 408552 496188
rect 498200 496136 498252 496188
rect 520096 496136 520148 496188
rect 285680 496068 285732 496120
rect 320364 496068 320416 496120
rect 374000 496068 374052 496120
rect 479708 496068 479760 496120
rect 491300 496068 491352 496120
rect 520924 496068 520976 496120
rect 299388 494980 299440 495032
rect 302332 494980 302384 495032
rect 484400 494776 484452 494828
rect 520372 494776 520424 494828
rect 284300 494708 284352 494760
rect 284944 494708 284996 494760
rect 287060 494708 287112 494760
rect 287888 494708 287940 494760
rect 289820 494708 289872 494760
rect 290832 494708 290884 494760
rect 292580 494708 292632 494760
rect 319076 494708 319128 494760
rect 358360 494708 358412 494760
rect 376024 494708 376076 494760
rect 478512 494708 478564 494760
rect 563060 494708 563112 494760
rect 299480 494640 299532 494692
rect 300400 494640 300452 494692
rect 307760 494096 307812 494148
rect 308496 494096 308548 494148
rect 254584 494028 254636 494080
rect 261576 494028 261628 494080
rect 478972 493484 479024 493536
rect 488540 493484 488592 493536
rect 378692 493416 378744 493468
rect 455420 493416 455472 493468
rect 483296 493416 483348 493468
rect 552020 493416 552072 493468
rect 441620 493348 441672 493400
rect 522212 493348 522264 493400
rect 264980 493280 265032 493332
rect 320456 493280 320508 493332
rect 396080 493280 396132 493332
rect 522028 493280 522080 493332
rect 500224 493008 500276 493060
rect 505100 493008 505152 493060
rect 479248 492056 479300 492108
rect 516140 492056 516192 492108
rect 478604 491988 478656 492040
rect 558184 491988 558236 492040
rect 297364 491920 297416 491972
rect 351920 491920 351972 491972
rect 353300 491920 353352 491972
rect 519636 491920 519688 491972
rect 288440 491512 288492 491564
rect 289360 491512 289412 491564
rect 407120 490560 407172 490612
rect 520004 490560 520056 490612
rect 254584 488520 254636 488572
rect 279516 488520 279568 488572
rect 49608 487840 49660 487892
rect 50344 487840 50396 487892
rect 307852 487840 307904 487892
rect 349712 487840 349764 487892
rect 478696 487840 478748 487892
rect 582380 487840 582432 487892
rect 267740 487772 267792 487824
rect 318984 487772 319036 487824
rect 355508 487772 355560 487824
rect 494152 487772 494204 487824
rect 276020 486412 276072 486464
rect 320272 486412 320324 486464
rect 479340 486412 479392 486464
rect 534080 486412 534132 486464
rect 525156 485732 525208 485784
rect 580172 485732 580224 485784
rect 479156 483624 479208 483676
rect 569960 483624 570012 483676
rect 289912 482264 289964 482316
rect 332600 482264 332652 482316
rect 254584 481652 254636 481704
rect 268476 481652 268528 481704
rect 49424 481584 49476 481636
rect 50436 481584 50488 481636
rect 364340 480904 364392 480956
rect 460204 480904 460256 480956
rect 389180 479476 389232 479528
rect 515404 479476 515456 479528
rect 371240 478116 371292 478168
rect 503904 478116 503956 478168
rect 254216 476076 254268 476128
rect 265716 476076 265768 476128
rect 363604 475328 363656 475380
rect 481916 475328 481968 475380
rect 46388 473288 46440 473340
rect 48964 473288 49016 473340
rect 338764 471928 338816 471980
rect 580172 471928 580224 471980
rect 254584 470568 254636 470620
rect 264336 470568 264388 470620
rect 45468 467780 45520 467832
rect 48780 467780 48832 467832
rect 49056 467780 49108 467832
rect 254584 465060 254636 465112
rect 271328 465060 271380 465112
rect 46480 462272 46532 462324
rect 50804 462272 50856 462324
rect 254584 458192 254636 458244
rect 278228 458192 278280 458244
rect 359832 458124 359884 458176
rect 580172 458124 580224 458176
rect 46572 456356 46624 456408
rect 49792 456356 49844 456408
rect 299572 453976 299624 454028
rect 300952 453976 301004 454028
rect 254308 452616 254360 452668
rect 289084 452616 289136 452668
rect 254676 447108 254728 447160
rect 275468 447108 275520 447160
rect 46664 445680 46716 445732
rect 48320 445680 48372 445732
rect 254400 441736 254452 441788
rect 257528 441736 257580 441788
rect 46756 438812 46808 438864
rect 48320 438812 48372 438864
rect 254400 434732 254452 434784
rect 291844 434732 291896 434784
rect 46848 433236 46900 433288
rect 49148 433236 49200 433288
rect 477868 431876 477920 431928
rect 579804 431876 579856 431928
rect 254584 429156 254636 429208
rect 350908 429156 350960 429208
rect 254584 423648 254636 423700
rect 323584 423648 323636 423700
rect 324964 419432 325016 419484
rect 580172 419432 580224 419484
rect 254584 418140 254636 418192
rect 282184 418140 282236 418192
rect 254584 411272 254636 411324
rect 349988 411272 350040 411324
rect 3148 409844 3200 409896
rect 50528 409844 50580 409896
rect 376024 405628 376076 405680
rect 580172 405628 580224 405680
rect 254032 400188 254084 400240
rect 350816 400188 350868 400240
rect 46848 397468 46900 397520
rect 49424 397468 49476 397520
rect 254676 394748 254728 394800
rect 260288 394748 260340 394800
rect 46756 391960 46808 392012
rect 48320 391960 48372 392012
rect 254676 389172 254728 389224
rect 317420 389172 317472 389224
rect 46664 385024 46716 385076
rect 48320 385024 48372 385076
rect 254400 382236 254452 382288
rect 289176 382236 289228 382288
rect 46572 379516 46624 379568
rect 49424 379516 49476 379568
rect 544384 379448 544436 379500
rect 580172 379448 580224 379500
rect 254124 376728 254176 376780
rect 351092 376728 351144 376780
rect 254676 371220 254728 371272
rect 301504 371220 301556 371272
rect 281540 369112 281592 369164
rect 283564 369112 283616 369164
rect 254676 365712 254728 365764
rect 282276 365712 282328 365764
rect 320824 365644 320876 365696
rect 580172 365644 580224 365696
rect 253940 358844 253992 358896
rect 256240 358844 256292 358896
rect 3148 357416 3200 357468
rect 50620 357416 50672 357468
rect 288532 353948 288584 354000
rect 352196 353948 352248 354000
rect 498752 353948 498804 354000
rect 540980 353948 541032 354000
rect 254216 353268 254268 353320
rect 289268 353268 289320 353320
rect 362224 353200 362276 353252
rect 580172 353200 580224 353252
rect 385040 352520 385092 352572
rect 521936 352520 521988 352572
rect 297640 351228 297692 351280
rect 313372 351228 313424 351280
rect 298008 351160 298060 351212
rect 320180 351160 320232 351212
rect 287152 349800 287204 349852
rect 350080 349800 350132 349852
rect 254492 347760 254544 347812
rect 346492 347760 346544 347812
rect 299664 345652 299716 345704
rect 314660 345652 314712 345704
rect 3332 345040 3384 345092
rect 50252 345040 50304 345092
rect 284392 344292 284444 344344
rect 352012 344292 352064 344344
rect 254584 342864 254636 342916
rect 351368 342864 351420 342916
rect 254584 342252 254636 342304
rect 287704 342252 287756 342304
rect 296996 341572 297048 341624
rect 311992 341572 312044 341624
rect 289820 341504 289872 341556
rect 349804 341504 349856 341556
rect 271880 340212 271932 340264
rect 318892 340212 318944 340264
rect 285772 340144 285824 340196
rect 352288 340144 352340 340196
rect 282920 338784 282972 338836
rect 318800 338784 318852 338836
rect 310612 338716 310664 338768
rect 350264 338716 350316 338768
rect 289820 337424 289872 337476
rect 322296 337424 322348 337476
rect 288440 337356 288492 337408
rect 352104 337356 352156 337408
rect 299480 335996 299532 336048
rect 319352 335996 319404 336048
rect 254400 335316 254452 335368
rect 332232 335316 332284 335368
rect 310520 334704 310572 334756
rect 352564 334704 352616 334756
rect 291292 334636 291344 334688
rect 351276 334636 351328 334688
rect 260840 334568 260892 334620
rect 321560 334568 321612 334620
rect 298652 333344 298704 333396
rect 307760 333344 307812 333396
rect 306472 333276 306524 333328
rect 352472 333276 352524 333328
rect 283104 333208 283156 333260
rect 350172 333208 350224 333260
rect 301504 332936 301556 332988
rect 306472 332936 306524 332988
rect 297916 332596 297968 332648
rect 298100 332596 298152 332648
rect 299756 332528 299808 332580
rect 306380 332528 306432 332580
rect 323584 332324 323636 332376
rect 325148 332324 325200 332376
rect 298836 332256 298888 332308
rect 347688 332256 347740 332308
rect 294604 332188 294656 332240
rect 310336 332188 310388 332240
rect 296260 332052 296312 332104
rect 309232 332052 309284 332104
rect 303804 331984 303856 332036
rect 320640 331984 320692 332036
rect 294972 331916 295024 331968
rect 305092 331916 305144 331968
rect 309140 331916 309192 331968
rect 353760 331916 353812 331968
rect 295064 331848 295116 331900
rect 302424 331848 302476 331900
rect 303620 331848 303672 331900
rect 353852 331848 353904 331900
rect 285036 331780 285088 331832
rect 321928 331780 321980 331832
rect 296352 331712 296404 331764
rect 309048 331712 309100 331764
rect 253296 331644 253348 331696
rect 341892 331644 341944 331696
rect 294880 331576 294932 331628
rect 313556 331576 313608 331628
rect 296444 331508 296496 331560
rect 330944 331508 330996 331560
rect 339316 331508 339368 331560
rect 354128 331508 354180 331560
rect 287796 331440 287848 331492
rect 323216 331440 323268 331492
rect 336096 331440 336148 331492
rect 352656 331440 352708 331492
rect 298560 331372 298612 331424
rect 307760 331372 307812 331424
rect 327724 331372 327776 331424
rect 352748 331372 352800 331424
rect 253204 331304 253256 331356
rect 300676 331304 300728 331356
rect 338028 331304 338080 331356
rect 353668 331304 353720 331356
rect 295156 331236 295208 331288
rect 301964 331236 302016 331288
rect 345112 331236 345164 331288
rect 349896 331236 349948 331288
rect 299020 330148 299072 330200
rect 326436 330148 326488 330200
rect 299112 330080 299164 330132
rect 329012 330080 329064 330132
rect 299204 330012 299256 330064
rect 334532 330012 334584 330064
rect 298928 329944 298980 329996
rect 340236 329944 340288 329996
rect 254216 329876 254268 329928
rect 284944 329876 284996 329928
rect 299296 329876 299348 329928
rect 343640 329876 343692 329928
rect 254676 329808 254728 329860
rect 351460 329808 351512 329860
rect 254492 325592 254544 325644
rect 285036 325592 285088 325644
rect 490564 325592 490616 325644
rect 580172 325592 580224 325644
rect 283564 324232 283616 324284
rect 297824 324232 297876 324284
rect 254308 320084 254360 320136
rect 287796 320084 287848 320136
rect 282276 318724 282328 318776
rect 297732 318724 297784 318776
rect 349804 318724 349856 318776
rect 349988 318656 350040 318708
rect 284944 317364 284996 317416
rect 297732 317364 297784 317416
rect 292764 313216 292816 313268
rect 297916 313216 297968 313268
rect 356980 313216 357032 313268
rect 580172 313216 580224 313268
rect 349988 312128 350040 312180
rect 349804 312060 349856 312112
rect 297916 311040 297968 311092
rect 298744 311040 298796 311092
rect 351184 310564 351236 310616
rect 351920 310564 351972 310616
rect 350264 309068 350316 309120
rect 351920 309068 351972 309120
rect 260288 307708 260340 307760
rect 297272 307708 297324 307760
rect 254216 306348 254268 306400
rect 293316 306348 293368 306400
rect 256240 306280 256292 306332
rect 298008 306280 298060 306332
rect 293960 303560 294012 303612
rect 298008 303560 298060 303612
rect 254676 300840 254728 300892
rect 294696 300840 294748 300892
rect 383200 299412 383252 299464
rect 580172 299412 580224 299464
rect 254676 295332 254728 295384
rect 284944 295332 284996 295384
rect 297824 295128 297876 295180
rect 299848 295128 299900 295180
rect 284300 292476 284352 292528
rect 298008 292476 298060 292528
rect 351368 291660 351420 291712
rect 353576 291660 353628 291712
rect 295432 289416 295484 289468
rect 298008 289416 298060 289468
rect 254400 288396 254452 288448
rect 296168 288396 296220 288448
rect 292028 288328 292080 288380
rect 298008 288328 298060 288380
rect 297824 287376 297876 287428
rect 297824 287036 297876 287088
rect 297824 285880 297876 285932
rect 297824 285676 297876 285728
rect 289176 285608 289228 285660
rect 297916 285608 297968 285660
rect 254308 282888 254360 282940
rect 264428 282888 264480 282940
rect 50620 282004 50672 282056
rect 298100 282004 298152 282056
rect 46664 281936 46716 281988
rect 279792 281936 279844 281988
rect 49148 281868 49200 281920
rect 278320 281868 278372 281920
rect 3516 281460 3568 281512
rect 519544 281460 519596 281512
rect 3424 281392 3476 281444
rect 485780 281392 485832 281444
rect 50528 281324 50580 281376
rect 521844 281324 521896 281376
rect 48964 281256 49016 281308
rect 53104 281256 53156 281308
rect 284944 281256 284996 281308
rect 352012 281256 352064 281308
rect 49056 281188 49108 281240
rect 54484 281188 54536 281240
rect 54576 281188 54628 281240
rect 279700 281188 279752 281240
rect 52092 281120 52144 281172
rect 280988 281120 281040 281172
rect 48688 281052 48740 281104
rect 280804 281052 280856 281104
rect 49240 280984 49292 281036
rect 276664 280984 276716 281036
rect 48044 280916 48096 280968
rect 54576 280916 54628 280968
rect 48780 280848 48832 280900
rect 272524 280916 272576 280968
rect 49332 280712 49384 280764
rect 287336 280712 287388 280764
rect 297732 280576 297784 280628
rect 300124 280576 300176 280628
rect 3608 280100 3660 280152
rect 468576 280100 468628 280152
rect 50252 280032 50304 280084
rect 507676 280032 507728 280084
rect 48228 279964 48280 280016
rect 279608 279964 279660 280016
rect 296168 279964 296220 280016
rect 351920 279964 351972 280016
rect 298560 279896 298612 279948
rect 303804 279896 303856 279948
rect 294880 279420 294932 279472
rect 310520 279420 310572 279472
rect 321652 279420 321704 279472
rect 354128 279420 354180 279472
rect 289268 279012 289320 279064
rect 315488 279012 315540 279064
rect 282276 278944 282328 278996
rect 321284 278944 321336 278996
rect 287704 278876 287756 278928
rect 330944 278876 330996 278928
rect 294696 278808 294748 278860
rect 342536 278808 342588 278860
rect 293316 278740 293368 278792
rect 349620 278740 349672 278792
rect 295984 278672 296036 278724
rect 301320 278672 301372 278724
rect 308404 278672 308456 278724
rect 313372 278672 313424 278724
rect 316776 278672 316828 278724
rect 323124 278672 323176 278724
rect 347044 278672 347096 278724
rect 353852 278672 353904 278724
rect 296536 278604 296588 278656
rect 305184 278604 305236 278656
rect 339960 278604 340012 278656
rect 353760 278604 353812 278656
rect 295340 278536 295392 278588
rect 335452 278536 335504 278588
rect 292672 278468 292724 278520
rect 319996 278468 320048 278520
rect 296260 278400 296312 278452
rect 322572 278400 322624 278452
rect 299756 278332 299808 278384
rect 318064 278332 318116 278384
rect 337384 278332 337436 278384
rect 341248 278332 341300 278384
rect 287060 278264 287112 278316
rect 303896 278264 303948 278316
rect 294972 278196 295024 278248
rect 338028 278196 338080 278248
rect 298744 278128 298796 278180
rect 303712 278128 303764 278180
rect 334164 278060 334216 278112
rect 338212 278060 338264 278112
rect 59452 277992 59504 278044
rect 297364 277992 297416 278044
rect 317420 277992 317472 278044
rect 343824 277992 343876 278044
rect 295064 277924 295116 277976
rect 345756 277924 345808 277976
rect 300032 277584 300084 277636
rect 305644 277584 305696 277636
rect 323860 277516 323912 277568
rect 326344 277516 326396 277568
rect 324320 277380 324372 277432
rect 327080 277380 327132 277432
rect 297456 276768 297508 276820
rect 309140 276768 309192 276820
rect 314752 276768 314804 276820
rect 351092 276768 351144 276820
rect 59268 276700 59320 276752
rect 352104 276700 352156 276752
rect 3424 276632 3476 276684
rect 519452 276632 519504 276684
rect 299664 276088 299716 276140
rect 305000 276088 305052 276140
rect 297640 276020 297692 276072
rect 298836 276020 298888 276072
rect 297180 275340 297232 275392
rect 311164 275340 311216 275392
rect 7564 275272 7616 275324
rect 501880 275272 501932 275324
rect 297548 273980 297600 274032
rect 335360 273980 335412 274032
rect 3700 273912 3752 273964
rect 520740 273912 520792 273964
rect 499948 273164 500000 273216
rect 580172 273164 580224 273216
rect 333980 272620 334032 272672
rect 349804 272620 349856 272672
rect 58900 272552 58952 272604
rect 352380 272552 352432 272604
rect 4804 272484 4856 272536
rect 496728 272484 496780 272536
rect 299572 271124 299624 271176
rect 318800 271124 318852 271176
rect 9680 268336 9732 268388
rect 478236 268336 478288 268388
rect 13820 266976 13872 267028
rect 457444 266976 457496 267028
rect 318892 260108 318944 260160
rect 351000 260108 351052 260160
rect 301504 258680 301556 258732
rect 350908 258680 350960 258732
rect 302332 257320 302384 257372
rect 384488 257320 384540 257372
rect 3148 255212 3200 255264
rect 436836 255212 436888 255264
rect 59084 253172 59136 253224
rect 347780 253172 347832 253224
rect 359648 245556 359700 245608
rect 580172 245556 580224 245608
rect 3516 241408 3568 241460
rect 423036 241408 423088 241460
rect 58992 236648 59044 236700
rect 352288 236648 352340 236700
rect 59636 235220 59688 235272
rect 311900 235220 311952 235272
rect 58808 233860 58860 233912
rect 310612 233860 310664 233912
rect 534724 233180 534776 233232
rect 579988 233180 580040 233232
rect 8944 231072 8996 231124
rect 487068 231072 487120 231124
rect 60004 229712 60056 229764
rect 507124 229712 507176 229764
rect 57336 228420 57388 228472
rect 256148 228420 256200 228472
rect 59544 228352 59596 228404
rect 324412 228352 324464 228404
rect 326068 228352 326120 228404
rect 349712 228352 349764 228404
rect 31024 226992 31076 227044
rect 478144 226992 478196 227044
rect 59176 225632 59228 225684
rect 283196 225632 283248 225684
rect 57796 225564 57848 225616
rect 296076 225564 296128 225616
rect 308864 225564 308916 225616
rect 332600 225564 332652 225616
rect 318800 224272 318852 224324
rect 319628 224272 319680 224324
rect 3792 224204 3844 224256
rect 454776 224204 454828 224256
rect 305644 223524 305696 223576
rect 307852 223524 307904 223576
rect 299940 223456 299992 223508
rect 306840 223456 306892 223508
rect 302240 223184 302292 223236
rect 314936 223184 314988 223236
rect 329104 223184 329156 223236
rect 309232 223116 309284 223168
rect 323032 223116 323084 223168
rect 328092 223116 328144 223168
rect 337200 223184 337252 223236
rect 350080 223184 350132 223236
rect 296352 223048 296404 223100
rect 299848 222980 299900 223032
rect 321008 222980 321060 223032
rect 326344 223048 326396 223100
rect 333152 223048 333204 223100
rect 331128 222980 331180 223032
rect 352656 223116 352708 223168
rect 334164 223048 334216 223100
rect 349896 223048 349948 223100
rect 353668 222980 353720 223032
rect 57520 222912 57572 222964
rect 253296 222912 253348 222964
rect 295156 222912 295208 222964
rect 330116 222912 330168 222964
rect 332140 222912 332192 222964
rect 352748 222912 352800 222964
rect 57060 222844 57112 222896
rect 267096 222844 267148 222896
rect 296444 222844 296496 222896
rect 311164 222844 311216 222896
rect 312912 222844 312964 222896
rect 316960 222844 317012 222896
rect 351184 222844 351236 222896
rect 311900 222776 311952 222828
rect 222844 222232 222896 222284
rect 301504 222232 301556 222284
rect 224408 222164 224460 222216
rect 339224 222164 339276 222216
rect 299480 222096 299532 222148
rect 300768 222096 300820 222148
rect 297364 221552 297416 221604
rect 336924 221552 336976 221604
rect 57244 221484 57296 221536
rect 254584 221484 254636 221536
rect 297456 221484 297508 221536
rect 337384 221484 337436 221536
rect 58716 221416 58768 221468
rect 352840 221416 352892 221468
rect 226064 220804 226116 220856
rect 300768 220804 300820 220856
rect 578884 220804 578936 220856
rect 299388 220260 299440 220312
rect 306380 220260 306432 220312
rect 57152 220192 57204 220244
rect 291936 220192 291988 220244
rect 298836 220192 298888 220244
rect 313280 220192 313332 220244
rect 60556 220124 60608 220176
rect 293224 220124 293276 220176
rect 298744 220124 298796 220176
rect 328460 220124 328512 220176
rect 3608 220056 3660 220108
rect 520648 220056 520700 220108
rect 57888 218832 57940 218884
rect 253204 218832 253256 218884
rect 57428 218764 57480 218816
rect 258816 218764 258868 218816
rect 57612 218696 57664 218748
rect 294604 218696 294656 218748
rect 222936 216656 222988 216708
rect 297916 216656 297968 216708
rect 247684 215296 247736 215348
rect 297916 215296 297968 215348
rect 57244 214548 57296 214600
rect 57704 214548 57756 214600
rect 246304 213936 246356 213988
rect 297916 213936 297968 213988
rect 222292 212984 222344 213036
rect 226064 212984 226116 213036
rect 242164 212508 242216 212560
rect 297916 212508 297968 212560
rect 239404 211148 239456 211200
rect 297916 211148 297968 211200
rect 238024 209788 238076 209840
rect 297916 209788 297968 209840
rect 235264 208360 235316 208412
rect 296812 208360 296864 208412
rect 287704 207000 287756 207052
rect 297916 207000 297968 207052
rect 409144 206932 409196 206984
rect 579804 206932 579856 206984
rect 284944 205640 284996 205692
rect 296812 205640 296864 205692
rect 223212 205572 223264 205624
rect 229744 205572 229796 205624
rect 282184 202852 282236 202904
rect 297916 202852 297968 202904
rect 253204 201492 253256 201544
rect 297916 201492 297968 201544
rect 51080 201424 51132 201476
rect 57336 201424 57388 201476
rect 228364 200132 228416 200184
rect 297916 200132 297968 200184
rect 225604 198704 225656 198756
rect 297916 198704 297968 198756
rect 224316 197344 224368 197396
rect 297916 197344 297968 197396
rect 50436 197276 50488 197328
rect 57336 197276 57388 197328
rect 224224 195984 224276 196036
rect 297916 195984 297968 196036
rect 223488 194556 223540 194608
rect 233976 194556 234028 194608
rect 250444 194556 250496 194608
rect 297916 194556 297968 194608
rect 243544 193196 243596 193248
rect 297916 193196 297968 193248
rect 229744 193128 229796 193180
rect 297732 193128 297784 193180
rect 516876 193128 516928 193180
rect 580172 193128 580224 193180
rect 50988 192924 51040 192976
rect 57336 192924 57388 192976
rect 223488 191836 223540 191888
rect 232504 191836 232556 191888
rect 233884 190476 233936 190528
rect 297916 190476 297968 190528
rect 222844 190408 222896 190460
rect 297732 190408 297784 190460
rect 223488 189048 223540 189100
rect 230388 189048 230440 189100
rect 50896 188980 50948 189032
rect 57336 188980 57388 189032
rect 223028 188980 223080 189032
rect 297916 188980 297968 189032
rect 223488 186328 223540 186380
rect 295984 186328 296036 186380
rect 222936 186260 222988 186312
rect 296812 186260 296864 186312
rect 51172 184832 51224 184884
rect 56692 184832 56744 184884
rect 233976 184832 234028 184884
rect 297916 184832 297968 184884
rect 222292 184152 222344 184204
rect 225696 184152 225748 184204
rect 232504 183472 232556 183524
rect 297916 183472 297968 183524
rect 230388 182112 230440 182164
rect 297916 182112 297968 182164
rect 51264 180752 51316 180804
rect 56692 180752 56744 180804
rect 225696 179324 225748 179376
rect 297916 179324 297968 179376
rect 356888 179324 356940 179376
rect 580172 179324 580224 179376
rect 223488 177964 223540 178016
rect 297916 177964 297968 178016
rect 357624 177352 357676 177404
rect 473452 177352 473504 177404
rect 382280 177284 382332 177336
rect 521752 177284 521804 177336
rect 50344 176604 50396 176656
rect 57336 176604 57388 176656
rect 222660 176604 222712 176656
rect 297916 176604 297968 176656
rect 358544 175924 358596 175976
rect 426440 175924 426492 175976
rect 222660 175176 222712 175228
rect 297916 175176 297968 175228
rect 48872 173340 48924 173392
rect 57244 173340 57296 173392
rect 222384 173136 222436 173188
rect 297916 173136 297968 173188
rect 222476 171096 222528 171148
rect 297916 171096 297968 171148
rect 222936 169736 222988 169788
rect 296812 169736 296864 169788
rect 49516 169668 49568 169720
rect 57336 169668 57388 169720
rect 223488 167016 223540 167068
rect 297916 167016 297968 167068
rect 405096 166948 405148 167000
rect 580172 166948 580224 167000
rect 223028 165588 223080 165640
rect 297916 165588 297968 165640
rect 222936 164228 222988 164280
rect 297916 164228 297968 164280
rect 223488 162868 223540 162920
rect 297916 162868 297968 162920
rect 229100 161440 229152 161492
rect 297916 161440 297968 161492
rect 54576 161372 54628 161424
rect 57060 161372 57112 161424
rect 225788 158720 225840 158772
rect 297916 158720 297968 158772
rect 232596 157360 232648 157412
rect 297916 157360 297968 157412
rect 53104 157292 53156 157344
rect 57060 157292 57112 157344
rect 222660 157292 222712 157344
rect 229100 157292 229152 157344
rect 229836 155932 229888 155984
rect 297916 155932 297968 155984
rect 222936 154572 222988 154624
rect 297916 154572 297968 154624
rect 222844 153212 222896 153264
rect 297916 153212 297968 153264
rect 54484 153144 54536 153196
rect 57336 153144 57388 153196
rect 518624 153144 518676 153196
rect 580172 153144 580224 153196
rect 231124 151784 231176 151836
rect 296812 151784 296864 151836
rect 223212 151036 223264 151088
rect 295984 151036 296036 151088
rect 2780 150288 2832 150340
rect 4804 150288 4856 150340
rect 228456 149064 228508 149116
rect 297916 149064 297968 149116
rect 50804 148996 50856 149048
rect 57336 148996 57388 149048
rect 222568 147092 222620 147144
rect 225788 147092 225840 147144
rect 225696 146276 225748 146328
rect 297916 146276 297968 146328
rect 229744 144916 229796 144968
rect 297916 144916 297968 144968
rect 223488 144848 223540 144900
rect 232596 144848 232648 144900
rect 50712 144508 50764 144560
rect 57336 144508 57388 144560
rect 232504 143556 232556 143608
rect 297916 143556 297968 143608
rect 257344 142060 257396 142112
rect 297916 142060 297968 142112
rect 223488 141448 223540 141500
rect 229836 141448 229888 141500
rect 51356 140700 51408 140752
rect 57428 140700 57480 140752
rect 257436 140700 257488 140752
rect 297916 140700 297968 140752
rect 269856 139340 269908 139392
rect 297916 139340 297968 139392
rect 354036 139340 354088 139392
rect 580172 139340 580224 139392
rect 222660 137912 222712 137964
rect 231124 137912 231176 137964
rect 275376 137912 275428 137964
rect 297916 137912 297968 137964
rect 273996 136552 274048 136604
rect 297916 136552 297968 136604
rect 274088 135192 274140 135244
rect 297916 135192 297968 135244
rect 222844 133152 222896 133204
rect 296076 133152 296128 133204
rect 258724 132404 258776 132456
rect 296812 132404 296864 132456
rect 271236 131044 271288 131096
rect 297916 131044 297968 131096
rect 223028 130024 223080 130076
rect 228456 130024 228508 130076
rect 269948 129684 270000 129736
rect 296812 129684 296864 129736
rect 222292 128256 222344 128308
rect 225696 128256 225748 128308
rect 262864 128256 262916 128308
rect 297916 128256 297968 128308
rect 261576 126896 261628 126948
rect 297916 126896 297968 126948
rect 372896 126896 372948 126948
rect 580172 126896 580224 126948
rect 279516 125536 279568 125588
rect 297916 125536 297968 125588
rect 268476 124108 268528 124160
rect 297916 124108 297968 124160
rect 265716 122748 265768 122800
rect 297916 122748 297968 122800
rect 264336 121388 264388 121440
rect 297916 121388 297968 121440
rect 223488 120640 223540 120692
rect 229744 120640 229796 120692
rect 271328 120028 271380 120080
rect 297916 120028 297968 120080
rect 223488 118600 223540 118652
rect 232504 118600 232556 118652
rect 278228 118600 278280 118652
rect 297916 118600 297968 118652
rect 289084 117240 289136 117292
rect 297916 117240 297968 117292
rect 342352 117240 342404 117292
rect 363604 117240 363656 117292
rect 223488 115880 223540 115932
rect 295984 115880 296036 115932
rect 275468 114452 275520 114504
rect 296812 114452 296864 114504
rect 257528 113092 257580 113144
rect 297916 113092 297968 113144
rect 530584 113092 530636 113144
rect 579804 113092 579856 113144
rect 222200 112956 222252 113008
rect 224408 112956 224460 113008
rect 223488 110372 223540 110424
rect 247684 110372 247736 110424
rect 357716 109692 357768 109744
rect 580264 109692 580316 109744
rect 342352 108944 342404 108996
rect 440884 108944 440936 108996
rect 222660 107584 222712 107636
rect 246304 107584 246356 107636
rect 342352 106224 342404 106276
rect 518256 106224 518308 106276
rect 222844 104796 222896 104848
rect 242164 104796 242216 104848
rect 223488 102076 223540 102128
rect 239404 102076 239456 102128
rect 223028 99288 223080 99340
rect 238024 99288 238076 99340
rect 223120 96568 223172 96620
rect 235264 96568 235316 96620
rect 223488 93780 223540 93832
rect 287704 93780 287756 93832
rect 223488 91740 223540 91792
rect 284944 91740 284996 91792
rect 267004 90312 267056 90364
rect 297364 90312 297416 90364
rect 264244 88952 264296 89004
rect 296812 88952 296864 89004
rect 357808 88952 357860 89004
rect 415400 88952 415452 89004
rect 223212 88272 223264 88324
rect 282184 88272 282236 88324
rect 291844 88272 291896 88324
rect 298008 88272 298060 88324
rect 260196 86912 260248 86964
rect 297180 86912 297232 86964
rect 223212 85484 223264 85536
rect 253204 85484 253256 85536
rect 3424 85008 3476 85060
rect 8944 85008 8996 85060
rect 273904 84124 273956 84176
rect 297916 84124 297968 84176
rect 271144 82764 271196 82816
rect 297916 82764 297968 82816
rect 223488 81336 223540 81388
rect 228364 81336 228416 81388
rect 269764 79976 269816 80028
rect 298008 79976 298060 80028
rect 275284 78616 275336 78668
rect 297548 78616 297600 78668
rect 222476 78548 222528 78600
rect 225604 78548 225656 78600
rect 260104 77188 260156 77240
rect 297180 77188 297232 77240
rect 255964 75828 256016 75880
rect 298008 75828 298060 75880
rect 222200 75692 222252 75744
rect 224316 75692 224368 75744
rect 278044 74468 278096 74520
rect 298008 74468 298060 74520
rect 256056 73108 256108 73160
rect 296812 73108 296864 73160
rect 543004 73108 543056 73160
rect 580172 73108 580224 73160
rect 222200 73040 222252 73092
rect 224224 73040 224276 73092
rect 279424 71680 279476 71732
rect 297732 71680 297784 71732
rect 223488 70320 223540 70372
rect 250444 70320 250496 70372
rect 265624 70320 265676 70372
rect 298008 70320 298060 70372
rect 342996 69028 343048 69080
rect 489920 69028 489972 69080
rect 268384 68960 268436 69012
rect 297180 68960 297232 69012
rect 223488 67532 223540 67584
rect 243544 67532 243596 67584
rect 261484 67532 261536 67584
rect 297548 67532 297600 67584
rect 342996 66240 343048 66292
rect 418896 66240 418948 66292
rect 222844 64812 222896 64864
rect 233884 64812 233936 64864
rect 278136 64812 278188 64864
rect 297916 64812 297968 64864
rect 342996 63520 343048 63572
rect 483020 63520 483072 63572
rect 342444 62840 342496 62892
rect 342996 62840 343048 62892
rect 342352 62092 342404 62144
rect 480260 62092 480312 62144
rect 264428 62024 264480 62076
rect 298008 62024 298060 62076
rect 215300 61480 215352 61532
rect 342628 61480 342680 61532
rect 158720 61412 158772 61464
rect 342812 61412 342864 61464
rect 154580 61344 154632 61396
rect 342904 61344 342956 61396
rect 353944 60664 353996 60716
rect 580172 60664 580224 60716
rect 296628 60324 296680 60376
rect 303620 60324 303672 60376
rect 295248 60256 295300 60308
rect 310520 60256 310572 60308
rect 314660 60256 314712 60308
rect 355600 60256 355652 60308
rect 211160 60188 211212 60240
rect 342720 60188 342772 60240
rect 197360 60120 197412 60172
rect 341340 60120 341392 60172
rect 168380 60052 168432 60104
rect 341708 60052 341760 60104
rect 133880 59984 133932 60036
rect 340512 59984 340564 60036
rect 247040 58828 247092 58880
rect 340144 58828 340196 58880
rect 172520 58760 172572 58812
rect 341616 58760 341668 58812
rect 151820 58692 151872 58744
rect 343180 58692 343232 58744
rect 140780 58624 140832 58676
rect 342444 58624 342496 58676
rect 233240 57332 233292 57384
rect 342996 57332 343048 57384
rect 179420 57264 179472 57316
rect 341432 57264 341484 57316
rect 176660 57196 176712 57248
rect 341524 57196 341576 57248
rect 236000 55904 236052 55956
rect 340236 55904 340288 55956
rect 190460 55836 190512 55888
rect 340420 55836 340472 55888
rect 218060 54476 218112 54528
rect 342536 54476 342588 54528
rect 226340 53048 226392 53100
rect 341156 53048 341208 53100
rect 251180 51688 251232 51740
rect 341064 51688 341116 51740
rect 201500 47540 201552 47592
rect 498844 47540 498896 47592
rect 359556 46860 359608 46912
rect 580172 46860 580224 46912
rect 242900 46180 242952 46232
rect 343088 46180 343140 46232
rect 3424 45500 3476 45552
rect 355508 45500 355560 45552
rect 204260 44820 204312 44872
rect 340328 44820 340380 44872
rect 222200 42168 222252 42220
rect 340052 42168 340104 42220
rect 193220 42100 193272 42152
rect 341248 42100 341300 42152
rect 99380 42032 99432 42084
rect 520556 42032 520608 42084
rect 120080 40672 120132 40724
rect 509700 40672 509752 40724
rect 85580 35164 85632 35216
rect 486424 35164 486476 35216
rect 510896 33056 510948 33108
rect 580172 33056 580224 33108
rect 77300 32376 77352 32428
rect 436744 32376 436796 32428
rect 74540 31016 74592 31068
rect 493324 31016 493376 31068
rect 349160 28296 349212 28348
rect 476856 28296 476908 28348
rect 113180 28228 113232 28280
rect 454684 28228 454736 28280
rect 63500 26868 63552 26920
rect 472624 26868 472676 26920
rect 60740 25508 60792 25560
rect 475476 25508 475528 25560
rect 391940 24080 391992 24132
rect 468484 24080 468536 24132
rect 346400 22720 346452 22772
rect 413284 22720 413336 22772
rect 392216 21428 392268 21480
rect 412640 21428 412692 21480
rect 2780 21360 2832 21412
rect 422944 21360 422996 21412
rect 3424 20612 3476 20664
rect 450544 20612 450596 20664
rect 356796 20544 356848 20596
rect 580172 20544 580224 20596
rect 1400 18572 1452 18624
rect 476764 18572 476816 18624
rect 378140 17212 378192 17264
rect 462964 17212 463016 17264
rect 390928 15920 390980 15972
rect 440240 15920 440292 15972
rect 95792 15852 95844 15904
rect 400864 15852 400916 15904
rect 367744 14492 367796 14544
rect 418804 14492 418856 14544
rect 102140 14424 102192 14476
rect 519912 14424 519964 14476
rect 258264 13064 258316 13116
rect 494704 13064 494756 13116
rect 240140 10276 240192 10328
rect 340880 10276 340932 10328
rect 427728 9052 427780 9104
rect 494704 9052 494756 9104
rect 110512 8984 110564 9036
rect 521108 8984 521160 9036
rect 82084 8916 82136 8968
rect 521016 8916 521068 8968
rect 396172 8236 396224 8288
rect 402520 8236 402572 8288
rect 229836 7624 229888 7676
rect 342260 7624 342312 7676
rect 418896 7624 418948 7676
rect 487620 7624 487672 7676
rect 39580 7556 39632 7608
rect 522580 7556 522632 7608
rect 359464 6808 359516 6860
rect 580172 6808 580224 6860
rect 3424 6604 3476 6656
rect 7564 6604 7616 6656
rect 32404 6128 32456 6180
rect 491576 6128 491628 6180
rect 208584 4836 208636 4888
rect 340972 4836 341024 4888
rect 357532 4836 357584 4888
rect 517980 4836 518032 4888
rect 50160 4768 50212 4820
rect 508320 4768 508372 4820
rect 332692 4088 332744 4140
rect 350632 4088 350684 4140
rect 499396 4088 499448 4140
rect 500224 4088 500276 4140
rect 336280 4020 336332 4072
rect 355416 4020 355468 4072
rect 325608 3952 325660 4004
rect 350540 3952 350592 4004
rect 322112 3884 322164 3936
rect 350724 3884 350776 3936
rect 307944 3816 307996 3868
rect 355324 3816 355376 3868
rect 361120 3816 361172 3868
rect 405004 3816 405056 3868
rect 117596 3748 117648 3800
rect 406384 3748 406436 3800
rect 124680 3680 124732 3732
rect 475384 3680 475436 3732
rect 491300 3680 491352 3732
rect 491944 3680 491996 3732
rect 46664 3612 46716 3664
rect 403716 3612 403768 3664
rect 478144 3612 478196 3664
rect 518164 3612 518216 3664
rect 540244 3612 540296 3664
rect 582196 3612 582248 3664
rect 28908 3544 28960 3596
rect 410524 3544 410576 3596
rect 415400 3544 415452 3596
rect 416688 3544 416740 3596
rect 423680 3544 423732 3596
rect 424968 3544 425020 3596
rect 440240 3544 440292 3596
rect 441528 3544 441580 3596
rect 449808 3544 449860 3596
rect 516784 3544 516836 3596
rect 525064 3544 525116 3596
rect 531320 3544 531372 3596
rect 536104 3544 536156 3596
rect 573916 3544 573968 3596
rect 57244 3476 57296 3528
rect 60004 3476 60056 3528
rect 102140 3476 102192 3528
rect 103336 3476 103388 3528
rect 106924 3476 106976 3528
rect 491300 3476 491352 3528
rect 526444 3476 526496 3528
rect 527824 3476 527876 3528
rect 527916 3476 527968 3528
rect 538404 3476 538456 3528
rect 538864 3476 538916 3528
rect 19432 3408 19484 3460
rect 31024 3408 31076 3460
rect 35992 3408 36044 3460
rect 48964 3408 49016 3460
rect 89168 3408 89220 3460
rect 489184 3408 489236 3460
rect 504456 3408 504508 3460
rect 577412 3408 577464 3460
rect 578884 3476 578936 3528
rect 579804 3476 579856 3528
rect 581000 3408 581052 3460
rect 168380 3340 168432 3392
rect 169576 3340 169628 3392
rect 193220 3340 193272 3392
rect 194416 3340 194468 3392
rect 218060 3340 218112 3392
rect 219256 3340 219308 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 339868 3340 339920 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 473360 3340 473412 3392
rect 474188 3340 474240 3392
rect 558184 3340 558236 3392
rect 559748 3340 559800 3392
rect 353484 3272 353536 3324
rect 343364 3204 343416 3256
rect 353392 3204 353444 3256
<< metal2 >>
rect 6932 703582 7972 703610
rect 3238 671256 3294 671265
rect 3238 671191 3294 671200
rect 3252 667214 3280 671191
rect 3240 667208 3292 667214
rect 3240 667150 3292 667156
rect 6932 661706 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700330 24348 703520
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 40052 665854 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 665848 40092 665854
rect 40040 665790 40092 665796
rect 46572 663808 46624 663814
rect 46572 663750 46624 663756
rect 46480 662652 46532 662658
rect 46480 662594 46532 662600
rect 45468 662584 45520 662590
rect 45468 662526 45520 662532
rect 6920 661700 6972 661706
rect 6920 661642 6972 661648
rect 3516 661088 3568 661094
rect 3516 661030 3568 661036
rect 3424 659932 3476 659938
rect 3424 659874 3476 659880
rect 3332 659864 3384 659870
rect 3332 659806 3384 659812
rect 3344 658209 3372 659806
rect 3330 658200 3386 658209
rect 3330 658135 3386 658144
rect 3332 567180 3384 567186
rect 3332 567122 3384 567128
rect 3344 566953 3372 567122
rect 3330 566944 3386 566953
rect 3330 566879 3386 566888
rect 2964 554736 3016 554742
rect 2964 554678 3016 554684
rect 2976 553897 3004 554678
rect 2962 553888 3018 553897
rect 2962 553823 3018 553832
rect 3436 449585 3464 659874
rect 3528 462641 3556 661030
rect 3606 659968 3662 659977
rect 3606 659903 3662 659912
rect 3620 514865 3648 659903
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 45480 467838 45508 662526
rect 46388 662448 46440 662454
rect 46388 662390 46440 662396
rect 46400 473346 46428 662390
rect 46388 473340 46440 473346
rect 46388 473282 46440 473288
rect 45468 467832 45520 467838
rect 45468 467774 45520 467780
rect 3514 462632 3570 462641
rect 3514 462567 3570 462576
rect 46492 462330 46520 662594
rect 46480 462324 46532 462330
rect 46480 462266 46532 462272
rect 46584 456414 46612 663750
rect 47950 663232 48006 663241
rect 47950 663167 48006 663176
rect 52000 663196 52052 663202
rect 46664 663060 46716 663066
rect 46664 663002 46716 663008
rect 46572 456408 46624 456414
rect 46572 456350 46624 456356
rect 3422 449576 3478 449585
rect 3422 449511 3478 449520
rect 46676 445738 46704 663002
rect 46846 662960 46902 662969
rect 46846 662895 46902 662904
rect 46754 662824 46810 662833
rect 46754 662759 46810 662768
rect 46664 445732 46716 445738
rect 46664 445674 46716 445680
rect 46768 438870 46796 662759
rect 46756 438864 46808 438870
rect 46756 438806 46808 438812
rect 46860 433294 46888 662895
rect 47860 662856 47912 662862
rect 47860 662798 47912 662804
rect 47872 590646 47900 662798
rect 47860 590640 47912 590646
rect 47860 590582 47912 590588
rect 46848 433288 46900 433294
rect 46848 433230 46900 433236
rect 47964 427145 47992 663167
rect 52000 663138 52052 663144
rect 51908 663128 51960 663134
rect 51908 663070 51960 663076
rect 51172 662924 51224 662930
rect 51172 662866 51224 662872
rect 51080 662788 51132 662794
rect 51080 662730 51132 662736
rect 50988 662720 51040 662726
rect 50988 662662 51040 662668
rect 49974 661872 50030 661881
rect 49974 661807 50030 661816
rect 48872 661632 48924 661638
rect 48872 661574 48924 661580
rect 49330 661600 49386 661609
rect 48504 661564 48556 661570
rect 48504 661506 48556 661512
rect 48136 660204 48188 660210
rect 48136 660146 48188 660152
rect 48044 660136 48096 660142
rect 48044 660078 48096 660084
rect 47950 427136 48006 427145
rect 47950 427071 48006 427080
rect 48056 421297 48084 660078
rect 48042 421288 48098 421297
rect 48042 421223 48098 421232
rect 48148 415449 48176 660146
rect 48228 660068 48280 660074
rect 48228 660010 48280 660016
rect 48134 415440 48190 415449
rect 48134 415375 48190 415384
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 48240 409601 48268 660010
rect 48516 612785 48544 661506
rect 48594 660104 48650 660113
rect 48594 660039 48650 660048
rect 48608 620129 48636 660039
rect 48688 652792 48740 652798
rect 48688 652734 48740 652740
rect 48594 620120 48650 620129
rect 48594 620055 48650 620064
rect 48502 612776 48558 612785
rect 48502 612711 48558 612720
rect 48700 579193 48728 652734
rect 48884 631825 48912 661574
rect 49330 661535 49386 661544
rect 49054 661328 49110 661337
rect 49054 661263 49110 661272
rect 48962 661056 49018 661065
rect 48962 660991 49018 661000
rect 48870 631816 48926 631825
rect 48870 631751 48926 631760
rect 48872 618996 48924 619002
rect 48872 618938 48924 618944
rect 48780 612808 48832 612814
rect 48780 612750 48832 612756
rect 48686 579184 48742 579193
rect 48686 579119 48742 579128
rect 48792 555801 48820 612750
rect 48778 555792 48834 555801
rect 48778 555727 48834 555736
rect 48884 549953 48912 618938
rect 48976 596737 49004 660991
rect 48962 596728 49018 596737
rect 48962 596663 49018 596672
rect 49068 590889 49096 661263
rect 49238 660376 49294 660385
rect 49238 660311 49294 660320
rect 49148 641776 49200 641782
rect 49148 641718 49200 641724
rect 49054 590880 49110 590889
rect 49054 590815 49110 590824
rect 48964 590640 49016 590646
rect 48964 590582 49016 590588
rect 48870 549944 48926 549953
rect 48870 549879 48926 549888
rect 48976 499574 49004 590582
rect 49160 567497 49188 641718
rect 49252 585041 49280 660311
rect 49344 655110 49372 661535
rect 49608 660612 49660 660618
rect 49608 660554 49660 660560
rect 49424 660408 49476 660414
rect 49424 660350 49476 660356
rect 49332 655104 49384 655110
rect 49332 655046 49384 655052
rect 49436 649369 49464 660350
rect 49516 660272 49568 660278
rect 49516 660214 49568 660220
rect 49422 649360 49478 649369
rect 49422 649295 49478 649304
rect 49424 648576 49476 648582
rect 49424 648518 49476 648524
rect 49332 629740 49384 629746
rect 49332 629682 49384 629688
rect 49238 585032 49294 585041
rect 49238 584967 49294 584976
rect 49146 567488 49202 567497
rect 49146 567423 49202 567432
rect 49344 544105 49372 629682
rect 49436 561649 49464 648518
rect 49528 643521 49556 660214
rect 49620 655217 49648 660554
rect 49884 660340 49936 660346
rect 49884 660282 49936 660288
rect 49896 659705 49924 660282
rect 49882 659696 49938 659705
rect 49882 659631 49938 659640
rect 49988 658034 50016 661807
rect 50158 661736 50214 661745
rect 50158 661671 50214 661680
rect 50066 661464 50122 661473
rect 50066 661399 50122 661408
rect 49976 658028 50028 658034
rect 49976 657970 50028 657976
rect 49606 655208 49662 655217
rect 49606 655143 49662 655152
rect 49608 655104 49660 655110
rect 49608 655046 49660 655052
rect 49514 643512 49570 643521
rect 49514 643447 49570 643456
rect 49516 594856 49568 594862
rect 49516 594798 49568 594804
rect 49422 561640 49478 561649
rect 49422 561575 49478 561584
rect 49330 544096 49386 544105
rect 49330 544031 49386 544040
rect 49422 532400 49478 532409
rect 49422 532335 49478 532344
rect 48884 499546 49004 499574
rect 48884 497321 48912 499546
rect 48870 497312 48926 497321
rect 48870 497247 48926 497256
rect 48778 468072 48834 468081
rect 48778 468007 48834 468016
rect 48792 467838 48820 468007
rect 48780 467832 48832 467838
rect 48780 467774 48832 467780
rect 48320 445732 48372 445738
rect 48320 445674 48372 445680
rect 48332 444689 48360 445674
rect 48318 444680 48374 444689
rect 48318 444615 48374 444624
rect 48320 438864 48372 438870
rect 48318 438832 48320 438841
rect 48372 438832 48374 438841
rect 48318 438767 48374 438776
rect 48226 409592 48282 409601
rect 48226 409527 48282 409536
rect 46848 397520 46900 397526
rect 3422 397488 3478 397497
rect 46848 397462 46900 397468
rect 3422 397423 3478 397432
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3436 281450 3464 397423
rect 46756 392012 46808 392018
rect 46756 391954 46808 391960
rect 46664 385076 46716 385082
rect 46664 385018 46716 385024
rect 46572 379568 46624 379574
rect 46572 379510 46624 379516
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3528 281518 3556 306167
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 3516 281512 3568 281518
rect 3516 281454 3568 281460
rect 3424 281444 3476 281450
rect 3424 281386 3476 281392
rect 3620 280158 3648 293111
rect 3608 280152 3660 280158
rect 3608 280094 3660 280100
rect 46584 279993 46612 379510
rect 46676 281994 46704 385018
rect 46664 281988 46716 281994
rect 46664 281930 46716 281936
rect 46768 280129 46796 391954
rect 46860 280673 46888 397462
rect 48318 392048 48374 392057
rect 48318 391983 48320 391992
rect 48372 391983 48374 391992
rect 48320 391954 48372 391960
rect 48318 386200 48374 386209
rect 48318 386135 48374 386144
rect 48332 385082 48360 386135
rect 48320 385076 48372 385082
rect 48320 385018 48372 385024
rect 48226 374504 48282 374513
rect 48226 374439 48282 374448
rect 48134 368656 48190 368665
rect 48134 368591 48190 368600
rect 48042 362808 48098 362817
rect 48042 362743 48098 362752
rect 47950 351112 48006 351121
rect 47950 351047 48006 351056
rect 47858 345264 47914 345273
rect 47858 345199 47914 345208
rect 47872 281353 47900 345199
rect 47858 281344 47914 281353
rect 47858 281279 47914 281288
rect 47964 281217 47992 351047
rect 47950 281208 48006 281217
rect 47950 281143 48006 281152
rect 48056 280974 48084 362743
rect 48044 280968 48096 280974
rect 48044 280910 48096 280916
rect 46846 280664 46902 280673
rect 46846 280599 46902 280608
rect 48148 280537 48176 368591
rect 48134 280528 48190 280537
rect 48134 280463 48190 280472
rect 46754 280120 46810 280129
rect 46754 280055 46810 280064
rect 48240 280022 48268 374439
rect 48686 298480 48742 298489
rect 48686 298415 48742 298424
rect 48700 281110 48728 298415
rect 48778 292632 48834 292641
rect 48778 292567 48834 292576
rect 48688 281104 48740 281110
rect 48688 281046 48740 281052
rect 48792 280906 48820 292567
rect 48780 280900 48832 280906
rect 48780 280842 48832 280848
rect 48228 280016 48280 280022
rect 46570 279984 46626 279993
rect 48228 279958 48280 279964
rect 46570 279919 46626 279928
rect 3424 276684 3476 276690
rect 3424 276626 3476 276632
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 2780 150340 2832 150346
rect 2780 150282 2832 150288
rect 2792 149841 2820 150282
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3436 97617 3464 276626
rect 7564 275324 7616 275330
rect 7564 275266 7616 275272
rect 3700 273964 3752 273970
rect 3700 273906 3752 273912
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3514 224224 3570 224233
rect 3514 224159 3570 224168
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3424 85060 3476 85066
rect 3424 85002 3476 85008
rect 3436 84697 3464 85002
rect 3422 84688 3478 84697
rect 3422 84623 3478 84632
rect 3528 58585 3556 224159
rect 3608 220108 3660 220114
rect 3608 220050 3660 220056
rect 3620 136785 3648 220050
rect 3712 201929 3740 273906
rect 4804 272536 4856 272542
rect 4804 272478 4856 272484
rect 3792 224256 3844 224262
rect 3792 224198 3844 224204
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3804 188873 3832 224198
rect 3790 188864 3846 188873
rect 3790 188799 3846 188808
rect 4816 150346 4844 272478
rect 4804 150340 4856 150346
rect 4804 150282 4856 150288
rect 3606 136776 3662 136785
rect 3606 136711 3662 136720
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2780 21412 2832 21418
rect 2780 21354 2832 21360
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 542 -960 654 480
rect 1412 354 1440 18566
rect 2792 16574 2820 21354
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2792 16546 2912 16574
rect 2884 480 2912 16546
rect 7576 6662 7604 275266
rect 9680 268388 9732 268394
rect 9680 268330 9732 268336
rect 8944 231124 8996 231130
rect 8944 231066 8996 231072
rect 8956 85066 8984 231066
rect 8944 85060 8996 85066
rect 8944 85002 8996 85008
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 268330
rect 13820 267028 13872 267034
rect 13820 266970 13872 266976
rect 13832 16574 13860 266970
rect 31024 227044 31076 227050
rect 31024 226986 31076 226992
rect 13832 16546 14320 16574
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 24214 8936 24270 8945
rect 24214 8871 24270 8880
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19444 480 19472 3402
rect 24228 480 24256 8871
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28920 480 28948 3538
rect 31036 3466 31064 226986
rect 42798 226944 42854 226953
rect 42798 226879 42854 226888
rect 39580 7608 39632 7614
rect 39580 7550 39632 7556
rect 32404 6180 32456 6186
rect 32404 6122 32456 6128
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 32416 480 32444 6122
rect 35992 3460 36044 3466
rect 35992 3402 36044 3408
rect 36004 480 36032 3402
rect 39592 480 39620 7550
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42812 354 42840 226879
rect 48884 173398 48912 497247
rect 49436 481642 49464 532335
rect 49528 491473 49556 594798
rect 49620 573345 49648 655046
rect 50080 648582 50108 661399
rect 50172 652798 50200 661671
rect 50896 661496 50948 661502
rect 50896 661438 50948 661444
rect 50804 661428 50856 661434
rect 50804 661370 50856 661376
rect 50620 661360 50672 661366
rect 50620 661302 50672 661308
rect 50344 661224 50396 661230
rect 50344 661166 50396 661172
rect 50252 660000 50304 660006
rect 50252 659942 50304 659948
rect 50264 659705 50292 659942
rect 50250 659696 50306 659705
rect 50250 659631 50306 659640
rect 50252 658028 50304 658034
rect 50252 657970 50304 657976
rect 50160 652792 50212 652798
rect 50160 652734 50212 652740
rect 50068 648576 50120 648582
rect 50068 648518 50120 648524
rect 50264 641782 50292 657970
rect 50252 641776 50304 641782
rect 50252 641718 50304 641724
rect 49606 573336 49662 573345
rect 49606 573271 49662 573280
rect 50356 554742 50384 661166
rect 50528 661156 50580 661162
rect 50528 661098 50580 661104
rect 50436 660476 50488 660482
rect 50436 660418 50488 660424
rect 50448 659841 50476 660418
rect 50434 659832 50490 659841
rect 50434 659767 50490 659776
rect 50540 657642 50568 661098
rect 50448 657614 50568 657642
rect 50448 567186 50476 657614
rect 50528 657552 50580 657558
rect 50528 657494 50580 657500
rect 50540 637537 50568 657494
rect 50526 637528 50582 637537
rect 50526 637463 50582 637472
rect 50436 567180 50488 567186
rect 50436 567122 50488 567128
rect 50344 554736 50396 554742
rect 50344 554678 50396 554684
rect 49606 503160 49662 503169
rect 49606 503095 49662 503104
rect 49514 491464 49570 491473
rect 49514 491399 49570 491408
rect 49424 481636 49476 481642
rect 49424 481578 49476 481584
rect 48962 473920 49018 473929
rect 48962 473855 49018 473864
rect 48976 473346 49004 473855
rect 48964 473340 49016 473346
rect 48964 473282 49016 473288
rect 48976 281314 49004 473282
rect 49056 467832 49108 467838
rect 49056 467774 49108 467780
rect 48964 281308 49016 281314
rect 48964 281250 49016 281256
rect 49068 281246 49096 467774
rect 49148 433288 49200 433294
rect 49148 433230 49200 433236
rect 49160 432993 49188 433230
rect 49146 432984 49202 432993
rect 49146 432919 49202 432928
rect 49422 397896 49478 397905
rect 49422 397831 49478 397840
rect 49436 397526 49464 397831
rect 49424 397520 49476 397526
rect 49424 397462 49476 397468
rect 49422 380352 49478 380361
rect 49422 380287 49478 380296
rect 49436 379574 49464 380287
rect 49424 379568 49476 379574
rect 49424 379510 49476 379516
rect 49422 327720 49478 327729
rect 49422 327655 49478 327664
rect 49330 321872 49386 321881
rect 49330 321807 49386 321816
rect 49238 316024 49294 316033
rect 49238 315959 49294 315968
rect 49146 304328 49202 304337
rect 49146 304263 49202 304272
rect 49160 281926 49188 304263
rect 49148 281920 49200 281926
rect 49148 281862 49200 281868
rect 49056 281240 49108 281246
rect 49056 281182 49108 281188
rect 49252 281042 49280 315959
rect 49240 281036 49292 281042
rect 49240 280978 49292 280984
rect 49344 280770 49372 321807
rect 49436 281081 49464 327655
rect 49422 281072 49478 281081
rect 49422 281007 49478 281016
rect 49332 280764 49384 280770
rect 49332 280706 49384 280712
rect 48962 224360 49018 224369
rect 48962 224295 49018 224304
rect 48872 173392 48924 173398
rect 48872 173334 48924 173340
rect 46664 3664 46716 3670
rect 46664 3606 46716 3612
rect 46676 480 46704 3606
rect 48976 3466 49004 224295
rect 49528 169726 49556 491399
rect 49620 487898 49648 503095
rect 49608 487892 49660 487898
rect 49608 487834 49660 487840
rect 50344 487892 50396 487898
rect 50344 487834 50396 487840
rect 49606 485616 49662 485625
rect 49606 485551 49662 485560
rect 49620 484401 49648 485551
rect 49606 484392 49662 484401
rect 49606 484327 49662 484336
rect 49792 456408 49844 456414
rect 49790 456376 49792 456385
rect 49844 456376 49846 456385
rect 49790 456311 49846 456320
rect 50252 345092 50304 345098
rect 50252 345034 50304 345040
rect 50264 280090 50292 345034
rect 50252 280084 50304 280090
rect 50252 280026 50304 280032
rect 50356 176662 50384 487834
rect 50436 481636 50488 481642
rect 50436 481578 50488 481584
rect 50448 197334 50476 481578
rect 50632 450537 50660 661302
rect 50712 660544 50764 660550
rect 50712 660486 50764 660492
rect 50724 625977 50752 660486
rect 50710 625968 50766 625977
rect 50710 625903 50766 625912
rect 50816 508774 50844 661370
rect 50908 657558 50936 661438
rect 50896 657552 50948 657558
rect 50896 657494 50948 657500
rect 51000 654134 51028 662662
rect 50908 654106 51028 654134
rect 50908 520713 50936 654106
rect 50988 651432 51040 651438
rect 50988 651374 51040 651380
rect 51000 526561 51028 651374
rect 51092 538257 51120 662730
rect 51078 538248 51134 538257
rect 51078 538183 51134 538192
rect 50986 526552 51042 526561
rect 50986 526487 51042 526496
rect 50894 520704 50950 520713
rect 50894 520639 50950 520648
rect 50804 508768 50856 508774
rect 50804 508710 50856 508716
rect 50804 462324 50856 462330
rect 50804 462266 50856 462272
rect 50816 462233 50844 462266
rect 50802 462224 50858 462233
rect 50802 462159 50858 462168
rect 50710 456376 50766 456385
rect 50710 456311 50766 456320
rect 50618 450528 50674 450537
rect 50618 450463 50674 450472
rect 50528 409896 50580 409902
rect 50528 409838 50580 409844
rect 50540 281382 50568 409838
rect 50620 357468 50672 357474
rect 50620 357410 50672 357416
rect 50632 282062 50660 357410
rect 50620 282056 50672 282062
rect 50620 281998 50672 282004
rect 50528 281376 50580 281382
rect 50528 281318 50580 281324
rect 50436 197328 50488 197334
rect 50436 197270 50488 197276
rect 50344 176656 50396 176662
rect 50344 176598 50396 176604
rect 49516 169720 49568 169726
rect 49516 169662 49568 169668
rect 50724 144566 50752 456311
rect 50816 149054 50844 462159
rect 50908 189038 50936 520639
rect 51000 192982 51028 526487
rect 51092 201482 51120 538183
rect 51184 514865 51212 662866
rect 51816 662516 51868 662522
rect 51816 662458 51868 662464
rect 51724 661292 51776 661298
rect 51724 661234 51776 661240
rect 51446 660648 51502 660657
rect 51446 660583 51502 660592
rect 51170 514856 51226 514865
rect 51170 514791 51226 514800
rect 51080 201476 51132 201482
rect 51080 201418 51132 201424
rect 50988 192976 51040 192982
rect 50988 192918 51040 192924
rect 50896 189032 50948 189038
rect 50896 188974 50948 188980
rect 51184 184890 51212 514791
rect 51262 509008 51318 509017
rect 51262 508943 51318 508952
rect 51276 508774 51304 508943
rect 51264 508768 51316 508774
rect 51264 508710 51316 508716
rect 51172 184884 51224 184890
rect 51172 184826 51224 184832
rect 51276 180810 51304 508710
rect 51354 450528 51410 450537
rect 51354 450463 51410 450472
rect 51264 180804 51316 180810
rect 51264 180746 51316 180752
rect 50804 149048 50856 149054
rect 50804 148990 50856 148996
rect 50712 144560 50764 144566
rect 50712 144502 50764 144508
rect 51368 140758 51396 450463
rect 51460 403753 51488 660583
rect 51736 594862 51764 661234
rect 51828 607209 51856 662458
rect 51920 612814 51948 663070
rect 52012 619002 52040 663138
rect 71792 663105 71820 702986
rect 89180 700398 89208 703520
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 105464 697610 105492 703520
rect 137848 700466 137876 703520
rect 154132 700534 154160 703520
rect 202800 700602 202828 703520
rect 202788 700596 202840 700602
rect 202788 700538 202840 700544
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 137836 700460 137888 700466
rect 137836 700402 137888 700408
rect 105452 697604 105504 697610
rect 105452 697546 105504 697552
rect 71778 663096 71834 663105
rect 71778 663031 71834 663040
rect 52184 662992 52236 662998
rect 52184 662934 52236 662940
rect 52092 661836 52144 661842
rect 52092 661778 52144 661784
rect 52104 629746 52132 661778
rect 52196 651438 52224 662934
rect 218072 661774 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 253204 700664 253256 700670
rect 253204 700606 253256 700612
rect 218060 661768 218112 661774
rect 218060 661710 218112 661716
rect 52184 651432 52236 651438
rect 52184 651374 52236 651380
rect 52092 629740 52144 629746
rect 52092 629682 52144 629688
rect 52000 618996 52052 619002
rect 52000 618938 52052 618944
rect 51908 612808 51960 612814
rect 51908 612750 51960 612756
rect 51814 607200 51870 607209
rect 51814 607135 51870 607144
rect 51724 594856 51776 594862
rect 51724 594798 51776 594804
rect 253216 562358 253244 700606
rect 253296 700596 253348 700602
rect 253296 700538 253348 700544
rect 253308 595474 253336 700538
rect 260104 700528 260156 700534
rect 260104 700470 260156 700476
rect 253388 700460 253440 700466
rect 253388 700402 253440 700408
rect 253400 596902 253428 700402
rect 254766 658200 254822 658209
rect 254766 658135 254822 658144
rect 254582 652352 254638 652361
rect 254582 652287 254638 652296
rect 254306 646504 254362 646513
rect 254306 646439 254362 646448
rect 254320 645930 254348 646439
rect 254308 645924 254360 645930
rect 254308 645866 254360 645872
rect 254306 640656 254362 640665
rect 254306 640591 254362 640600
rect 254320 640490 254348 640591
rect 254308 640484 254360 640490
rect 254308 640426 254360 640432
rect 254398 617264 254454 617273
rect 254398 617199 254454 617208
rect 254412 616894 254440 617199
rect 254400 616888 254452 616894
rect 254400 616830 254452 616836
rect 254490 611416 254546 611425
rect 254490 611351 254492 611360
rect 254544 611351 254546 611360
rect 254492 611322 254544 611328
rect 254214 605568 254270 605577
rect 254214 605503 254270 605512
rect 254228 604518 254256 605503
rect 254216 604512 254268 604518
rect 254216 604454 254268 604460
rect 254596 599622 254624 652287
rect 254674 634808 254730 634817
rect 254674 634743 254730 634752
rect 254688 633486 254716 634743
rect 254676 633480 254728 633486
rect 254676 633422 254728 633428
rect 254674 628960 254730 628969
rect 254674 628895 254730 628904
rect 254688 627978 254716 628895
rect 254676 627972 254728 627978
rect 254676 627914 254728 627920
rect 254674 623112 254730 623121
rect 254674 623047 254730 623056
rect 254584 599616 254636 599622
rect 254584 599558 254636 599564
rect 253388 596896 253440 596902
rect 253388 596838 253440 596844
rect 253296 595468 253348 595474
rect 253296 595410 253348 595416
rect 254490 593872 254546 593881
rect 254490 593807 254546 593816
rect 254504 593434 254532 593807
rect 254492 593428 254544 593434
rect 254492 593370 254544 593376
rect 254582 588024 254638 588033
rect 254582 587959 254584 587968
rect 254636 587959 254638 587968
rect 254584 587930 254636 587936
rect 253938 582176 253994 582185
rect 253938 582111 253994 582120
rect 253952 581330 253980 582111
rect 253940 581324 253992 581330
rect 253940 581266 253992 581272
rect 254214 576328 254270 576337
rect 254214 576263 254270 576272
rect 254228 575550 254256 576263
rect 254216 575544 254268 575550
rect 254216 575486 254268 575492
rect 253938 570480 253994 570489
rect 253938 570415 253994 570424
rect 253952 570042 253980 570415
rect 253940 570036 253992 570042
rect 253940 569978 253992 569984
rect 254582 564632 254638 564641
rect 254582 564567 254638 564576
rect 254596 564466 254624 564567
rect 254584 564460 254636 564466
rect 254584 564402 254636 564408
rect 253204 562352 253256 562358
rect 253204 562294 253256 562300
rect 254582 558784 254638 558793
rect 254582 558719 254638 558728
rect 254596 557598 254624 558719
rect 254584 557592 254636 557598
rect 254584 557534 254636 557540
rect 254582 552936 254638 552945
rect 254582 552871 254638 552880
rect 254596 552090 254624 552871
rect 254584 552084 254636 552090
rect 254584 552026 254636 552032
rect 254582 547088 254638 547097
rect 254582 547023 254638 547032
rect 254596 546514 254624 547023
rect 254584 546508 254636 546514
rect 254584 546450 254636 546456
rect 254688 545086 254716 623047
rect 254780 598942 254808 658135
rect 257344 645924 257396 645930
rect 257344 645866 257396 645872
rect 254858 599720 254914 599729
rect 254858 599655 254914 599664
rect 254768 598936 254820 598942
rect 254768 598878 254820 598884
rect 254872 592686 254900 599655
rect 254860 592680 254912 592686
rect 254860 592622 254912 592628
rect 255964 581324 256016 581330
rect 255964 581266 256016 581272
rect 254676 545080 254728 545086
rect 254676 545022 254728 545028
rect 254398 541240 254454 541249
rect 254398 541175 254454 541184
rect 254412 541006 254440 541175
rect 254400 541000 254452 541006
rect 254400 540942 254452 540948
rect 254582 535392 254638 535401
rect 254582 535327 254638 535336
rect 254596 534138 254624 535327
rect 254584 534132 254636 534138
rect 254584 534074 254636 534080
rect 254582 529544 254638 529553
rect 254582 529479 254638 529488
rect 254596 528630 254624 529479
rect 254584 528624 254636 528630
rect 254584 528566 254636 528572
rect 254306 523696 254362 523705
rect 254306 523631 254362 523640
rect 254320 523054 254348 523631
rect 254308 523048 254360 523054
rect 254308 522990 254360 522996
rect 254582 517848 254638 517857
rect 254582 517783 254584 517792
rect 254636 517783 254638 517792
rect 254584 517754 254636 517760
rect 254398 512000 254454 512009
rect 254398 511935 254454 511944
rect 254412 510678 254440 511935
rect 254400 510672 254452 510678
rect 254400 510614 254452 510620
rect 254306 506152 254362 506161
rect 254306 506087 254362 506096
rect 254320 505170 254348 506087
rect 254308 505164 254360 505170
rect 254308 505106 254360 505112
rect 254582 500304 254638 500313
rect 254582 500239 254638 500248
rect 254596 499594 254624 500239
rect 254584 499588 254636 499594
rect 254584 499530 254636 499536
rect 254582 494456 254638 494465
rect 254582 494391 254638 494400
rect 254596 494086 254624 494391
rect 254584 494080 254636 494086
rect 254584 494022 254636 494028
rect 254582 488608 254638 488617
rect 254582 488543 254584 488552
rect 254636 488543 254638 488552
rect 254584 488514 254636 488520
rect 254582 482760 254638 482769
rect 254582 482695 254638 482704
rect 254596 481710 254624 482695
rect 254584 481704 254636 481710
rect 254584 481646 254636 481652
rect 254214 476912 254270 476921
rect 254214 476847 254270 476856
rect 254228 476134 254256 476847
rect 254216 476128 254268 476134
rect 254216 476070 254268 476076
rect 254582 471064 254638 471073
rect 254582 470999 254638 471008
rect 254596 470626 254624 470999
rect 254584 470620 254636 470626
rect 254584 470562 254636 470568
rect 254582 465216 254638 465225
rect 254582 465151 254638 465160
rect 254596 465118 254624 465151
rect 254584 465112 254636 465118
rect 254584 465054 254636 465060
rect 254582 459368 254638 459377
rect 254582 459303 254638 459312
rect 254596 458250 254624 459303
rect 254584 458244 254636 458250
rect 254584 458186 254636 458192
rect 254306 453520 254362 453529
rect 254306 453455 254362 453464
rect 254320 452674 254348 453455
rect 254308 452668 254360 452674
rect 254308 452610 254360 452616
rect 254674 447672 254730 447681
rect 254674 447607 254730 447616
rect 254688 447166 254716 447607
rect 254676 447160 254728 447166
rect 254676 447102 254728 447108
rect 254398 441824 254454 441833
rect 254398 441759 254400 441768
rect 254452 441759 254454 441768
rect 254400 441730 254452 441736
rect 254398 435976 254454 435985
rect 254398 435911 254454 435920
rect 254412 434790 254440 435911
rect 254400 434784 254452 434790
rect 254400 434726 254452 434732
rect 254582 430128 254638 430137
rect 254582 430063 254638 430072
rect 254596 429214 254624 430063
rect 254584 429208 254636 429214
rect 254584 429150 254636 429156
rect 254582 424280 254638 424289
rect 254582 424215 254638 424224
rect 254596 423706 254624 424215
rect 254584 423700 254636 423706
rect 254584 423642 254636 423648
rect 254582 418432 254638 418441
rect 254582 418367 254638 418376
rect 254596 418198 254624 418367
rect 254584 418192 254636 418198
rect 254584 418134 254636 418140
rect 254582 412584 254638 412593
rect 254582 412519 254638 412528
rect 254596 411330 254624 412519
rect 254584 411324 254636 411330
rect 254584 411266 254636 411272
rect 254582 406736 254638 406745
rect 254582 406671 254638 406680
rect 51446 403744 51502 403753
rect 51446 403679 51502 403688
rect 254030 400888 254086 400897
rect 254030 400823 254086 400832
rect 254044 400246 254072 400823
rect 254032 400240 254084 400246
rect 254032 400182 254084 400188
rect 254398 383344 254454 383353
rect 254398 383279 254454 383288
rect 254412 382294 254440 383279
rect 254400 382288 254452 382294
rect 254400 382230 254452 382236
rect 254122 377496 254178 377505
rect 254122 377431 254178 377440
rect 254136 376786 254164 377431
rect 254124 376780 254176 376786
rect 254124 376722 254176 376728
rect 253938 359952 253994 359961
rect 253938 359887 253994 359896
rect 253952 358902 253980 359887
rect 253940 358896 253992 358902
rect 253940 358838 253992 358844
rect 51446 356960 51502 356969
rect 51446 356895 51502 356904
rect 51460 282033 51488 356895
rect 254214 354104 254270 354113
rect 254214 354039 254270 354048
rect 254228 353326 254256 354039
rect 254216 353320 254268 353326
rect 254216 353262 254268 353268
rect 254490 348256 254546 348265
rect 254490 348191 254546 348200
rect 254504 347818 254532 348191
rect 254492 347812 254544 347818
rect 254492 347754 254544 347760
rect 254596 342922 254624 406671
rect 254674 395040 254730 395049
rect 254674 394975 254730 394984
rect 254688 394806 254716 394975
rect 254676 394800 254728 394806
rect 254676 394742 254728 394748
rect 254676 389224 254728 389230
rect 254674 389192 254676 389201
rect 254728 389192 254730 389201
rect 254674 389127 254730 389136
rect 254674 371648 254730 371657
rect 254674 371583 254730 371592
rect 254688 371278 254716 371583
rect 254676 371272 254728 371278
rect 254676 371214 254728 371220
rect 254674 365800 254730 365809
rect 254674 365735 254676 365744
rect 254728 365735 254730 365744
rect 254676 365706 254728 365712
rect 254584 342916 254636 342922
rect 254584 342858 254636 342864
rect 254582 342408 254638 342417
rect 254582 342343 254638 342352
rect 254596 342310 254624 342343
rect 254584 342304 254636 342310
rect 254584 342246 254636 342252
rect 51538 339416 51594 339425
rect 51538 339351 51594 339360
rect 51446 282024 51502 282033
rect 51446 281959 51502 281968
rect 51552 280945 51580 339351
rect 254398 336560 254454 336569
rect 254398 336495 254454 336504
rect 254412 335374 254440 336495
rect 254400 335368 254452 335374
rect 254400 335310 254452 335316
rect 51722 333568 51778 333577
rect 51722 333503 51778 333512
rect 51630 310176 51686 310185
rect 51630 310111 51686 310120
rect 51644 281897 51672 310111
rect 51630 281888 51686 281897
rect 51630 281823 51686 281832
rect 51538 280936 51594 280945
rect 51538 280871 51594 280880
rect 51736 280809 51764 333503
rect 253296 331696 253348 331702
rect 253296 331638 253348 331644
rect 253204 331356 253256 331362
rect 253204 331298 253256 331304
rect 52090 286512 52146 286521
rect 52090 286447 52146 286456
rect 52104 281178 52132 286447
rect 53104 281308 53156 281314
rect 53104 281250 53156 281256
rect 52092 281172 52144 281178
rect 52092 281114 52144 281120
rect 51722 280800 51778 280809
rect 51722 280735 51778 280744
rect 53116 157350 53144 281250
rect 54484 281240 54536 281246
rect 54484 281182 54536 281188
rect 54576 281240 54628 281246
rect 54576 281182 54628 281188
rect 53104 157344 53156 157350
rect 53104 157286 53156 157292
rect 54496 153202 54524 281182
rect 54588 280974 54616 281182
rect 54576 280968 54628 280974
rect 54576 280910 54628 280916
rect 59358 279440 59414 279449
rect 59358 279375 59414 279384
rect 54574 278760 54630 278769
rect 54574 278695 54630 278704
rect 54588 161430 54616 278695
rect 59268 276752 59320 276758
rect 59268 276694 59320 276700
rect 58900 272604 58952 272610
rect 58900 272546 58952 272552
rect 58808 233912 58860 233918
rect 58808 233854 58860 233860
rect 57336 228472 57388 228478
rect 57336 228414 57388 228420
rect 55862 223544 55918 223553
rect 55862 223479 55918 223488
rect 55876 164393 55904 223479
rect 57060 222896 57112 222902
rect 57060 222838 57112 222844
rect 57072 217433 57100 222838
rect 57244 221536 57296 221542
rect 57244 221478 57296 221484
rect 57152 220244 57204 220250
rect 57152 220186 57204 220192
rect 57058 217424 57114 217433
rect 57058 217359 57114 217368
rect 57164 209273 57192 220186
rect 57256 214606 57284 221478
rect 57244 214600 57296 214606
rect 57244 214542 57296 214548
rect 57150 209264 57206 209273
rect 57150 209199 57206 209208
rect 57348 205193 57376 228414
rect 57796 225616 57848 225622
rect 57796 225558 57848 225564
rect 57520 222964 57572 222970
rect 57520 222906 57572 222912
rect 57428 218816 57480 218822
rect 57428 218758 57480 218764
rect 57334 205184 57390 205193
rect 57334 205119 57390 205128
rect 57336 201476 57388 201482
rect 57336 201418 57388 201424
rect 57348 201113 57376 201418
rect 57334 201104 57390 201113
rect 57334 201039 57390 201048
rect 57336 197328 57388 197334
rect 57336 197270 57388 197276
rect 57348 197033 57376 197270
rect 57334 197024 57390 197033
rect 57334 196959 57390 196968
rect 57336 192976 57388 192982
rect 57334 192944 57336 192953
rect 57388 192944 57390 192953
rect 57334 192879 57390 192888
rect 57336 189032 57388 189038
rect 57336 188974 57388 188980
rect 57348 188873 57376 188974
rect 57334 188864 57390 188873
rect 57334 188799 57390 188808
rect 56692 184884 56744 184890
rect 56692 184826 56744 184832
rect 56704 184793 56732 184826
rect 56690 184784 56746 184793
rect 56690 184719 56746 184728
rect 56692 180804 56744 180810
rect 56692 180746 56744 180752
rect 56704 180713 56732 180746
rect 56690 180704 56746 180713
rect 56690 180639 56746 180648
rect 57336 176656 57388 176662
rect 57334 176624 57336 176633
rect 57388 176624 57390 176633
rect 57334 176559 57390 176568
rect 57244 173392 57296 173398
rect 57244 173334 57296 173340
rect 57256 172553 57284 173334
rect 57242 172544 57298 172553
rect 57242 172479 57298 172488
rect 57336 169720 57388 169726
rect 57336 169662 57388 169668
rect 57348 168473 57376 169662
rect 57334 168464 57390 168473
rect 57334 168399 57390 168408
rect 55862 164384 55918 164393
rect 55862 164319 55918 164328
rect 54576 161424 54628 161430
rect 54576 161366 54628 161372
rect 57060 161424 57112 161430
rect 57060 161366 57112 161372
rect 57072 160313 57100 161366
rect 57058 160304 57114 160313
rect 57058 160239 57114 160248
rect 57060 157344 57112 157350
rect 57060 157286 57112 157292
rect 57072 156233 57100 157286
rect 57058 156224 57114 156233
rect 57058 156159 57114 156168
rect 54484 153196 54536 153202
rect 54484 153138 54536 153144
rect 57336 153196 57388 153202
rect 57336 153138 57388 153144
rect 57348 152153 57376 153138
rect 57334 152144 57390 152153
rect 57334 152079 57390 152088
rect 57336 149048 57388 149054
rect 57336 148990 57388 148996
rect 57348 148073 57376 148990
rect 57334 148064 57390 148073
rect 57334 147999 57390 148008
rect 57336 144560 57388 144566
rect 57336 144502 57388 144508
rect 57348 143993 57376 144502
rect 57334 143984 57390 143993
rect 57334 143919 57390 143928
rect 57440 142154 57468 218758
rect 57348 142126 57468 142154
rect 51356 140752 51408 140758
rect 51356 140694 51408 140700
rect 57348 135833 57376 142126
rect 57428 140752 57480 140758
rect 57428 140694 57480 140700
rect 57440 139913 57468 140694
rect 57426 139904 57482 139913
rect 57426 139839 57482 139848
rect 57334 135824 57390 135833
rect 57334 135759 57390 135768
rect 57532 123593 57560 222906
rect 57612 218748 57664 218754
rect 57612 218690 57664 218696
rect 57518 123584 57574 123593
rect 57518 123519 57574 123528
rect 57624 107273 57652 218690
rect 57704 214600 57756 214606
rect 57704 214542 57756 214548
rect 57610 107264 57666 107273
rect 57610 107199 57666 107208
rect 57716 103193 57744 214542
rect 57702 103184 57758 103193
rect 57702 103119 57758 103128
rect 57808 86873 57836 225558
rect 58716 221468 58768 221474
rect 58716 221410 58768 221416
rect 57888 218884 57940 218890
rect 57888 218826 57940 218832
rect 57794 86864 57850 86873
rect 57794 86799 57850 86808
rect 57900 78713 57928 218826
rect 58728 111353 58756 221410
rect 58820 119513 58848 233854
rect 58912 127673 58940 272546
rect 59084 253224 59136 253230
rect 59084 253166 59136 253172
rect 58992 236700 59044 236706
rect 58992 236642 59044 236648
rect 58898 127664 58954 127673
rect 58898 127599 58954 127608
rect 58806 119504 58862 119513
rect 58806 119439 58862 119448
rect 58714 111344 58770 111353
rect 58714 111279 58770 111288
rect 59004 82793 59032 236642
rect 59096 90953 59124 253166
rect 59176 225684 59228 225690
rect 59176 225626 59228 225632
rect 59082 90944 59138 90953
rect 59082 90879 59138 90888
rect 58990 82784 59046 82793
rect 58990 82719 59046 82728
rect 57886 78704 57942 78713
rect 57886 78639 57942 78648
rect 59188 62393 59216 225626
rect 59280 99113 59308 276694
rect 59266 99104 59322 99113
rect 59266 99039 59322 99048
rect 59372 70553 59400 279375
rect 59452 278044 59504 278050
rect 59452 277986 59504 277992
rect 59464 115433 59492 277986
rect 59636 235272 59688 235278
rect 59636 235214 59688 235220
rect 59544 228404 59596 228410
rect 59544 228346 59596 228352
rect 59450 115424 59506 115433
rect 59450 115359 59506 115368
rect 59358 70544 59414 70553
rect 59358 70479 59414 70488
rect 59556 66473 59584 228346
rect 59648 74633 59676 235214
rect 60004 229764 60056 229770
rect 60004 229706 60056 229712
rect 59726 225584 59782 225593
rect 59726 225519 59782 225528
rect 59740 95033 59768 225519
rect 59726 95024 59782 95033
rect 59726 94959 59782 94968
rect 59634 74624 59690 74633
rect 59634 74559 59690 74568
rect 59542 66464 59598 66473
rect 59542 66399 59598 66408
rect 59174 62384 59230 62393
rect 59174 62319 59230 62328
rect 53746 4856 53802 4865
rect 50160 4820 50212 4826
rect 53746 4791 53802 4800
rect 50160 4762 50212 4768
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 50172 480 50200 4762
rect 53760 480 53788 4791
rect 60016 3534 60044 229706
rect 222844 222284 222896 222290
rect 222844 222226 222896 222232
rect 60556 220176 60608 220182
rect 60556 220118 60608 220124
rect 60568 213897 60596 220118
rect 222856 215665 222884 222226
rect 224408 222216 224460 222222
rect 224408 222158 224460 222164
rect 222936 216708 222988 216714
rect 222936 216650 222988 216656
rect 222842 215656 222898 215665
rect 222842 215591 222898 215600
rect 60554 213888 60610 213897
rect 60554 213823 60610 213832
rect 222292 213036 222344 213042
rect 222292 212978 222344 212984
rect 222304 212809 222332 212978
rect 222290 212800 222346 212809
rect 222290 212735 222346 212744
rect 222948 207097 222976 216650
rect 223210 209944 223266 209953
rect 223210 209879 223266 209888
rect 222934 207088 222990 207097
rect 222934 207023 222990 207032
rect 223224 205630 223252 209879
rect 223212 205624 223264 205630
rect 223212 205566 223264 205572
rect 222842 204232 222898 204241
rect 222842 204167 222898 204176
rect 222856 190466 222884 204167
rect 223026 201376 223082 201385
rect 223026 201311 223082 201320
rect 222934 198520 222990 198529
rect 222934 198455 222990 198464
rect 222844 190460 222896 190466
rect 222844 190402 222896 190408
rect 222948 186318 222976 198455
rect 223040 189038 223068 201311
rect 224316 197396 224368 197402
rect 224316 197338 224368 197344
rect 224224 196036 224276 196042
rect 224224 195978 224276 195984
rect 223486 195664 223542 195673
rect 223486 195599 223542 195608
rect 223500 194614 223528 195599
rect 223488 194608 223540 194614
rect 223488 194550 223540 194556
rect 223486 192808 223542 192817
rect 223486 192743 223542 192752
rect 223500 191894 223528 192743
rect 223488 191888 223540 191894
rect 223488 191830 223540 191836
rect 223486 189952 223542 189961
rect 223486 189887 223542 189896
rect 223500 189106 223528 189887
rect 223488 189100 223540 189106
rect 223488 189042 223540 189048
rect 223028 189032 223080 189038
rect 223028 188974 223080 188980
rect 223486 187096 223542 187105
rect 223486 187031 223542 187040
rect 223500 186386 223528 187031
rect 223488 186380 223540 186386
rect 223488 186322 223540 186328
rect 222936 186312 222988 186318
rect 222936 186254 222988 186260
rect 222290 184240 222346 184249
rect 222290 184175 222292 184184
rect 222344 184175 222346 184184
rect 222292 184146 222344 184152
rect 223486 181384 223542 181393
rect 223486 181319 223542 181328
rect 222658 178528 222714 178537
rect 222658 178463 222714 178472
rect 222672 176662 222700 178463
rect 223500 178022 223528 181319
rect 223488 178016 223540 178022
rect 223488 177958 223540 177964
rect 222660 176656 222712 176662
rect 222660 176598 222712 176604
rect 222658 175672 222714 175681
rect 222658 175607 222714 175616
rect 222672 175234 222700 175607
rect 222660 175228 222712 175234
rect 222660 175170 222712 175176
rect 222384 173188 222436 173194
rect 222384 173130 222436 173136
rect 222396 172825 222424 173130
rect 222382 172816 222438 172825
rect 222382 172751 222438 172760
rect 222476 171148 222528 171154
rect 222476 171090 222528 171096
rect 222488 169969 222516 171090
rect 222474 169960 222530 169969
rect 222474 169895 222530 169904
rect 222936 169788 222988 169794
rect 222936 169730 222988 169736
rect 222948 167113 222976 169730
rect 222934 167104 222990 167113
rect 222934 167039 222990 167048
rect 223488 167068 223540 167074
rect 223488 167010 223540 167016
rect 223028 165640 223080 165646
rect 223028 165582 223080 165588
rect 222936 164280 222988 164286
rect 222936 164222 222988 164228
rect 222948 158545 222976 164222
rect 223040 161401 223068 165582
rect 223500 164257 223528 167010
rect 223486 164248 223542 164257
rect 223486 164183 223542 164192
rect 223488 162920 223540 162926
rect 223488 162862 223540 162868
rect 223026 161392 223082 161401
rect 223026 161327 223082 161336
rect 222934 158536 222990 158545
rect 222934 158471 222990 158480
rect 222660 157344 222712 157350
rect 222660 157286 222712 157292
rect 222672 152833 222700 157286
rect 223500 155689 223528 162862
rect 223486 155680 223542 155689
rect 223486 155615 223542 155624
rect 222936 154624 222988 154630
rect 222936 154566 222988 154572
rect 222844 153264 222896 153270
rect 222844 153206 222896 153212
rect 222658 152824 222714 152833
rect 222658 152759 222714 152768
rect 222568 147144 222620 147150
rect 222566 147112 222568 147121
rect 222620 147112 222622 147121
rect 222566 147047 222622 147056
rect 222660 137964 222712 137970
rect 222660 137906 222712 137912
rect 222672 132841 222700 137906
rect 222856 135697 222884 153206
rect 222948 138553 222976 154566
rect 223212 151088 223264 151094
rect 223212 151030 223264 151036
rect 223224 149977 223252 151030
rect 223210 149968 223266 149977
rect 223210 149903 223266 149912
rect 223488 144900 223540 144906
rect 223488 144842 223540 144848
rect 223500 144265 223528 144842
rect 223486 144256 223542 144265
rect 223486 144191 223542 144200
rect 223488 141500 223540 141506
rect 223488 141442 223540 141448
rect 223500 141409 223528 141442
rect 223486 141400 223542 141409
rect 223486 141335 223542 141344
rect 222934 138544 222990 138553
rect 222934 138479 222990 138488
rect 222842 135688 222898 135697
rect 222842 135623 222898 135632
rect 222844 133204 222896 133210
rect 222844 133146 222896 133152
rect 222658 132832 222714 132841
rect 222658 132767 222714 132776
rect 222292 128308 222344 128314
rect 222292 128250 222344 128256
rect 222304 124273 222332 128250
rect 222856 127129 222884 133146
rect 223028 130076 223080 130082
rect 223028 130018 223080 130024
rect 223040 129985 223068 130018
rect 223026 129976 223082 129985
rect 223026 129911 223082 129920
rect 222842 127120 222898 127129
rect 222842 127055 222898 127064
rect 222290 124264 222346 124273
rect 222290 124199 222346 124208
rect 223486 121408 223542 121417
rect 223486 121343 223542 121352
rect 223500 120698 223528 121343
rect 223488 120692 223540 120698
rect 223488 120634 223540 120640
rect 223488 118652 223540 118658
rect 223488 118594 223540 118600
rect 223500 118561 223528 118594
rect 223486 118552 223542 118561
rect 223486 118487 223542 118496
rect 223488 115932 223540 115938
rect 223488 115874 223540 115880
rect 223500 115705 223528 115874
rect 223486 115696 223542 115705
rect 223486 115631 223542 115640
rect 222200 113008 222252 113014
rect 222200 112950 222252 112956
rect 222212 112849 222240 112950
rect 222198 112840 222254 112849
rect 222198 112775 222254 112784
rect 223488 110424 223540 110430
rect 223488 110366 223540 110372
rect 223500 109993 223528 110366
rect 223486 109984 223542 109993
rect 223486 109919 223542 109928
rect 222660 107636 222712 107642
rect 222660 107578 222712 107584
rect 222672 107137 222700 107578
rect 222658 107128 222714 107137
rect 222658 107063 222714 107072
rect 222844 104848 222896 104854
rect 222844 104790 222896 104796
rect 222856 104281 222884 104790
rect 222842 104272 222898 104281
rect 222842 104207 222898 104216
rect 223488 102128 223540 102134
rect 223488 102070 223540 102076
rect 223500 101425 223528 102070
rect 223486 101416 223542 101425
rect 223486 101351 223542 101360
rect 223028 99340 223080 99346
rect 223028 99282 223080 99288
rect 223040 98569 223068 99282
rect 223026 98560 223082 98569
rect 223026 98495 223082 98504
rect 223120 96620 223172 96626
rect 223120 96562 223172 96568
rect 223132 95713 223160 96562
rect 223118 95704 223174 95713
rect 223118 95639 223174 95648
rect 223488 93832 223540 93838
rect 223488 93774 223540 93780
rect 223500 92857 223528 93774
rect 223486 92848 223542 92857
rect 223486 92783 223542 92792
rect 223488 91792 223540 91798
rect 223488 91734 223540 91740
rect 223500 90001 223528 91734
rect 223486 89992 223542 90001
rect 223486 89927 223542 89936
rect 223212 88324 223264 88330
rect 223212 88266 223264 88272
rect 223224 87145 223252 88266
rect 223210 87136 223266 87145
rect 223210 87071 223266 87080
rect 223212 85536 223264 85542
rect 223212 85478 223264 85484
rect 223224 84289 223252 85478
rect 223210 84280 223266 84289
rect 223210 84215 223266 84224
rect 223486 81424 223542 81433
rect 223486 81359 223488 81368
rect 223540 81359 223542 81368
rect 223488 81330 223540 81336
rect 222476 78600 222528 78606
rect 222474 78568 222476 78577
rect 222528 78568 222530 78577
rect 222474 78503 222530 78512
rect 222200 75744 222252 75750
rect 222198 75712 222200 75721
rect 222252 75712 222254 75721
rect 222198 75647 222254 75656
rect 224236 73098 224264 195978
rect 224328 75750 224356 197338
rect 224420 113014 224448 222158
rect 226064 220856 226116 220862
rect 226064 220798 226116 220804
rect 226076 213042 226104 220798
rect 253216 218890 253244 331298
rect 253308 222970 253336 331638
rect 254582 331528 254638 331537
rect 254582 331463 254638 331472
rect 254214 330712 254270 330721
rect 254214 330647 254270 330656
rect 254228 329934 254256 330647
rect 254216 329928 254268 329934
rect 254216 329870 254268 329876
rect 254492 325644 254544 325650
rect 254492 325586 254544 325592
rect 254504 324873 254532 325586
rect 254490 324864 254546 324873
rect 254490 324799 254546 324808
rect 254308 320136 254360 320142
rect 254308 320078 254360 320084
rect 254320 319025 254348 320078
rect 254306 319016 254362 319025
rect 254306 318951 254362 318960
rect 254214 307320 254270 307329
rect 254214 307255 254270 307264
rect 254228 306406 254256 307255
rect 254216 306400 254268 306406
rect 254216 306342 254268 306348
rect 254398 289776 254454 289785
rect 254398 289711 254454 289720
rect 254412 288454 254440 289711
rect 254400 288448 254452 288454
rect 254400 288390 254452 288396
rect 254306 283928 254362 283937
rect 254306 283863 254362 283872
rect 254320 282946 254348 283863
rect 254308 282940 254360 282946
rect 254308 282882 254360 282888
rect 253296 222964 253348 222970
rect 253296 222906 253348 222912
rect 254596 221542 254624 331463
rect 254676 329860 254728 329866
rect 254676 329802 254728 329808
rect 254688 313177 254716 329802
rect 254674 313168 254730 313177
rect 254674 313103 254730 313112
rect 254674 301472 254730 301481
rect 254674 301407 254730 301416
rect 254688 300898 254716 301407
rect 254676 300892 254728 300898
rect 254676 300834 254728 300840
rect 254674 295624 254730 295633
rect 254674 295559 254730 295568
rect 254688 295390 254716 295559
rect 254676 295384 254728 295390
rect 254676 295326 254728 295332
rect 254584 221536 254636 221542
rect 254584 221478 254636 221484
rect 253204 218884 253256 218890
rect 253204 218826 253256 218832
rect 247684 215348 247736 215354
rect 247684 215290 247736 215296
rect 246304 213988 246356 213994
rect 246304 213930 246356 213936
rect 226064 213036 226116 213042
rect 226064 212978 226116 212984
rect 242164 212560 242216 212566
rect 242164 212502 242216 212508
rect 239404 211200 239456 211206
rect 239404 211142 239456 211148
rect 238024 209840 238076 209846
rect 238024 209782 238076 209788
rect 235264 208412 235316 208418
rect 235264 208354 235316 208360
rect 229744 205624 229796 205630
rect 229744 205566 229796 205572
rect 228364 200184 228416 200190
rect 228364 200126 228416 200132
rect 225604 198756 225656 198762
rect 225604 198698 225656 198704
rect 224408 113008 224460 113014
rect 224408 112950 224460 112956
rect 225616 78606 225644 198698
rect 225696 184204 225748 184210
rect 225696 184146 225748 184152
rect 225708 179382 225736 184146
rect 225696 179376 225748 179382
rect 225696 179318 225748 179324
rect 225788 158772 225840 158778
rect 225788 158714 225840 158720
rect 225800 147150 225828 158714
rect 225788 147144 225840 147150
rect 225788 147086 225840 147092
rect 225696 146328 225748 146334
rect 225696 146270 225748 146276
rect 225708 128314 225736 146270
rect 225696 128308 225748 128314
rect 225696 128250 225748 128256
rect 228376 81394 228404 200126
rect 229756 193186 229784 205566
rect 233976 194608 234028 194614
rect 233976 194550 234028 194556
rect 229744 193180 229796 193186
rect 229744 193122 229796 193128
rect 232504 191888 232556 191894
rect 232504 191830 232556 191836
rect 230388 189100 230440 189106
rect 230388 189042 230440 189048
rect 230400 182170 230428 189042
rect 232516 183530 232544 191830
rect 233884 190528 233936 190534
rect 233884 190470 233936 190476
rect 232504 183524 232556 183530
rect 232504 183466 232556 183472
rect 230388 182164 230440 182170
rect 230388 182106 230440 182112
rect 229100 161492 229152 161498
rect 229100 161434 229152 161440
rect 229112 157350 229140 161434
rect 232596 157412 232648 157418
rect 232596 157354 232648 157360
rect 229100 157344 229152 157350
rect 229100 157286 229152 157292
rect 229836 155984 229888 155990
rect 229836 155926 229888 155932
rect 228456 149116 228508 149122
rect 228456 149058 228508 149064
rect 228468 130082 228496 149058
rect 229744 144968 229796 144974
rect 229744 144910 229796 144916
rect 228456 130076 228508 130082
rect 228456 130018 228508 130024
rect 229756 120698 229784 144910
rect 229848 141506 229876 155926
rect 231124 151836 231176 151842
rect 231124 151778 231176 151784
rect 229836 141500 229888 141506
rect 229836 141442 229888 141448
rect 231136 137970 231164 151778
rect 232608 144906 232636 157354
rect 232596 144900 232648 144906
rect 232596 144842 232648 144848
rect 232504 143608 232556 143614
rect 232504 143550 232556 143556
rect 231124 137964 231176 137970
rect 231124 137906 231176 137912
rect 229744 120692 229796 120698
rect 229744 120634 229796 120640
rect 232516 118658 232544 143550
rect 232504 118652 232556 118658
rect 232504 118594 232556 118600
rect 228364 81388 228416 81394
rect 228364 81330 228416 81336
rect 225604 78600 225656 78606
rect 225604 78542 225656 78548
rect 224316 75744 224368 75750
rect 224316 75686 224368 75692
rect 222200 73092 222252 73098
rect 222200 73034 222252 73040
rect 224224 73092 224276 73098
rect 224224 73034 224276 73040
rect 222212 72865 222240 73034
rect 222198 72856 222254 72865
rect 222198 72791 222254 72800
rect 223488 70372 223540 70378
rect 223488 70314 223540 70320
rect 223500 70009 223528 70314
rect 223486 70000 223542 70009
rect 223486 69935 223542 69944
rect 223488 67584 223540 67590
rect 223488 67526 223540 67532
rect 223500 67153 223528 67526
rect 223486 67144 223542 67153
rect 223486 67079 223542 67088
rect 233896 64870 233924 190470
rect 233988 184890 234016 194550
rect 233976 184884 234028 184890
rect 233976 184826 234028 184832
rect 235276 96626 235304 208354
rect 238036 99346 238064 209782
rect 239416 102134 239444 211142
rect 242176 104854 242204 212502
rect 243544 193248 243596 193254
rect 243544 193190 243596 193196
rect 242164 104848 242216 104854
rect 242164 104790 242216 104796
rect 239404 102128 239456 102134
rect 239404 102070 239456 102076
rect 238024 99340 238076 99346
rect 238024 99282 238076 99288
rect 235264 96620 235316 96626
rect 235264 96562 235316 96568
rect 243556 67590 243584 193190
rect 246316 107642 246344 213930
rect 247696 110430 247724 215290
rect 253204 201544 253256 201550
rect 253204 201486 253256 201492
rect 250444 194608 250496 194614
rect 250444 194550 250496 194556
rect 247684 110424 247736 110430
rect 247684 110366 247736 110372
rect 246304 107636 246356 107642
rect 246304 107578 246356 107584
rect 250456 70378 250484 194550
rect 253216 85542 253244 201486
rect 253204 85536 253256 85542
rect 253204 85478 253256 85484
rect 255976 75886 256004 581266
rect 256056 570036 256108 570042
rect 256056 569978 256108 569984
rect 255964 75880 256016 75886
rect 255964 75822 256016 75828
rect 256068 73166 256096 569978
rect 256148 497548 256200 497554
rect 256148 497490 256200 497496
rect 256160 228478 256188 497490
rect 256240 358896 256292 358902
rect 256240 358838 256292 358844
rect 256252 306338 256280 358838
rect 256240 306332 256292 306338
rect 256240 306274 256292 306280
rect 256148 228472 256200 228478
rect 256148 228414 256200 228420
rect 257356 142118 257384 645866
rect 257436 640484 257488 640490
rect 257436 640426 257488 640432
rect 257344 142112 257396 142118
rect 257344 142054 257396 142060
rect 257448 140758 257476 640426
rect 260116 591326 260144 700470
rect 267660 694822 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 694816 267700 694822
rect 267648 694758 267700 694764
rect 276664 663196 276716 663202
rect 276664 663138 276716 663144
rect 269856 633480 269908 633486
rect 269856 633422 269908 633428
rect 264244 616888 264296 616894
rect 264244 616830 264296 616836
rect 260104 591320 260156 591326
rect 260104 591262 260156 591268
rect 260104 587988 260156 587994
rect 260104 587930 260156 587936
rect 258724 517812 258776 517818
rect 258724 517754 258776 517760
rect 257620 497480 257672 497486
rect 257620 497422 257672 497428
rect 257528 441788 257580 441794
rect 257528 441730 257580 441736
rect 257436 140752 257488 140758
rect 257436 140694 257488 140700
rect 257540 113150 257568 441730
rect 257632 227089 257660 497422
rect 257618 227080 257674 227089
rect 257618 227015 257674 227024
rect 258736 132462 258764 517754
rect 258816 497684 258868 497690
rect 258816 497626 258868 497632
rect 258828 218822 258856 497626
rect 258816 218816 258868 218822
rect 258816 218758 258868 218764
rect 258724 132456 258776 132462
rect 258724 132398 258776 132404
rect 257528 113144 257580 113150
rect 257528 113086 257580 113092
rect 260116 77246 260144 587930
rect 261484 546508 261536 546514
rect 261484 546450 261536 546456
rect 260196 545080 260248 545086
rect 260196 545022 260248 545028
rect 260208 86970 260236 545022
rect 260288 394800 260340 394806
rect 260288 394742 260340 394748
rect 260300 307766 260328 394742
rect 260840 334620 260892 334626
rect 260840 334562 260892 334568
rect 260288 307760 260340 307766
rect 260288 307702 260340 307708
rect 260196 86964 260248 86970
rect 260196 86906 260248 86912
rect 260104 77240 260156 77246
rect 260104 77182 260156 77188
rect 256056 73160 256108 73166
rect 256056 73102 256108 73108
rect 250444 70372 250496 70378
rect 250444 70314 250496 70320
rect 243544 67584 243596 67590
rect 243544 67526 243596 67532
rect 222844 64864 222896 64870
rect 222844 64806 222896 64812
rect 233884 64864 233936 64870
rect 233884 64806 233936 64812
rect 222856 64297 222884 64806
rect 222842 64288 222898 64297
rect 222842 64223 222898 64232
rect 165618 61568 165674 61577
rect 165618 61503 165674 61512
rect 215300 61532 215352 61538
rect 158720 61464 158772 61470
rect 126978 61432 127034 61441
rect 158720 61406 158772 61412
rect 126978 61367 127034 61376
rect 154580 61396 154632 61402
rect 99380 42084 99432 42090
rect 99380 42026 99432 42032
rect 85580 35216 85632 35222
rect 85580 35158 85632 35164
rect 77300 32428 77352 32434
rect 77300 32370 77352 32376
rect 74540 31068 74592 31074
rect 74540 31010 74592 31016
rect 63500 26920 63552 26926
rect 63500 26862 63552 26868
rect 60740 25560 60792 25566
rect 60740 25502 60792 25508
rect 60752 16574 60780 25502
rect 63512 16574 63540 26862
rect 74552 16574 74580 31010
rect 77312 16574 77340 32370
rect 85592 16574 85620 35158
rect 92478 24168 92534 24177
rect 92478 24103 92534 24112
rect 60752 16546 60872 16574
rect 63512 16546 64368 16574
rect 74552 16546 75040 16574
rect 77312 16546 78168 16574
rect 85592 16546 85712 16574
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 60004 3528 60056 3534
rect 60004 3470 60056 3476
rect 57256 480 57284 3470
rect 60844 480 60872 16546
rect 64340 480 64368 16546
rect 71502 7576 71558 7585
rect 71502 7511 71558 7520
rect 67914 6216 67970 6225
rect 67914 6151 67970 6160
rect 67928 480 67956 6151
rect 71516 480 71544 7511
rect 75012 480 75040 16546
rect 43046 354 43158 480
rect 42812 326 43158 354
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78140 354 78168 16546
rect 82084 8968 82136 8974
rect 82084 8910 82136 8916
rect 82096 480 82124 8910
rect 85684 480 85712 16546
rect 89168 3460 89220 3466
rect 89168 3402 89220 3408
rect 89180 480 89208 3402
rect 78558 354 78670 480
rect 78140 326 78670 354
rect 78558 -960 78670 326
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92492 354 92520 24103
rect 99392 16574 99420 42026
rect 120080 40724 120132 40730
rect 120080 40666 120132 40672
rect 113180 28280 113232 28286
rect 113180 28222 113232 28228
rect 113192 16574 113220 28222
rect 120092 16574 120120 40666
rect 99392 16546 99880 16574
rect 113192 16546 114048 16574
rect 120092 16546 120672 16574
rect 95792 15904 95844 15910
rect 95792 15846 95844 15852
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 95804 354 95832 15846
rect 99852 480 99880 16546
rect 102140 14476 102192 14482
rect 102140 14418 102192 14424
rect 102152 3534 102180 14418
rect 110512 9036 110564 9042
rect 110512 8978 110564 8984
rect 102140 3528 102192 3534
rect 102140 3470 102192 3476
rect 103336 3528 103388 3534
rect 103336 3470 103388 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 103348 480 103376 3470
rect 106936 480 106964 3470
rect 110524 480 110552 8978
rect 114020 480 114048 16546
rect 117596 3800 117648 3806
rect 117596 3742 117648 3748
rect 117608 480 117636 3742
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 124680 3732 124732 3738
rect 124680 3674 124732 3680
rect 124692 480 124720 3674
rect 126992 480 127020 61367
rect 154580 61338 154632 61344
rect 133880 60036 133932 60042
rect 133880 59978 133932 59984
rect 129738 55856 129794 55865
rect 129738 55791 129794 55800
rect 129752 16574 129780 55791
rect 129752 16546 130608 16574
rect 130580 480 130608 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 133892 354 133920 59978
rect 136638 59936 136694 59945
rect 136638 59871 136694 59880
rect 136652 16574 136680 59871
rect 151820 58744 151872 58750
rect 151820 58686 151872 58692
rect 140780 58676 140832 58682
rect 140780 58618 140832 58624
rect 140792 16574 140820 58618
rect 147678 57216 147734 57225
rect 147678 57151 147734 57160
rect 147692 16574 147720 57151
rect 136652 16546 137232 16574
rect 140792 16546 141280 16574
rect 147692 16546 147904 16574
rect 134126 354 134238 480
rect 133892 326 134238 354
rect 134126 -960 134238 326
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137204 354 137232 16546
rect 141252 480 141280 16546
rect 144734 5128 144790 5137
rect 144734 5063 144790 5072
rect 144748 480 144776 5063
rect 137622 354 137734 480
rect 137204 326 137734 354
rect 137622 -960 137734 326
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 151832 480 151860 58686
rect 154592 16574 154620 61338
rect 158732 16574 158760 61406
rect 165632 16574 165660 61503
rect 215300 61474 215352 61480
rect 211160 60240 211212 60246
rect 211160 60182 211212 60188
rect 197360 60172 197412 60178
rect 197360 60114 197412 60120
rect 168380 60104 168432 60110
rect 168380 60046 168432 60052
rect 154592 16546 155448 16574
rect 158732 16546 158944 16574
rect 165632 16546 166120 16574
rect 155420 480 155448 16546
rect 158916 480 158944 16546
rect 162490 3360 162546 3369
rect 162490 3295 162546 3304
rect 162504 480 162532 3295
rect 166092 480 166120 16546
rect 168392 3398 168420 60046
rect 172520 58812 172572 58818
rect 172520 58754 172572 58760
rect 172532 16574 172560 58754
rect 179420 57316 179472 57322
rect 179420 57258 179472 57264
rect 176660 57248 176712 57254
rect 176660 57190 176712 57196
rect 172532 16546 172744 16574
rect 168380 3392 168432 3398
rect 168380 3334 168432 3340
rect 169576 3392 169628 3398
rect 169576 3334 169628 3340
rect 169588 480 169616 3334
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 176672 480 176700 57190
rect 179432 16574 179460 57258
rect 190460 55888 190512 55894
rect 190460 55830 190512 55836
rect 186318 39264 186374 39273
rect 186318 39199 186374 39208
rect 186332 16574 186360 39199
rect 179432 16546 180288 16574
rect 186332 16546 186912 16574
rect 180260 480 180288 16546
rect 183742 3496 183798 3505
rect 183742 3431 183798 3440
rect 183756 480 183784 3431
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 55830
rect 193220 42152 193272 42158
rect 193220 42094 193272 42100
rect 193232 3398 193260 42094
rect 197372 16574 197400 60114
rect 201500 47592 201552 47598
rect 201500 47534 201552 47540
rect 197372 16546 197952 16574
rect 193220 3392 193272 3398
rect 193220 3334 193272 3340
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 194428 480 194456 3334
rect 197924 480 197952 16546
rect 201512 480 201540 47534
rect 204260 44872 204312 44878
rect 204260 44814 204312 44820
rect 204272 16574 204300 44814
rect 211172 16574 211200 60182
rect 204272 16546 205128 16574
rect 211172 16546 211752 16574
rect 205100 480 205128 16546
rect 208584 4888 208636 4894
rect 208584 4830 208636 4836
rect 208596 480 208624 4830
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 61474
rect 247040 58880 247092 58886
rect 247040 58822 247092 58828
rect 233240 57384 233292 57390
rect 233240 57326 233292 57332
rect 218060 54528 218112 54534
rect 218060 54470 218112 54476
rect 218072 3398 218100 54470
rect 226340 53100 226392 53106
rect 226340 53042 226392 53048
rect 222200 42220 222252 42226
rect 222200 42162 222252 42168
rect 222212 16574 222240 42162
rect 222212 16546 222792 16574
rect 218060 3392 218112 3398
rect 218060 3334 218112 3340
rect 219256 3392 219308 3398
rect 219256 3334 219308 3340
rect 219268 480 219296 3334
rect 222764 480 222792 16546
rect 226352 480 226380 53042
rect 233252 16574 233280 57326
rect 236000 55956 236052 55962
rect 236000 55898 236052 55904
rect 236012 16574 236040 55898
rect 242900 46232 242952 46238
rect 242900 46174 242952 46180
rect 233252 16546 233464 16574
rect 236012 16546 236592 16574
rect 229836 7676 229888 7682
rect 229836 7618 229888 7624
rect 229848 480 229876 7618
rect 233436 480 233464 16546
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 16546
rect 240140 10328 240192 10334
rect 240140 10270 240192 10276
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 354 240180 10270
rect 242912 3398 242940 46174
rect 247052 16574 247080 58822
rect 251180 51740 251232 51746
rect 251180 51682 251232 51688
rect 247052 16546 247632 16574
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 244108 480 244136 3334
rect 247604 480 247632 16546
rect 251192 480 251220 51682
rect 260852 16574 260880 334562
rect 261496 67590 261524 546450
rect 262864 499588 262916 499594
rect 262864 499530 262916 499536
rect 261576 494080 261628 494086
rect 261576 494022 261628 494028
rect 261588 126954 261616 494022
rect 262876 128314 262904 499530
rect 262864 128308 262916 128314
rect 262864 128250 262916 128256
rect 261576 126948 261628 126954
rect 261576 126890 261628 126896
rect 264256 89010 264284 616830
rect 269764 592680 269816 592686
rect 269764 592622 269816 592628
rect 265624 557592 265676 557598
rect 265624 557534 265676 557540
rect 264980 493332 265032 493338
rect 264980 493274 265032 493280
rect 264336 470620 264388 470626
rect 264336 470562 264388 470568
rect 264348 121446 264376 470562
rect 264428 282940 264480 282946
rect 264428 282882 264480 282888
rect 264336 121440 264388 121446
rect 264336 121382 264388 121388
rect 264244 89004 264296 89010
rect 264244 88946 264296 88952
rect 261484 67584 261536 67590
rect 261484 67526 261536 67532
rect 264440 62082 264468 282882
rect 264428 62076 264480 62082
rect 264428 62018 264480 62024
rect 260852 16546 261800 16574
rect 258264 13116 258316 13122
rect 258264 13058 258316 13064
rect 254674 4992 254730 5001
rect 254674 4927 254730 4936
rect 254688 480 254716 4927
rect 258276 480 258304 13058
rect 261772 480 261800 16546
rect 240478 354 240590 480
rect 240152 326 240590 354
rect 240478 -960 240590 326
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 354 265020 493274
rect 265636 70378 265664 557534
rect 268384 552084 268436 552090
rect 268384 552026 268436 552032
rect 267004 541000 267056 541006
rect 267004 540942 267056 540948
rect 265716 476128 265768 476134
rect 265716 476070 265768 476076
rect 265728 122806 265756 476070
rect 265716 122800 265768 122806
rect 265716 122742 265768 122748
rect 267016 90370 267044 540942
rect 267096 497616 267148 497622
rect 267096 497558 267148 497564
rect 267108 222902 267136 497558
rect 267740 487824 267792 487830
rect 267740 487766 267792 487772
rect 267096 222896 267148 222902
rect 267096 222838 267148 222844
rect 267004 90364 267056 90370
rect 267004 90306 267056 90312
rect 265624 70372 265676 70378
rect 265624 70314 265676 70320
rect 267752 16574 267780 487766
rect 268396 69018 268424 552026
rect 268476 481704 268528 481710
rect 268476 481646 268528 481652
rect 268488 124166 268516 481646
rect 268476 124160 268528 124166
rect 268476 124102 268528 124108
rect 269776 80034 269804 592622
rect 269868 139398 269896 633422
rect 275376 627972 275428 627978
rect 275376 627914 275428 627920
rect 273904 611380 273956 611386
rect 273904 611322 273956 611328
rect 271144 604512 271196 604518
rect 271144 604454 271196 604460
rect 269948 505164 270000 505170
rect 269948 505106 270000 505112
rect 269856 139392 269908 139398
rect 269856 139334 269908 139340
rect 269960 129742 269988 505106
rect 269948 129736 270000 129742
rect 269948 129678 270000 129684
rect 271156 82822 271184 604454
rect 272522 542872 272578 542881
rect 272522 542807 272578 542816
rect 271236 510672 271288 510678
rect 271236 510614 271288 510620
rect 271248 131102 271276 510614
rect 271328 465112 271380 465118
rect 271328 465054 271380 465060
rect 271236 131096 271288 131102
rect 271236 131038 271288 131044
rect 271340 120086 271368 465054
rect 271880 340264 271932 340270
rect 271880 340206 271932 340212
rect 271328 120080 271380 120086
rect 271328 120022 271380 120028
rect 271144 82816 271196 82822
rect 271144 82758 271196 82764
rect 269764 80028 269816 80034
rect 269764 79970 269816 79976
rect 268384 69012 268436 69018
rect 268384 68954 268436 68960
rect 271892 16574 271920 340206
rect 272536 280974 272564 542807
rect 272524 280968 272576 280974
rect 272524 280910 272576 280916
rect 273916 84182 273944 611322
rect 275284 593428 275336 593434
rect 275284 593370 275336 593376
rect 273996 528624 274048 528630
rect 273996 528566 274048 528572
rect 274008 136610 274036 528566
rect 274088 523048 274140 523054
rect 274088 522990 274140 522996
rect 273996 136604 274048 136610
rect 273996 136546 274048 136552
rect 274100 135250 274128 522990
rect 274088 135244 274140 135250
rect 274088 135186 274140 135192
rect 273904 84176 273956 84182
rect 273904 84118 273956 84124
rect 275296 78674 275324 593370
rect 275388 137970 275416 627914
rect 276676 543114 276704 663138
rect 276756 663128 276808 663134
rect 276756 663070 276808 663076
rect 276768 543386 276796 663070
rect 276848 663060 276900 663066
rect 276848 663002 276900 663008
rect 276860 545902 276888 663002
rect 279516 661836 279568 661842
rect 279516 661778 279568 661784
rect 278136 660612 278188 660618
rect 278136 660554 278188 660560
rect 278044 575544 278096 575550
rect 278044 575486 278096 575492
rect 276848 545896 276900 545902
rect 276848 545838 276900 545844
rect 276756 543380 276808 543386
rect 276756 543322 276808 543328
rect 276664 543108 276716 543114
rect 276664 543050 276716 543056
rect 276664 539640 276716 539646
rect 276664 539582 276716 539588
rect 276020 486464 276072 486470
rect 276020 486406 276072 486412
rect 275468 447160 275520 447166
rect 275468 447102 275520 447108
rect 275376 137964 275428 137970
rect 275376 137906 275428 137912
rect 275480 114510 275508 447102
rect 275468 114504 275520 114510
rect 275468 114446 275520 114452
rect 275284 78668 275336 78674
rect 275284 78610 275336 78616
rect 267752 16546 268424 16574
rect 271892 16546 272472 16574
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 272444 480 272472 16546
rect 276032 480 276060 486406
rect 276676 281042 276704 539582
rect 276664 281036 276716 281042
rect 276664 280978 276716 280984
rect 278056 74526 278084 575486
rect 278148 543182 278176 660554
rect 279148 660408 279200 660414
rect 279148 660350 279200 660356
rect 278688 641028 278740 641034
rect 278688 640970 278740 640976
rect 278700 610065 278728 640970
rect 278780 638988 278832 638994
rect 278780 638930 278832 638936
rect 278792 630057 278820 638930
rect 278778 630048 278834 630057
rect 278778 629983 278834 629992
rect 278686 610056 278742 610065
rect 278686 609991 278742 610000
rect 279160 543318 279188 660350
rect 279332 660204 279384 660210
rect 279332 660146 279384 660152
rect 279240 660136 279292 660142
rect 279240 660078 279292 660084
rect 279252 543522 279280 660078
rect 279344 543590 279372 660146
rect 279424 564460 279476 564466
rect 279424 564402 279476 564408
rect 279332 543584 279384 543590
rect 279332 543526 279384 543532
rect 279240 543516 279292 543522
rect 279240 543458 279292 543464
rect 279148 543312 279200 543318
rect 279148 543254 279200 543260
rect 278136 543176 278188 543182
rect 278136 543118 278188 543124
rect 278320 542428 278372 542434
rect 278320 542370 278372 542376
rect 278136 534132 278188 534138
rect 278136 534074 278188 534080
rect 278044 74520 278096 74526
rect 278044 74462 278096 74468
rect 278148 64870 278176 534074
rect 278228 458244 278280 458250
rect 278228 458186 278280 458192
rect 278240 118658 278268 458186
rect 278332 281926 278360 542370
rect 278780 498840 278832 498846
rect 278780 498782 278832 498788
rect 278320 281920 278372 281926
rect 278320 281862 278372 281868
rect 278228 118652 278280 118658
rect 278228 118594 278280 118600
rect 278136 64864 278188 64870
rect 278136 64806 278188 64812
rect 278792 16574 278820 498782
rect 279436 71738 279464 564402
rect 279528 543454 279556 661778
rect 279608 661632 279660 661638
rect 279608 661574 279660 661580
rect 279620 545766 279648 661574
rect 279700 660544 279752 660550
rect 279700 660486 279752 660492
rect 279974 660512 280030 660521
rect 279712 545834 279740 660486
rect 279974 660447 280030 660456
rect 279884 660068 279936 660074
rect 279884 660010 279936 660016
rect 279700 545828 279752 545834
rect 279700 545770 279752 545776
rect 279608 545760 279660 545766
rect 279608 545702 279660 545708
rect 279896 543726 279924 660010
rect 279884 543720 279936 543726
rect 279884 543662 279936 543668
rect 279516 543448 279568 543454
rect 279516 543390 279568 543396
rect 279988 543046 280016 660447
rect 280068 660272 280120 660278
rect 280068 660214 280120 660220
rect 280080 543250 280108 660214
rect 282932 643754 282960 702406
rect 300136 700369 300164 703520
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 317420 700460 317472 700466
rect 317420 700402 317472 700408
rect 300122 700360 300178 700369
rect 300122 700295 300178 700304
rect 316132 683188 316184 683194
rect 316132 683130 316184 683136
rect 310520 661564 310572 661570
rect 310520 661506 310572 661512
rect 310532 661473 310560 661506
rect 310518 661464 310574 661473
rect 310518 661399 310574 661408
rect 316144 654134 316172 683130
rect 317432 654134 317460 700402
rect 331232 660414 331260 702986
rect 348804 700602 348832 703520
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 397472 698970 397500 703520
rect 409236 700596 409288 700602
rect 409236 700538 409288 700544
rect 405004 700528 405056 700534
rect 405004 700470 405056 700476
rect 397460 698964 397512 698970
rect 397460 698906 397512 698912
rect 337384 697604 337436 697610
rect 337384 697546 337436 697552
rect 331220 660408 331272 660414
rect 331220 660350 331272 660356
rect 316144 654106 316724 654134
rect 317432 654106 317828 654134
rect 282920 643748 282972 643754
rect 282920 643690 282972 643696
rect 287612 642388 287664 642394
rect 287612 642330 287664 642336
rect 286508 642116 286560 642122
rect 286508 642058 286560 642064
rect 282092 642048 282144 642054
rect 282092 641990 282144 641996
rect 282104 639962 282132 641990
rect 282736 641980 282788 641986
rect 282736 641922 282788 641928
rect 281796 639934 282132 639962
rect 282748 639826 282776 641922
rect 284208 641912 284260 641918
rect 284208 641854 284260 641860
rect 284220 639962 284248 641854
rect 286520 639962 286548 642058
rect 287624 639962 287652 642330
rect 293776 642320 293828 642326
rect 293776 642262 293828 642268
rect 310058 642288 310114 642297
rect 284004 639934 284248 639962
rect 286212 639934 286548 639962
rect 287316 639934 287652 639962
rect 293788 639826 293816 642262
rect 300768 642252 300820 642258
rect 310058 642223 310114 642232
rect 300768 642194 300820 642200
rect 295248 642184 295300 642190
rect 295248 642126 295300 642132
rect 295260 639962 295288 642126
rect 297548 641844 297600 641850
rect 297548 641786 297600 641792
rect 297560 639962 297588 641786
rect 299296 641776 299348 641782
rect 299296 641718 299348 641724
rect 295044 639934 295288 639962
rect 297252 639934 297588 639962
rect 299308 639826 299336 641718
rect 300780 639962 300808 642194
rect 310072 641034 310100 642223
rect 310060 641028 310112 641034
rect 310060 640970 310112 640976
rect 315856 641028 315908 641034
rect 315856 640970 315908 640976
rect 314108 640960 314160 640966
rect 314108 640902 314160 640908
rect 313004 640688 313056 640694
rect 307482 640656 307538 640665
rect 313004 640630 313056 640636
rect 307482 640591 307538 640600
rect 309692 640620 309744 640626
rect 304816 640552 304868 640558
rect 304170 640520 304226 640529
rect 301964 640484 302016 640490
rect 304816 640494 304868 640500
rect 304170 640455 304226 640464
rect 301964 640426 302016 640432
rect 301976 639962 302004 640426
rect 304184 639962 304212 640455
rect 300564 639934 300808 639962
rect 301668 639934 302004 639962
rect 303876 639934 304212 639962
rect 304828 639962 304856 640494
rect 307496 639962 307524 640591
rect 309692 640562 309744 640568
rect 309704 639962 309732 640562
rect 310336 640348 310388 640354
rect 310336 640290 310388 640296
rect 304828 639934 304980 639962
rect 307188 639934 307524 639962
rect 309396 639934 309732 639962
rect 310348 639962 310376 640290
rect 313016 639962 313044 640630
rect 314120 639962 314148 640902
rect 315212 640416 315264 640422
rect 315212 640358 315264 640364
rect 315224 639962 315252 640358
rect 310348 639934 310500 639962
rect 312708 639934 313044 639962
rect 313812 639934 314148 639962
rect 314916 639934 315252 639962
rect 315868 639826 315896 640970
rect 316696 639962 316724 654106
rect 317800 639962 317828 654106
rect 327724 642524 327776 642530
rect 327724 642466 327776 642472
rect 321192 642320 321244 642326
rect 321192 642262 321244 642268
rect 319536 642048 319588 642054
rect 319536 641990 319588 641996
rect 316696 639934 317124 639962
rect 317800 639934 318228 639962
rect 282748 639798 282900 639826
rect 293788 639798 293940 639826
rect 299308 639798 299460 639826
rect 315868 639798 316020 639826
rect 308586 639432 308642 639441
rect 302772 639402 303108 639418
rect 302772 639396 303120 639402
rect 302772 639390 303068 639396
rect 308292 639390 308586 639418
rect 308586 639367 308642 639376
rect 303068 639338 303120 639344
rect 296444 639328 296496 639334
rect 285402 639296 285458 639305
rect 280172 639254 280692 639282
rect 285108 639254 285402 639282
rect 280172 559609 280200 639254
rect 285402 639231 285458 639240
rect 288254 639296 288310 639305
rect 289634 639296 289690 639305
rect 288310 639254 288420 639282
rect 289524 639254 289634 639282
rect 288254 639231 288310 639240
rect 290922 639296 290978 639305
rect 290628 639254 290922 639282
rect 289634 639231 289690 639240
rect 292026 639296 292082 639305
rect 291732 639254 292026 639282
rect 290922 639231 290978 639240
rect 293130 639296 293186 639305
rect 292836 639254 293130 639282
rect 292026 639231 292082 639240
rect 296148 639276 296444 639282
rect 306288 639328 306340 639334
rect 298466 639296 298522 639305
rect 296148 639270 296496 639276
rect 296148 639254 296484 639270
rect 298356 639254 298466 639282
rect 293130 639231 293186 639240
rect 306084 639276 306288 639282
rect 311716 639328 311768 639334
rect 306084 639270 306340 639276
rect 311604 639276 311716 639282
rect 311604 639270 311768 639276
rect 306084 639254 306328 639270
rect 311604 639254 311756 639270
rect 319332 639254 319484 639282
rect 298466 639231 298522 639240
rect 303434 600672 303490 600681
rect 303324 600630 303434 600658
rect 304722 600672 304778 600681
rect 304428 600630 304722 600658
rect 303434 600607 303490 600616
rect 301410 600536 301466 600545
rect 301116 600494 301410 600522
rect 301410 600471 301466 600480
rect 300674 600128 300730 600137
rect 281552 600086 282348 600114
rect 282472 600086 282900 600114
rect 283024 600086 283452 600114
rect 283668 600086 284004 600114
rect 284312 600086 284556 600114
rect 280158 559600 280214 559609
rect 280158 559535 280214 559544
rect 281552 547874 281580 600086
rect 282472 586514 282500 600086
rect 283024 599010 283052 600086
rect 283012 599004 283064 599010
rect 283012 598946 283064 598952
rect 282920 597100 282972 597106
rect 282920 597042 282972 597048
rect 281644 586486 282500 586514
rect 281644 573345 281672 586486
rect 281630 573336 281686 573345
rect 281630 573271 281686 573280
rect 282932 563689 282960 597042
rect 283024 565146 283052 598946
rect 283668 597106 283696 600086
rect 283656 597100 283708 597106
rect 283656 597042 283708 597048
rect 283012 565140 283064 565146
rect 283012 565082 283064 565088
rect 282918 563680 282974 563689
rect 282918 563615 282974 563624
rect 284312 555490 284340 600086
rect 285094 599842 285122 600100
rect 285232 600086 285660 600114
rect 285876 600086 286212 600114
rect 286764 600086 286916 600114
rect 285094 599814 285168 599842
rect 285140 598466 285168 599814
rect 285128 598460 285180 598466
rect 285128 598402 285180 598408
rect 285232 586514 285260 600086
rect 285876 586514 285904 600086
rect 286888 598670 286916 600086
rect 287164 600086 287316 600114
rect 287532 600086 287868 600114
rect 287992 600086 288420 600114
rect 286876 598664 286928 598670
rect 286876 598606 286928 598612
rect 287060 598188 287112 598194
rect 287060 598130 287112 598136
rect 284404 586486 285260 586514
rect 285692 586486 285904 586514
rect 284404 570654 284432 586486
rect 285692 572082 285720 586486
rect 287072 576230 287100 598130
rect 287164 580281 287192 600086
rect 287532 598194 287560 600086
rect 287520 598188 287572 598194
rect 287520 598130 287572 598136
rect 287992 587178 288020 600086
rect 288958 599842 288986 600100
rect 289096 600086 289524 600114
rect 288958 599814 289032 599842
rect 289004 598398 289032 599814
rect 288992 598392 289044 598398
rect 288992 598334 289044 598340
rect 289096 598210 289124 600086
rect 290062 599842 290090 600100
rect 290200 600086 290628 600114
rect 290062 599814 290136 599842
rect 289176 598664 289228 598670
rect 289176 598606 289228 598612
rect 288452 598182 289124 598210
rect 288452 594114 288480 598182
rect 288440 594108 288492 594114
rect 288440 594050 288492 594056
rect 287980 587172 288032 587178
rect 287980 587114 288032 587120
rect 289188 586514 289216 598606
rect 290108 598262 290136 599814
rect 290096 598256 290148 598262
rect 290096 598198 290148 598204
rect 290200 586514 290228 600086
rect 291166 599842 291194 600100
rect 291120 599814 291194 599842
rect 291396 600086 291732 600114
rect 292284 600086 292528 600114
rect 291120 598194 291148 599814
rect 291108 598188 291160 598194
rect 291108 598130 291160 598136
rect 291396 588606 291424 600086
rect 292500 598670 292528 600086
rect 292684 600086 292836 600114
rect 293388 600086 293540 600114
rect 292488 598664 292540 598670
rect 292488 598606 292540 598612
rect 291844 598188 291896 598194
rect 291844 598130 291896 598136
rect 291384 588600 291436 588606
rect 291384 588542 291436 588548
rect 289096 586486 289216 586514
rect 289832 586486 290228 586514
rect 287150 580272 287206 580281
rect 287150 580207 287206 580216
rect 287060 576224 287112 576230
rect 287060 576166 287112 576172
rect 285680 572076 285732 572082
rect 285680 572018 285732 572024
rect 284392 570648 284444 570654
rect 284392 570590 284444 570596
rect 289096 567866 289124 586486
rect 289084 567860 289136 567866
rect 289084 567802 289136 567808
rect 284300 555484 284352 555490
rect 284300 555426 284352 555432
rect 289832 555393 289860 586486
rect 291856 558210 291884 598130
rect 292580 596080 292632 596086
rect 292580 596022 292632 596028
rect 292592 569226 292620 596022
rect 292684 587217 292712 600086
rect 293512 592686 293540 600086
rect 293604 600086 293940 600114
rect 294156 600086 294492 600114
rect 294616 600086 295044 600114
rect 295352 600086 295596 600114
rect 295812 600086 296148 600114
rect 296364 600086 296700 600114
rect 297252 600086 297588 600114
rect 293604 596086 293632 600086
rect 293592 596080 293644 596086
rect 293592 596022 293644 596028
rect 293500 592680 293552 592686
rect 293500 592622 293552 592628
rect 294156 592034 294184 600086
rect 293972 592006 294184 592034
rect 292670 587208 292726 587217
rect 292670 587143 292726 587152
rect 293972 581670 294000 592006
rect 294616 589966 294644 600086
rect 294604 589960 294656 589966
rect 294604 589902 294656 589908
rect 293960 581664 294012 581670
rect 293960 581606 294012 581612
rect 292580 569220 292632 569226
rect 292580 569162 292632 569168
rect 291844 558204 291896 558210
rect 291844 558146 291896 558152
rect 289818 555384 289874 555393
rect 289818 555319 289874 555328
rect 295352 551410 295380 600086
rect 295812 592034 295840 600086
rect 295444 592006 295840 592034
rect 295340 551404 295392 551410
rect 295340 551346 295392 551352
rect 295444 551342 295472 592006
rect 296364 586514 296392 600086
rect 296720 599888 296772 599894
rect 296720 599830 296772 599836
rect 295536 586486 296392 586514
rect 295536 551478 295564 586486
rect 296732 573442 296760 599830
rect 297456 598664 297508 598670
rect 297456 598606 297508 598612
rect 297468 598398 297496 598606
rect 297456 598392 297508 598398
rect 297456 598334 297508 598340
rect 297560 595542 297588 600086
rect 297790 599894 297818 600100
rect 298356 600086 298692 600114
rect 298908 600086 299336 600114
rect 297778 599888 297830 599894
rect 298100 599888 298152 599894
rect 297830 599836 297864 599842
rect 297778 599830 297864 599836
rect 298100 599830 298152 599836
rect 297790 599814 297864 599830
rect 297836 599282 297864 599814
rect 297824 599276 297876 599282
rect 297824 599218 297876 599224
rect 297548 595536 297600 595542
rect 297548 595478 297600 595484
rect 296720 573436 296772 573442
rect 296720 573378 296772 573384
rect 295524 551472 295576 551478
rect 298112 551449 298140 599830
rect 298664 598126 298692 600086
rect 299308 598913 299336 600086
rect 299446 599894 299474 600100
rect 300012 600086 300348 600114
rect 300564 600086 300674 600114
rect 299434 599888 299486 599894
rect 299400 599836 299434 599842
rect 299400 599830 299486 599836
rect 299400 599814 299474 599830
rect 299400 599078 299428 599814
rect 299388 599072 299440 599078
rect 299388 599014 299440 599020
rect 299294 598904 299350 598913
rect 299294 598839 299350 598848
rect 298652 598120 298704 598126
rect 298652 598062 298704 598068
rect 299308 592034 299336 598839
rect 300320 598058 300348 600086
rect 300730 600086 300808 600114
rect 301668 600086 302096 600114
rect 300674 600063 300730 600072
rect 300688 600003 300716 600063
rect 300676 598120 300728 598126
rect 300676 598062 300728 598068
rect 300308 598052 300360 598058
rect 300308 597994 300360 598000
rect 300584 598052 300636 598058
rect 300584 597994 300636 598000
rect 299308 592006 299428 592034
rect 299400 589937 299428 592006
rect 299386 589928 299442 589937
rect 299386 589863 299442 589872
rect 300596 580417 300624 597994
rect 300582 580408 300638 580417
rect 300582 580343 300638 580352
rect 300688 578921 300716 598062
rect 300674 578912 300730 578921
rect 300674 578847 300730 578856
rect 300780 563718 300808 600086
rect 301964 599956 302016 599962
rect 301964 599898 302016 599904
rect 301976 599214 302004 599898
rect 302068 599842 302096 600086
rect 302206 599962 302234 600100
rect 302772 600086 303108 600114
rect 302194 599956 302246 599962
rect 302194 599898 302246 599904
rect 302068 599814 302188 599842
rect 300860 599208 300912 599214
rect 300860 599150 300912 599156
rect 301964 599208 302016 599214
rect 301964 599150 302016 599156
rect 300872 583001 300900 599150
rect 302160 598874 302188 599814
rect 302148 598868 302200 598874
rect 302148 598810 302200 598816
rect 300858 582992 300914 583001
rect 300858 582927 300914 582936
rect 300768 563712 300820 563718
rect 300768 563654 300820 563660
rect 295524 551414 295576 551420
rect 298098 551440 298154 551449
rect 298098 551375 298154 551384
rect 295432 551336 295484 551342
rect 295432 551278 295484 551284
rect 302160 548554 302188 598810
rect 303080 598398 303108 600086
rect 303068 598392 303120 598398
rect 303068 598334 303120 598340
rect 303448 577590 303476 600607
rect 303876 600086 304212 600114
rect 303528 598800 303580 598806
rect 303528 598742 303580 598748
rect 303540 598398 303568 598742
rect 304184 598534 304212 600086
rect 304172 598528 304224 598534
rect 304172 598470 304224 598476
rect 303528 598392 303580 598398
rect 303528 598334 303580 598340
rect 303620 598392 303672 598398
rect 303620 598334 303672 598340
rect 303436 577584 303488 577590
rect 303436 577526 303488 577532
rect 302148 548548 302200 548554
rect 302148 548490 302200 548496
rect 281540 547868 281592 547874
rect 281540 547810 281592 547816
rect 301872 545896 301924 545902
rect 301872 545838 301924 545844
rect 298192 543720 298244 543726
rect 298192 543662 298244 543668
rect 297086 543416 297142 543425
rect 297086 543351 297142 543360
rect 280068 543244 280120 543250
rect 280068 543186 280120 543192
rect 279976 543040 280028 543046
rect 279976 542982 280028 542988
rect 297100 542881 297128 543351
rect 297454 543144 297510 543153
rect 297454 543079 297510 543088
rect 283470 542872 283526 542881
rect 283470 542807 283526 542816
rect 297086 542872 297142 542881
rect 297086 542807 297142 542816
rect 279700 542632 279752 542638
rect 279700 542574 279752 542580
rect 279608 542564 279660 542570
rect 279608 542506 279660 542512
rect 279516 488572 279568 488578
rect 279516 488514 279568 488520
rect 279528 125594 279556 488514
rect 279620 280022 279648 542506
rect 279712 281246 279740 542574
rect 279792 542496 279844 542502
rect 279792 542438 279844 542444
rect 279804 281994 279832 542438
rect 283484 539866 283512 542807
rect 296902 542736 296958 542745
rect 296902 542671 296958 542680
rect 292764 542564 292816 542570
rect 292764 542506 292816 542512
rect 284944 542428 284996 542434
rect 284944 542370 284996 542376
rect 284956 539866 284984 542370
rect 283484 539838 283820 539866
rect 284956 539838 285292 539866
rect 287886 539744 287942 539753
rect 289358 539744 289414 539753
rect 287942 539702 288236 539730
rect 287886 539679 287942 539688
rect 290830 539744 290886 539753
rect 289414 539702 289708 539730
rect 289358 539679 289414 539688
rect 290886 539702 291180 539730
rect 290830 539679 290886 539688
rect 286416 539640 286468 539646
rect 283378 539608 283434 539617
rect 280804 539572 280856 539578
rect 280804 539514 280856 539520
rect 281460 539566 282348 539594
rect 283084 539566 283378 539594
rect 279792 281988 279844 281994
rect 279792 281930 279844 281936
rect 279700 281240 279752 281246
rect 279700 281182 279752 281188
rect 280816 281110 280844 539514
rect 281460 528554 281488 539566
rect 286138 539608 286194 539617
rect 284220 539578 284556 539594
rect 283378 539543 283434 539552
rect 284208 539572 284556 539578
rect 284260 539566 284556 539572
rect 286028 539566 286138 539594
rect 287610 539608 287666 539617
rect 286468 539588 286764 539594
rect 286416 539582 286764 539588
rect 286428 539566 286764 539582
rect 287500 539566 287610 539594
rect 286138 539543 286194 539552
rect 287610 539543 287666 539552
rect 288622 539608 288678 539617
rect 290738 539608 290794 539617
rect 288678 539566 288972 539594
rect 290444 539566 290738 539594
rect 288622 539543 288678 539552
rect 290738 539543 290794 539552
rect 291566 539608 291622 539617
rect 292776 539594 292804 542506
rect 293960 542496 294012 542502
rect 293960 542438 294012 542444
rect 293972 539866 294000 542438
rect 295340 542428 295392 542434
rect 295340 542370 295392 542376
rect 295352 539866 295380 542370
rect 296916 539866 296944 542671
rect 297468 539866 297496 543079
rect 298204 539866 298232 543662
rect 298928 543584 298980 543590
rect 298928 543526 298980 543532
rect 298940 539866 298968 543526
rect 299664 543516 299716 543522
rect 299664 543458 299716 543464
rect 299676 539866 299704 543458
rect 300398 543280 300454 543289
rect 300398 543215 300454 543224
rect 300412 539866 300440 543215
rect 301134 542872 301190 542881
rect 301134 542807 301190 542816
rect 301148 539866 301176 542807
rect 301884 539866 301912 545838
rect 302608 543448 302660 543454
rect 302608 543390 302660 543396
rect 302620 539866 302648 543390
rect 303540 540258 303568 598334
rect 303632 598126 303660 598334
rect 304184 598126 304212 598470
rect 303620 598120 303672 598126
rect 303620 598062 303672 598068
rect 304172 598120 304224 598126
rect 304172 598062 304224 598068
rect 304644 551546 304672 600630
rect 306194 600672 306250 600681
rect 306084 600630 306194 600658
rect 304722 600607 304778 600616
rect 306194 600607 306250 600616
rect 304966 599842 304994 600100
rect 305532 600086 305868 600114
rect 304920 599814 304994 599842
rect 304920 598670 304948 599814
rect 304908 598664 304960 598670
rect 304908 598606 304960 598612
rect 304920 598346 304948 598606
rect 305840 598602 305868 600086
rect 305828 598596 305880 598602
rect 305828 598538 305880 598544
rect 304736 598318 304948 598346
rect 304736 585886 304764 598318
rect 304816 598120 304868 598126
rect 304816 598062 304868 598068
rect 304724 585880 304776 585886
rect 304724 585822 304776 585828
rect 304828 574802 304856 598062
rect 304816 574796 304868 574802
rect 304816 574738 304868 574744
rect 306208 565214 306236 600607
rect 306636 600086 306788 600114
rect 306760 599146 306788 600086
rect 306852 600086 307188 600114
rect 307404 600086 307740 600114
rect 306380 599140 306432 599146
rect 306380 599082 306432 599088
rect 306748 599140 306800 599146
rect 306748 599082 306800 599088
rect 306288 598596 306340 598602
rect 306288 598538 306340 598544
rect 306196 565208 306248 565214
rect 306196 565150 306248 565156
rect 304632 551540 304684 551546
rect 304632 551482 304684 551488
rect 304998 543416 305054 543425
rect 304080 543380 304132 543386
rect 304998 543351 305054 543360
rect 304080 543322 304132 543328
rect 303620 543108 303672 543114
rect 303620 543050 303672 543056
rect 303528 540252 303580 540258
rect 303528 540194 303580 540200
rect 303632 540138 303660 543050
rect 303632 540110 303706 540138
rect 293972 539838 294124 539866
rect 295352 539838 295596 539866
rect 296916 539838 297068 539866
rect 297468 539838 297804 539866
rect 298204 539838 298540 539866
rect 298940 539838 299276 539866
rect 299676 539838 300012 539866
rect 300412 539838 300748 539866
rect 301148 539838 301484 539866
rect 301884 539838 302220 539866
rect 302620 539838 302956 539866
rect 303678 539852 303706 540110
rect 304092 539866 304120 543322
rect 305012 539866 305040 543351
rect 305550 543008 305606 543017
rect 305550 542943 305606 542952
rect 305564 539866 305592 542943
rect 306300 540326 306328 598538
rect 306392 545086 306420 599082
rect 306472 598120 306524 598126
rect 306472 598062 306524 598068
rect 306484 576162 306512 598062
rect 306852 591394 306880 600086
rect 307404 598126 307432 600086
rect 308278 599842 308306 600100
rect 308416 600086 308844 600114
rect 309244 600086 309396 600114
rect 309612 600086 309948 600114
rect 310164 600086 310500 600114
rect 310624 600086 311052 600114
rect 311176 600086 311604 600114
rect 312004 600086 312156 600114
rect 312372 600086 312708 600114
rect 308278 599814 308352 599842
rect 307392 598120 307444 598126
rect 307392 598062 307444 598068
rect 308324 597990 308352 599814
rect 308312 597984 308364 597990
rect 308312 597926 308364 597932
rect 307022 597680 307078 597689
rect 307022 597615 307078 597624
rect 307036 594182 307064 597615
rect 307024 594176 307076 594182
rect 307024 594118 307076 594124
rect 306840 591388 306892 591394
rect 306840 591330 306892 591336
rect 308416 586514 308444 600086
rect 309140 598120 309192 598126
rect 309140 598062 309192 598068
rect 307772 586486 308444 586514
rect 306472 576156 306524 576162
rect 306472 576098 306524 576104
rect 307772 567934 307800 586486
rect 307760 567928 307812 567934
rect 307760 567870 307812 567876
rect 306380 545080 306432 545086
rect 306380 545022 306432 545028
rect 309152 544406 309180 598062
rect 309244 552702 309272 600086
rect 309612 586514 309640 600086
rect 310164 598126 310192 600086
rect 310624 598210 310652 600086
rect 310532 598182 310652 598210
rect 310152 598120 310204 598126
rect 310152 598062 310204 598068
rect 309336 586486 309640 586514
rect 309336 556753 309364 586486
rect 310532 570722 310560 598182
rect 311176 586514 311204 600086
rect 311256 598868 311308 598874
rect 311256 598810 311308 598816
rect 311268 598058 311296 598810
rect 311900 598120 311952 598126
rect 311900 598062 311952 598068
rect 311256 598052 311308 598058
rect 311256 597994 311308 598000
rect 310624 586486 311204 586514
rect 310624 584458 310652 586486
rect 310612 584452 310664 584458
rect 310612 584394 310664 584400
rect 310520 570716 310572 570722
rect 310520 570658 310572 570664
rect 311912 561241 311940 598062
rect 312004 592754 312032 600086
rect 312372 598126 312400 600086
rect 313246 599842 313274 600100
rect 313200 599814 313274 599842
rect 313384 600086 313812 600114
rect 314028 600086 314364 600114
rect 312360 598120 312412 598126
rect 312360 598062 312412 598068
rect 313200 596970 313228 599814
rect 313280 598120 313332 598126
rect 313280 598062 313332 598068
rect 313188 596964 313240 596970
rect 313188 596906 313240 596912
rect 311992 592748 312044 592754
rect 311992 592690 312044 592696
rect 311898 561232 311954 561241
rect 311898 561167 311954 561176
rect 309322 556744 309378 556753
rect 309322 556679 309378 556688
rect 309232 552696 309284 552702
rect 309232 552638 309284 552644
rect 312912 545828 312964 545834
rect 312912 545770 312964 545776
rect 309140 544400 309192 544406
rect 309140 544342 309192 544348
rect 306378 543688 306434 543697
rect 306378 543623 306434 543632
rect 306288 540320 306340 540326
rect 306288 540262 306340 540268
rect 306392 539866 306420 543623
rect 307022 543552 307078 543561
rect 307022 543487 307078 543496
rect 307036 539866 307064 543487
rect 312266 543144 312322 543153
rect 312266 543079 312322 543088
rect 308402 542600 308458 542609
rect 308402 542535 308458 542544
rect 309966 542600 310022 542609
rect 309966 542535 310022 542544
rect 311438 542600 311494 542609
rect 311438 542535 311494 542544
rect 308416 539866 308444 542535
rect 308678 542464 308734 542473
rect 308678 542399 308734 542408
rect 309414 542464 309470 542473
rect 309414 542399 309470 542408
rect 304092 539838 304428 539866
rect 305012 539838 305164 539866
rect 305564 539838 305900 539866
rect 306392 539838 306636 539866
rect 307036 539838 307372 539866
rect 308108 539838 308444 539866
rect 308692 539730 308720 542399
rect 309428 539866 309456 542399
rect 309980 539866 310008 542535
rect 311070 542464 311126 542473
rect 311070 542399 311126 542408
rect 311084 540138 311112 542399
rect 311038 540110 311112 540138
rect 309428 539838 309580 539866
rect 309980 539838 310316 539866
rect 311038 539852 311066 540110
rect 311452 539866 311480 542535
rect 312280 539866 312308 543079
rect 312924 539866 312952 545770
rect 313292 541686 313320 598062
rect 313384 566506 313412 600086
rect 314028 598126 314056 600086
rect 314902 599842 314930 600100
rect 314856 599814 314930 599842
rect 315132 600086 315468 600114
rect 315684 600086 316020 600114
rect 316144 600086 316572 600114
rect 316788 600086 317124 600114
rect 317432 600086 317676 600114
rect 314016 598120 314068 598126
rect 314016 598062 314068 598068
rect 314660 598120 314712 598126
rect 314660 598062 314712 598068
rect 313372 566500 313424 566506
rect 313372 566442 313424 566448
rect 314672 554062 314700 598062
rect 314752 598052 314804 598058
rect 314752 597994 314804 598000
rect 314764 573374 314792 597994
rect 314856 588674 314884 599814
rect 315132 598126 315160 600086
rect 315120 598120 315172 598126
rect 315120 598062 315172 598068
rect 315684 598058 315712 600086
rect 316144 598210 316172 600086
rect 316052 598182 316172 598210
rect 315672 598052 315724 598058
rect 315672 597994 315724 598000
rect 314844 588668 314896 588674
rect 314844 588610 314896 588616
rect 314752 573368 314804 573374
rect 314752 573310 314804 573316
rect 314660 554056 314712 554062
rect 314660 553998 314712 554004
rect 313648 545760 313700 545766
rect 313648 545702 313700 545708
rect 313280 541680 313332 541686
rect 313280 541622 313332 541628
rect 313660 539866 313688 545702
rect 315120 543244 315172 543250
rect 315120 543186 315172 543192
rect 314844 543040 314896 543046
rect 314844 542982 314896 542988
rect 311452 539838 311788 539866
rect 312280 539838 312524 539866
rect 312924 539838 313260 539866
rect 313660 539838 313996 539866
rect 308692 539702 308844 539730
rect 291622 539566 291916 539594
rect 292652 539566 292804 539594
rect 293038 539608 293094 539617
rect 291566 539543 291622 539552
rect 294510 539608 294566 539617
rect 293094 539566 293388 539594
rect 293038 539543 293094 539552
rect 295982 539608 296038 539617
rect 294566 539566 294860 539594
rect 294510 539543 294566 539552
rect 314856 539594 314884 542982
rect 315132 539866 315160 543186
rect 316052 543046 316080 598182
rect 316788 586514 316816 600086
rect 316144 586486 316816 586514
rect 316144 559570 316172 586486
rect 316132 559564 316184 559570
rect 316132 559506 316184 559512
rect 317432 545766 317460 600086
rect 319456 580310 319484 639254
rect 319444 580304 319496 580310
rect 319444 580246 319496 580252
rect 319548 572014 319576 641990
rect 321008 641980 321060 641986
rect 321008 641922 321060 641928
rect 320824 640348 320876 640354
rect 320824 640290 320876 640296
rect 320180 599616 320232 599622
rect 320180 599558 320232 599564
rect 320192 596154 320220 599558
rect 320180 596148 320232 596154
rect 320180 596090 320232 596096
rect 319536 572008 319588 572014
rect 319536 571950 319588 571956
rect 317420 545760 317472 545766
rect 317420 545702 317472 545708
rect 317510 543688 317566 543697
rect 317510 543623 317566 543632
rect 316316 543312 316368 543318
rect 316316 543254 316368 543260
rect 316040 543040 316092 543046
rect 316040 542982 316092 542988
rect 315132 539838 315468 539866
rect 316328 539594 316356 543254
rect 316592 543176 316644 543182
rect 316592 543118 316644 543124
rect 316604 539866 316632 543118
rect 316604 539838 316940 539866
rect 296038 539566 296332 539594
rect 314732 539566 314884 539594
rect 316204 539566 316356 539594
rect 317524 539594 317552 543623
rect 317524 539566 317676 539594
rect 295982 539543 296038 539552
rect 284208 539514 284260 539520
rect 320192 537538 320220 596090
rect 320180 537532 320232 537538
rect 320180 537474 320232 537480
rect 320192 537373 320220 537474
rect 320178 537364 320234 537373
rect 320178 537299 320234 537308
rect 281000 528526 281488 528554
rect 281000 281178 281028 528526
rect 320088 511896 320140 511902
rect 320088 511838 320140 511844
rect 320100 510853 320128 511838
rect 320086 510844 320142 510853
rect 320086 510779 320142 510788
rect 320100 510678 320128 510779
rect 319076 510672 319128 510678
rect 319076 510614 319128 510620
rect 320088 510672 320140 510678
rect 320088 510614 320140 510620
rect 318892 508292 318944 508298
rect 318892 508234 318944 508240
rect 318904 508178 318932 508234
rect 318812 508150 318932 508178
rect 295248 500404 295300 500410
rect 295248 500346 295300 500352
rect 281552 500126 282348 500154
rect 281552 369170 281580 500126
rect 283070 499882 283098 500140
rect 283208 500126 283820 500154
rect 284404 500126 284556 500154
rect 284956 500126 285292 500154
rect 283070 499854 283144 499882
rect 282184 418192 282236 418198
rect 282184 418134 282236 418140
rect 281540 369164 281592 369170
rect 281540 369106 281592 369112
rect 282196 287054 282224 418134
rect 282276 365764 282328 365770
rect 282276 365706 282328 365712
rect 282288 318782 282316 365706
rect 282920 338836 282972 338842
rect 282920 338778 282972 338784
rect 282276 318776 282328 318782
rect 282276 318718 282328 318724
rect 282196 287026 282316 287054
rect 282182 281480 282238 281489
rect 282182 281415 282238 281424
rect 280988 281172 281040 281178
rect 280988 281114 281040 281120
rect 280804 281104 280856 281110
rect 280804 281046 280856 281052
rect 282196 280945 282224 281415
rect 282182 280936 282238 280945
rect 282182 280871 282238 280880
rect 279608 280016 279660 280022
rect 279608 279958 279660 279964
rect 282288 279002 282316 287026
rect 282276 278996 282328 279002
rect 282276 278938 282328 278944
rect 282184 202904 282236 202910
rect 282184 202846 282236 202852
rect 279516 125588 279568 125594
rect 279516 125530 279568 125536
rect 282196 88330 282224 202846
rect 282184 88324 282236 88330
rect 282184 88266 282236 88272
rect 279424 71732 279476 71738
rect 279424 71674 279476 71680
rect 282932 16574 282960 338778
rect 283116 333266 283144 499854
rect 283104 333260 283156 333266
rect 283104 333202 283156 333208
rect 283208 225690 283236 500126
rect 284300 494760 284352 494766
rect 284300 494702 284352 494708
rect 283564 369164 283616 369170
rect 283564 369106 283616 369112
rect 283576 324290 283604 369106
rect 283564 324284 283616 324290
rect 283564 324226 283616 324232
rect 284312 292534 284340 494702
rect 284404 344350 284432 500126
rect 284956 494766 284984 500126
rect 286014 499882 286042 500140
rect 286152 500126 286764 500154
rect 287164 500126 287500 500154
rect 287900 500126 288236 500154
rect 288544 500126 288972 500154
rect 289372 500126 289708 500154
rect 289924 500126 290444 500154
rect 290844 500126 291180 500154
rect 291304 500126 291916 500154
rect 286014 499854 286088 499882
rect 286060 497758 286088 499854
rect 286048 497752 286100 497758
rect 286048 497694 286100 497700
rect 285680 496120 285732 496126
rect 285680 496062 285732 496068
rect 284944 494760 284996 494766
rect 284944 494702 284996 494708
rect 284392 344344 284444 344350
rect 284392 344286 284444 344292
rect 285036 331832 285088 331838
rect 285036 331774 285088 331780
rect 284944 329928 284996 329934
rect 284944 329870 284996 329876
rect 284956 317422 284984 329870
rect 285048 325650 285076 331774
rect 285036 325644 285088 325650
rect 285036 325586 285088 325592
rect 284944 317416 284996 317422
rect 284944 317358 284996 317364
rect 284944 295384 284996 295390
rect 284944 295326 284996 295332
rect 284300 292528 284352 292534
rect 284300 292470 284352 292476
rect 284956 281314 284984 295326
rect 284944 281308 284996 281314
rect 284944 281250 284996 281256
rect 283196 225684 283248 225690
rect 283196 225626 283248 225632
rect 284944 205692 284996 205698
rect 284944 205634 284996 205640
rect 284956 91798 284984 205634
rect 284944 91792 284996 91798
rect 284944 91734 284996 91740
rect 285692 16574 285720 496062
rect 286152 489914 286180 500126
rect 287060 494760 287112 494766
rect 287060 494702 287112 494708
rect 285784 489886 286180 489914
rect 285784 340202 285812 489886
rect 285772 340196 285824 340202
rect 285772 340138 285824 340144
rect 287072 278322 287100 494702
rect 287164 349858 287192 500126
rect 287900 494766 287928 500126
rect 287888 494760 287940 494766
rect 287888 494702 287940 494708
rect 288440 491564 288492 491570
rect 288440 491506 288492 491512
rect 287152 349852 287204 349858
rect 287152 349794 287204 349800
rect 287704 342304 287756 342310
rect 287704 342246 287756 342252
rect 287334 280800 287390 280809
rect 287334 280735 287336 280744
rect 287388 280735 287390 280744
rect 287336 280706 287388 280712
rect 287716 278934 287744 342246
rect 288452 337414 288480 491506
rect 288544 354006 288572 500126
rect 289372 491570 289400 500126
rect 289820 494760 289872 494766
rect 289820 494702 289872 494708
rect 289360 491564 289412 491570
rect 289360 491506 289412 491512
rect 289084 452668 289136 452674
rect 289084 452610 289136 452616
rect 288532 354000 288584 354006
rect 288532 353942 288584 353948
rect 288440 337408 288492 337414
rect 288440 337350 288492 337356
rect 287796 331492 287848 331498
rect 287796 331434 287848 331440
rect 287808 320142 287836 331434
rect 287796 320136 287848 320142
rect 287796 320078 287848 320084
rect 287704 278928 287756 278934
rect 287704 278870 287756 278876
rect 287060 278316 287112 278322
rect 287060 278258 287112 278264
rect 287704 207052 287756 207058
rect 287704 206994 287756 207000
rect 287716 93838 287744 206994
rect 289096 117298 289124 452610
rect 289176 382288 289228 382294
rect 289176 382230 289228 382236
rect 289188 285666 289216 382230
rect 289268 353320 289320 353326
rect 289268 353262 289320 353268
rect 289176 285660 289228 285666
rect 289176 285602 289228 285608
rect 289280 279070 289308 353262
rect 289832 341562 289860 494702
rect 289924 482322 289952 500126
rect 290844 494766 290872 500126
rect 290832 494760 290884 494766
rect 290832 494702 290884 494708
rect 289912 482316 289964 482322
rect 289912 482258 289964 482264
rect 289820 341556 289872 341562
rect 289820 341498 289872 341504
rect 289820 337476 289872 337482
rect 289820 337418 289872 337424
rect 289268 279064 289320 279070
rect 289268 279006 289320 279012
rect 289084 117292 289136 117298
rect 289084 117234 289136 117240
rect 287704 93832 287756 93838
rect 287704 93774 287756 93780
rect 278792 16546 279096 16574
rect 282932 16546 283144 16574
rect 285692 16546 286640 16574
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 283116 480 283144 16546
rect 286612 480 286640 16546
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 337418
rect 291304 334694 291332 500126
rect 292638 499882 292666 500140
rect 292776 500126 293388 500154
rect 292638 499854 292712 499882
rect 291936 497820 291988 497826
rect 291936 497762 291988 497768
rect 291844 434784 291896 434790
rect 291844 434726 291896 434732
rect 291292 334688 291344 334694
rect 291292 334630 291344 334636
rect 291856 88330 291884 434726
rect 291948 220250 291976 497762
rect 292028 497752 292080 497758
rect 292028 497694 292080 497700
rect 292040 288386 292068 497694
rect 292580 494760 292632 494766
rect 292580 494702 292632 494708
rect 292028 288380 292080 288386
rect 292028 288322 292080 288328
rect 291936 220244 291988 220250
rect 291936 220186 291988 220192
rect 291844 88324 291896 88330
rect 291844 88266 291896 88272
rect 292592 16574 292620 494702
rect 292684 278526 292712 499854
rect 292776 313274 292804 500126
rect 294110 499882 294138 500140
rect 294248 500126 294860 500154
rect 294110 499854 294184 499882
rect 293224 497752 293276 497758
rect 293224 497694 293276 497700
rect 292764 313268 292816 313274
rect 292764 313210 292816 313216
rect 292672 278520 292724 278526
rect 292672 278462 292724 278468
rect 293236 220182 293264 497694
rect 294156 496398 294184 499854
rect 294144 496392 294196 496398
rect 294144 496334 294196 496340
rect 294248 489914 294276 500126
rect 293972 489886 294276 489914
rect 293316 306400 293368 306406
rect 293316 306342 293368 306348
rect 293328 278798 293356 306342
rect 293972 303618 294000 489886
rect 294604 332240 294656 332246
rect 294604 332182 294656 332188
rect 293960 303612 294012 303618
rect 293960 303554 294012 303560
rect 293316 278792 293368 278798
rect 293316 278734 293368 278740
rect 293224 220176 293276 220182
rect 293224 220118 293276 220124
rect 294616 218754 294644 332182
rect 294972 331968 295024 331974
rect 294972 331910 295024 331916
rect 294880 331628 294932 331634
rect 294880 331570 294932 331576
rect 294696 300892 294748 300898
rect 294696 300834 294748 300840
rect 294708 278866 294736 300834
rect 294892 279478 294920 331570
rect 294880 279472 294932 279478
rect 294880 279414 294932 279420
rect 294696 278860 294748 278866
rect 294696 278802 294748 278808
rect 294984 278254 295012 331910
rect 295064 331900 295116 331906
rect 295064 331842 295116 331848
rect 294972 278248 295024 278254
rect 294972 278190 295024 278196
rect 295076 277982 295104 331842
rect 295156 331288 295208 331294
rect 295156 331230 295208 331236
rect 295064 277976 295116 277982
rect 295064 277918 295116 277924
rect 295168 222970 295196 331230
rect 295156 222964 295208 222970
rect 295156 222906 295208 222912
rect 294604 218748 294656 218754
rect 294604 218690 294656 218696
rect 295260 60314 295288 500346
rect 296628 500268 296680 500274
rect 296628 500210 296680 500216
rect 295352 500126 295596 500154
rect 295812 500126 296332 500154
rect 295352 278594 295380 500126
rect 295812 489914 295840 500126
rect 296536 497956 296588 497962
rect 296536 497898 296588 497904
rect 295984 496392 296036 496398
rect 295984 496334 296036 496340
rect 295444 489886 295840 489914
rect 295444 289474 295472 489886
rect 295432 289468 295484 289474
rect 295432 289410 295484 289416
rect 295996 278730 296024 496334
rect 296260 332104 296312 332110
rect 296260 332046 296312 332052
rect 296074 331392 296130 331401
rect 296074 331327 296130 331336
rect 295984 278724 296036 278730
rect 295984 278666 296036 278672
rect 295340 278588 295392 278594
rect 295340 278530 295392 278536
rect 296088 225622 296116 331327
rect 296168 288448 296220 288454
rect 296168 288390 296220 288396
rect 296180 280022 296208 288390
rect 296168 280016 296220 280022
rect 296168 279958 296220 279964
rect 296272 278458 296300 332046
rect 296352 331764 296404 331770
rect 296352 331706 296404 331712
rect 296260 278452 296312 278458
rect 296260 278394 296312 278400
rect 296076 225616 296128 225622
rect 296076 225558 296128 225564
rect 296364 223106 296392 331706
rect 296444 331560 296496 331566
rect 296444 331502 296496 331508
rect 296352 223100 296404 223106
rect 296352 223042 296404 223048
rect 296456 222902 296484 331502
rect 296548 278662 296576 497898
rect 296536 278656 296588 278662
rect 296536 278598 296588 278604
rect 296444 222896 296496 222902
rect 296444 222838 296496 222844
rect 295984 186380 296036 186386
rect 295984 186322 296036 186328
rect 295996 180305 296024 186322
rect 295982 180296 296038 180305
rect 295982 180231 296038 180240
rect 295982 160848 296038 160857
rect 295982 160783 296038 160792
rect 295996 151094 296024 160783
rect 295984 151088 296036 151094
rect 295984 151030 296036 151036
rect 296074 148880 296130 148889
rect 296074 148815 296130 148824
rect 295982 142896 296038 142905
rect 295982 142831 296038 142840
rect 295996 115938 296024 142831
rect 296088 133210 296116 148815
rect 296076 133204 296128 133210
rect 296076 133146 296128 133152
rect 295984 115932 296036 115938
rect 295984 115874 296036 115880
rect 296640 60382 296668 500210
rect 297068 500126 297312 500154
rect 297284 496194 297312 500126
rect 297376 500126 297804 500154
rect 298112 500126 298540 500154
rect 299276 500126 299428 500154
rect 297272 496188 297324 496194
rect 297272 496130 297324 496136
rect 297376 491978 297404 500126
rect 297364 491972 297416 491978
rect 297364 491914 297416 491920
rect 297640 351280 297692 351286
rect 297640 351222 297692 351228
rect 296996 341624 297048 341630
rect 296996 341566 297048 341572
rect 297008 303929 297036 341566
rect 297362 329760 297418 329769
rect 297362 329695 297418 329704
rect 297086 320240 297142 320249
rect 297086 320175 297142 320184
rect 296994 303920 297050 303929
rect 296994 303855 297050 303864
rect 296994 301200 297050 301209
rect 296994 301135 297050 301144
rect 296810 208720 296866 208729
rect 296810 208655 296866 208664
rect 296824 208418 296852 208655
rect 296812 208412 296864 208418
rect 296812 208354 296864 208360
rect 296810 205728 296866 205737
rect 296810 205663 296812 205672
rect 296864 205663 296866 205672
rect 296812 205634 296864 205640
rect 296812 186312 296864 186318
rect 296810 186280 296812 186289
rect 296864 186280 296866 186289
rect 296810 186215 296866 186224
rect 296810 169824 296866 169833
rect 296810 169759 296812 169768
rect 296864 169759 296866 169768
rect 296812 169730 296864 169736
rect 296810 151872 296866 151881
rect 296810 151807 296812 151816
rect 296864 151807 296866 151816
rect 296812 151778 296864 151784
rect 296812 132456 296864 132462
rect 296810 132424 296812 132433
rect 296864 132424 296866 132433
rect 296810 132359 296866 132368
rect 296812 129736 296864 129742
rect 296812 129678 296864 129684
rect 296824 129441 296852 129678
rect 296810 129432 296866 129441
rect 296810 129367 296866 129376
rect 296812 114504 296864 114510
rect 296810 114472 296812 114481
rect 296864 114472 296866 114481
rect 296810 114407 296866 114416
rect 297008 102513 297036 301135
rect 296994 102504 297050 102513
rect 296994 102439 297050 102448
rect 297100 92041 297128 320175
rect 297178 318880 297234 318889
rect 297178 318815 297234 318824
rect 297192 275398 297220 318815
rect 297272 307760 297324 307766
rect 297272 307702 297324 307708
rect 297284 306649 297312 307702
rect 297270 306640 297326 306649
rect 297270 306575 297326 306584
rect 297376 278050 297404 329695
rect 297454 328400 297510 328409
rect 297454 328335 297510 328344
rect 297364 278044 297416 278050
rect 297364 277986 297416 277992
rect 297468 276826 297496 328335
rect 297546 326360 297602 326369
rect 297546 326295 297602 326304
rect 297456 276820 297508 276826
rect 297456 276762 297508 276768
rect 297180 275392 297232 275398
rect 297180 275334 297232 275340
rect 297560 274038 297588 326295
rect 297652 284209 297680 351222
rect 298008 351212 298060 351218
rect 298008 351154 298060 351160
rect 297916 332648 297968 332654
rect 297916 332590 297968 332596
rect 297730 325000 297786 325009
rect 297730 324935 297786 324944
rect 297744 318866 297772 324935
rect 297824 324284 297876 324290
rect 297824 324226 297876 324232
rect 297836 323649 297864 324226
rect 297822 323640 297878 323649
rect 297822 323575 297878 323584
rect 297744 318838 297864 318866
rect 297732 318776 297784 318782
rect 297732 318718 297784 318724
rect 297744 317529 297772 318718
rect 297730 317520 297786 317529
rect 297730 317455 297786 317464
rect 297732 317416 297784 317422
rect 297732 317358 297784 317364
rect 297744 316169 297772 317358
rect 297730 316160 297786 316169
rect 297730 316095 297786 316104
rect 297836 316034 297864 318838
rect 297744 316006 297864 316034
rect 297744 306374 297772 316006
rect 297928 314809 297956 332590
rect 297914 314800 297970 314809
rect 297914 314735 297970 314744
rect 297916 313268 297968 313274
rect 297916 313210 297968 313216
rect 297928 312769 297956 313210
rect 297914 312760 297970 312769
rect 297914 312695 297970 312704
rect 298020 311409 298048 351154
rect 298112 332654 298140 500126
rect 298744 497888 298796 497894
rect 298744 497830 298796 497836
rect 298652 333396 298704 333402
rect 298652 333338 298704 333344
rect 298100 332648 298152 332654
rect 298100 332590 298152 332596
rect 298560 331424 298612 331430
rect 298560 331366 298612 331372
rect 298006 311400 298062 311409
rect 298006 311335 298062 311344
rect 297916 311092 297968 311098
rect 297916 311034 297968 311040
rect 297744 306346 297864 306374
rect 297730 296440 297786 296449
rect 297730 296375 297786 296384
rect 297744 287178 297772 296375
rect 297836 295186 297864 306346
rect 297928 299169 297956 311034
rect 298008 306332 298060 306338
rect 298008 306274 298060 306280
rect 298020 305289 298048 306274
rect 298006 305280 298062 305289
rect 298006 305215 298062 305224
rect 298008 303612 298060 303618
rect 298008 303554 298060 303560
rect 298020 302569 298048 303554
rect 298006 302560 298062 302569
rect 298006 302495 298062 302504
rect 297914 299160 297970 299169
rect 297914 299095 297970 299104
rect 297824 295180 297876 295186
rect 297824 295122 297876 295128
rect 297822 295080 297878 295089
rect 297822 295015 297878 295024
rect 297836 287434 297864 295015
rect 298008 292528 298060 292534
rect 298008 292470 298060 292476
rect 298020 291689 298048 292470
rect 298006 291680 298062 291689
rect 298006 291615 298062 291624
rect 297914 290320 297970 290329
rect 297914 290255 297970 290264
rect 297928 287450 297956 290255
rect 298008 289468 298060 289474
rect 298008 289410 298060 289416
rect 298020 288969 298048 289410
rect 298006 288960 298062 288969
rect 298006 288895 298062 288904
rect 298008 288380 298060 288386
rect 298008 288322 298060 288328
rect 298020 287609 298048 288322
rect 298006 287600 298062 287609
rect 298006 287535 298062 287544
rect 297824 287428 297876 287434
rect 297928 287422 298048 287450
rect 297824 287370 297876 287376
rect 297744 287150 297956 287178
rect 297824 287088 297876 287094
rect 297824 287030 297876 287036
rect 297836 285938 297864 287030
rect 297824 285932 297876 285938
rect 297824 285874 297876 285880
rect 297928 285818 297956 287150
rect 297744 285790 297956 285818
rect 297638 284200 297694 284209
rect 297638 284135 297694 284144
rect 297744 280634 297772 285790
rect 297824 285728 297876 285734
rect 297824 285670 297876 285676
rect 297732 280628 297784 280634
rect 297732 280570 297784 280576
rect 297640 276072 297692 276078
rect 297640 276014 297692 276020
rect 297548 274032 297600 274038
rect 297548 273974 297600 273980
rect 297364 221604 297416 221610
rect 297364 221546 297416 221552
rect 297376 109993 297404 221546
rect 297456 221536 297508 221542
rect 297456 221478 297508 221484
rect 297362 109984 297418 109993
rect 297362 109919 297418 109928
rect 297468 104009 297496 221478
rect 297546 216744 297602 216753
rect 297546 216679 297602 216688
rect 297454 104000 297510 104009
rect 297454 103935 297510 103944
rect 297560 99521 297588 216679
rect 297546 99512 297602 99521
rect 297546 99447 297602 99456
rect 297652 95033 297680 276014
rect 297732 193180 297784 193186
rect 297732 193122 297784 193128
rect 297744 192273 297772 193122
rect 297730 192264 297786 192273
rect 297730 192199 297786 192208
rect 297732 190460 297784 190466
rect 297732 190402 297784 190408
rect 297744 189281 297772 190402
rect 297730 189272 297786 189281
rect 297730 189207 297786 189216
rect 297836 96529 297864 285670
rect 297916 285660 297968 285666
rect 297916 285602 297968 285608
rect 297928 285569 297956 285602
rect 297914 285560 297970 285569
rect 297914 285495 297970 285504
rect 297914 217696 297970 217705
rect 297914 217631 297970 217640
rect 297928 216714 297956 217631
rect 297916 216708 297968 216714
rect 297916 216650 297968 216656
rect 297914 216200 297970 216209
rect 297914 216135 297970 216144
rect 297928 215354 297956 216135
rect 297916 215348 297968 215354
rect 297916 215290 297968 215296
rect 297914 214704 297970 214713
rect 297914 214639 297970 214648
rect 297928 213994 297956 214639
rect 297916 213988 297968 213994
rect 297916 213930 297968 213936
rect 297914 213208 297970 213217
rect 297914 213143 297970 213152
rect 297928 212566 297956 213143
rect 297916 212560 297968 212566
rect 297916 212502 297968 212508
rect 297914 211712 297970 211721
rect 297914 211647 297970 211656
rect 297928 211206 297956 211647
rect 297916 211200 297968 211206
rect 297916 211142 297968 211148
rect 297914 210216 297970 210225
rect 297914 210151 297970 210160
rect 297928 209846 297956 210151
rect 297916 209840 297968 209846
rect 297916 209782 297968 209788
rect 297914 207224 297970 207233
rect 297914 207159 297970 207168
rect 297928 207058 297956 207159
rect 297916 207052 297968 207058
rect 297916 206994 297968 207000
rect 297914 204232 297970 204241
rect 297914 204167 297970 204176
rect 297928 202910 297956 204167
rect 297916 202904 297968 202910
rect 297916 202846 297968 202852
rect 297914 202736 297970 202745
rect 297914 202671 297970 202680
rect 297928 201550 297956 202671
rect 297916 201544 297968 201550
rect 297916 201486 297968 201492
rect 297914 201240 297970 201249
rect 297914 201175 297970 201184
rect 297928 200190 297956 201175
rect 297916 200184 297968 200190
rect 297916 200126 297968 200132
rect 297914 199744 297970 199753
rect 297914 199679 297970 199688
rect 297928 198762 297956 199679
rect 297916 198756 297968 198762
rect 297916 198698 297968 198704
rect 297914 198248 297970 198257
rect 297914 198183 297970 198192
rect 297928 197402 297956 198183
rect 297916 197396 297968 197402
rect 297916 197338 297968 197344
rect 297914 196752 297970 196761
rect 297914 196687 297970 196696
rect 297928 196042 297956 196687
rect 297916 196036 297968 196042
rect 297916 195978 297968 195984
rect 297914 195256 297970 195265
rect 297914 195191 297970 195200
rect 297928 194614 297956 195191
rect 297916 194608 297968 194614
rect 297916 194550 297968 194556
rect 297914 193760 297970 193769
rect 297914 193695 297970 193704
rect 297928 193254 297956 193695
rect 297916 193248 297968 193254
rect 297916 193190 297968 193196
rect 297914 190768 297970 190777
rect 297914 190703 297970 190712
rect 297928 190534 297956 190703
rect 297916 190528 297968 190534
rect 297916 190470 297968 190476
rect 297916 189032 297968 189038
rect 297916 188974 297968 188980
rect 297928 187785 297956 188974
rect 297914 187776 297970 187785
rect 297914 187711 297970 187720
rect 297916 184884 297968 184890
rect 297916 184826 297968 184832
rect 297928 184793 297956 184826
rect 297914 184784 297970 184793
rect 297914 184719 297970 184728
rect 297916 183524 297968 183530
rect 297916 183466 297968 183472
rect 297928 183297 297956 183466
rect 297914 183288 297970 183297
rect 297914 183223 297970 183232
rect 297916 182164 297968 182170
rect 297916 182106 297968 182112
rect 297928 181801 297956 182106
rect 297914 181792 297970 181801
rect 297914 181727 297970 181736
rect 297916 179376 297968 179382
rect 297916 179318 297968 179324
rect 297928 178809 297956 179318
rect 297914 178800 297970 178809
rect 297914 178735 297970 178744
rect 297916 178016 297968 178022
rect 297916 177958 297968 177964
rect 297928 177313 297956 177958
rect 297914 177304 297970 177313
rect 297914 177239 297970 177248
rect 297916 176656 297968 176662
rect 297916 176598 297968 176604
rect 297928 175817 297956 176598
rect 297914 175808 297970 175817
rect 297914 175743 297970 175752
rect 297916 175228 297968 175234
rect 297916 175170 297968 175176
rect 297928 174321 297956 175170
rect 297914 174312 297970 174321
rect 297914 174247 297970 174256
rect 297916 173188 297968 173194
rect 297916 173130 297968 173136
rect 297928 172825 297956 173130
rect 297914 172816 297970 172825
rect 297914 172751 297970 172760
rect 297914 171320 297970 171329
rect 297914 171255 297970 171264
rect 297928 171154 297956 171255
rect 297916 171148 297968 171154
rect 297916 171090 297968 171096
rect 297914 168328 297970 168337
rect 297914 168263 297970 168272
rect 297928 167074 297956 168263
rect 297916 167068 297968 167074
rect 297916 167010 297968 167016
rect 297914 166832 297970 166841
rect 297914 166767 297970 166776
rect 297928 165646 297956 166767
rect 297916 165640 297968 165646
rect 297916 165582 297968 165588
rect 297914 165336 297970 165345
rect 297914 165271 297970 165280
rect 297928 164286 297956 165271
rect 297916 164280 297968 164286
rect 297916 164222 297968 164228
rect 297914 163840 297970 163849
rect 297914 163775 297970 163784
rect 297928 162926 297956 163775
rect 297916 162920 297968 162926
rect 297916 162862 297968 162868
rect 297914 162344 297970 162353
rect 297914 162279 297970 162288
rect 297928 161498 297956 162279
rect 297916 161492 297968 161498
rect 297916 161434 297968 161440
rect 297914 159352 297970 159361
rect 297914 159287 297970 159296
rect 297928 158778 297956 159287
rect 297916 158772 297968 158778
rect 297916 158714 297968 158720
rect 297914 157856 297970 157865
rect 297914 157791 297970 157800
rect 297928 157418 297956 157791
rect 297916 157412 297968 157418
rect 297916 157354 297968 157360
rect 297914 156360 297970 156369
rect 297914 156295 297970 156304
rect 297928 155990 297956 156295
rect 297916 155984 297968 155990
rect 297916 155926 297968 155932
rect 297914 154864 297970 154873
rect 297914 154799 297970 154808
rect 297928 154630 297956 154799
rect 297916 154624 297968 154630
rect 297916 154566 297968 154572
rect 297914 153368 297970 153377
rect 297914 153303 297970 153312
rect 297928 153270 297956 153303
rect 297916 153264 297968 153270
rect 297916 153206 297968 153212
rect 297914 150376 297970 150385
rect 297914 150311 297970 150320
rect 297928 149122 297956 150311
rect 297916 149116 297968 149122
rect 297916 149058 297968 149064
rect 297914 147384 297970 147393
rect 297914 147319 297970 147328
rect 297928 146334 297956 147319
rect 297916 146328 297968 146334
rect 297916 146270 297968 146276
rect 297914 145888 297970 145897
rect 297914 145823 297970 145832
rect 297928 144974 297956 145823
rect 297916 144968 297968 144974
rect 297916 144910 297968 144916
rect 297914 144392 297970 144401
rect 297914 144327 297970 144336
rect 297928 143614 297956 144327
rect 297916 143608 297968 143614
rect 297916 143550 297968 143556
rect 297916 142112 297968 142118
rect 297916 142054 297968 142060
rect 297928 141409 297956 142054
rect 297914 141400 297970 141409
rect 297914 141335 297970 141344
rect 297916 140752 297968 140758
rect 297916 140694 297968 140700
rect 297928 139913 297956 140694
rect 297914 139904 297970 139913
rect 297914 139839 297970 139848
rect 297916 139392 297968 139398
rect 297916 139334 297968 139340
rect 297928 138417 297956 139334
rect 297914 138408 297970 138417
rect 297914 138343 297970 138352
rect 297916 137964 297968 137970
rect 297916 137906 297968 137912
rect 297928 136921 297956 137906
rect 297914 136912 297970 136921
rect 297914 136847 297970 136856
rect 297916 136604 297968 136610
rect 297916 136546 297968 136552
rect 297928 135425 297956 136546
rect 297914 135416 297970 135425
rect 297914 135351 297970 135360
rect 297916 135244 297968 135250
rect 297916 135186 297968 135192
rect 297928 133929 297956 135186
rect 297914 133920 297970 133929
rect 297914 133855 297970 133864
rect 297916 131096 297968 131102
rect 297916 131038 297968 131044
rect 297928 130937 297956 131038
rect 297914 130928 297970 130937
rect 297914 130863 297970 130872
rect 297916 128308 297968 128314
rect 297916 128250 297968 128256
rect 297928 127945 297956 128250
rect 297914 127936 297970 127945
rect 297914 127871 297970 127880
rect 297916 126948 297968 126954
rect 297916 126890 297968 126896
rect 297928 126449 297956 126890
rect 297914 126440 297970 126449
rect 297914 126375 297970 126384
rect 297916 125588 297968 125594
rect 297916 125530 297968 125536
rect 297928 124953 297956 125530
rect 297914 124944 297970 124953
rect 297914 124879 297970 124888
rect 297916 124160 297968 124166
rect 297916 124102 297968 124108
rect 297928 123457 297956 124102
rect 297914 123448 297970 123457
rect 297914 123383 297970 123392
rect 297916 122800 297968 122806
rect 297916 122742 297968 122748
rect 297928 121961 297956 122742
rect 297914 121952 297970 121961
rect 297914 121887 297970 121896
rect 297916 121440 297968 121446
rect 297916 121382 297968 121388
rect 297928 120465 297956 121382
rect 297914 120456 297970 120465
rect 297914 120391 297970 120400
rect 297916 120080 297968 120086
rect 297916 120022 297968 120028
rect 297928 118969 297956 120022
rect 297914 118960 297970 118969
rect 297914 118895 297970 118904
rect 297916 118652 297968 118658
rect 297916 118594 297968 118600
rect 297928 117473 297956 118594
rect 297914 117464 297970 117473
rect 297914 117399 297970 117408
rect 297916 117292 297968 117298
rect 297916 117234 297968 117240
rect 297928 115977 297956 117234
rect 297914 115968 297970 115977
rect 297914 115903 297970 115912
rect 297916 113144 297968 113150
rect 297916 113086 297968 113092
rect 297928 112985 297956 113086
rect 297914 112976 297970 112985
rect 297914 112911 297970 112920
rect 297822 96520 297878 96529
rect 297822 96455 297878 96464
rect 297638 95024 297694 95033
rect 297638 94959 297694 94968
rect 297086 92032 297142 92041
rect 297086 91967 297142 91976
rect 298020 90545 298048 287422
rect 298098 282432 298154 282441
rect 298098 282367 298154 282376
rect 298112 282062 298140 282367
rect 298100 282056 298152 282062
rect 298100 281998 298152 282004
rect 298572 279954 298600 331366
rect 298664 281489 298692 333338
rect 298756 311098 298784 497830
rect 299400 495038 299428 500126
rect 299676 500126 300012 500154
rect 300412 500126 300748 500154
rect 300964 500126 301484 500154
rect 301884 500126 302220 500154
rect 302436 500126 302956 500154
rect 299388 495032 299440 495038
rect 299388 494974 299440 494980
rect 299480 494692 299532 494698
rect 299480 494634 299532 494640
rect 299492 336054 299520 494634
rect 299572 454028 299624 454034
rect 299572 453970 299624 453976
rect 299480 336048 299532 336054
rect 299480 335990 299532 335996
rect 298836 332308 298888 332314
rect 298836 332250 298888 332256
rect 298744 311092 298796 311098
rect 298744 311034 298796 311040
rect 298742 308680 298798 308689
rect 298742 308615 298798 308624
rect 298650 281480 298706 281489
rect 298650 281415 298706 281424
rect 298560 279948 298612 279954
rect 298560 279890 298612 279896
rect 298756 278186 298784 308615
rect 298744 278180 298796 278186
rect 298744 278122 298796 278128
rect 298848 276078 298876 332250
rect 299020 330200 299072 330206
rect 299020 330142 299072 330148
rect 298928 329996 298980 330002
rect 298928 329938 298980 329944
rect 298836 276072 298888 276078
rect 298836 276014 298888 276020
rect 298836 220244 298888 220250
rect 298836 220186 298888 220192
rect 298744 220176 298796 220182
rect 298744 220118 298796 220124
rect 298756 98025 298784 220118
rect 298742 98016 298798 98025
rect 298742 97951 298798 97960
rect 298848 93537 298876 220186
rect 298940 111489 298968 329938
rect 298926 111480 298982 111489
rect 298926 111415 298982 111424
rect 299032 108497 299060 330142
rect 299112 330132 299164 330138
rect 299112 330074 299164 330080
rect 299018 108488 299074 108497
rect 299018 108423 299074 108432
rect 299124 107001 299152 330074
rect 299204 330064 299256 330070
rect 299204 330006 299256 330012
rect 299110 106992 299166 107001
rect 299110 106927 299166 106936
rect 299216 105505 299244 330006
rect 299296 329928 299348 329934
rect 299296 329870 299348 329876
rect 299202 105496 299258 105505
rect 299202 105431 299258 105440
rect 299308 101017 299336 329870
rect 299386 311400 299442 311409
rect 299386 311335 299442 311344
rect 299400 281466 299428 311335
rect 299584 297809 299612 453970
rect 299676 345710 299704 500126
rect 300412 494698 300440 500126
rect 300400 494692 300452 494698
rect 300400 494634 300452 494640
rect 300964 454034 300992 500126
rect 301884 497690 301912 500126
rect 301872 497684 301924 497690
rect 301872 497626 301924 497632
rect 302332 495032 302384 495038
rect 302332 494974 302384 494980
rect 300952 454028 301004 454034
rect 300952 453970 301004 453976
rect 301504 371272 301556 371278
rect 301504 371214 301556 371220
rect 299664 345704 299716 345710
rect 299664 345646 299716 345652
rect 301516 332994 301544 371214
rect 301504 332988 301556 332994
rect 301504 332930 301556 332936
rect 299756 332580 299808 332586
rect 299756 332522 299808 332528
rect 299662 322280 299718 322289
rect 299662 322215 299718 322224
rect 299570 297800 299626 297809
rect 299570 297735 299626 297744
rect 299570 282840 299626 282849
rect 299570 282775 299626 282784
rect 299400 281438 299520 281466
rect 299492 222154 299520 281438
rect 299584 271182 299612 282775
rect 299676 276146 299704 322215
rect 299768 278390 299796 332522
rect 300676 331356 300728 331362
rect 300676 331298 300728 331304
rect 300688 329868 300716 331298
rect 301964 331288 302016 331294
rect 301964 331230 302016 331236
rect 301976 329868 302004 331230
rect 302344 330018 302372 494974
rect 302436 331906 302464 500126
rect 303678 499882 303706 500140
rect 303632 499854 303706 499882
rect 303816 500126 304428 500154
rect 303632 331906 303660 499854
rect 303816 332042 303844 500126
rect 305150 499882 305178 500140
rect 305104 499854 305178 499882
rect 305564 500126 305900 500154
rect 306392 500126 306636 500154
rect 306760 500126 307372 500154
rect 307864 500126 308108 500154
rect 308508 500126 308844 500154
rect 309152 500126 309580 500154
rect 309704 500126 310316 500154
rect 310532 500126 311052 500154
rect 311176 500126 311788 500154
rect 312188 500126 312524 500154
rect 312648 500126 313260 500154
rect 313384 500126 313996 500154
rect 303804 332036 303856 332042
rect 303804 331978 303856 331984
rect 305104 331974 305132 499854
rect 305564 497962 305592 500126
rect 305552 497956 305604 497962
rect 305552 497898 305604 497904
rect 306392 332586 306420 500126
rect 306760 489914 306788 500126
rect 307760 494148 307812 494154
rect 307760 494090 307812 494096
rect 306484 489886 306788 489914
rect 306484 333334 306512 489886
rect 307772 333402 307800 494090
rect 307864 487898 307892 500126
rect 308508 494154 308536 500126
rect 308496 494148 308548 494154
rect 308496 494090 308548 494096
rect 307852 487892 307904 487898
rect 307852 487834 307904 487840
rect 307760 333396 307812 333402
rect 307760 333338 307812 333344
rect 306472 333328 306524 333334
rect 306472 333270 306524 333276
rect 306472 332988 306524 332994
rect 306472 332930 306524 332936
rect 306380 332580 306432 332586
rect 306380 332522 306432 332528
rect 305092 331968 305144 331974
rect 305092 331910 305144 331916
rect 302424 331900 302476 331906
rect 302424 331842 302476 331848
rect 303620 331900 303672 331906
rect 303620 331842 303672 331848
rect 305182 331256 305238 331265
rect 305182 331191 305238 331200
rect 302344 329990 302832 330018
rect 302804 329882 302832 329990
rect 302804 329854 303278 329882
rect 305196 329868 305224 331191
rect 306484 329868 306512 332930
rect 309152 331974 309180 500126
rect 309704 489914 309732 500126
rect 309244 489886 309732 489914
rect 309244 332110 309272 489886
rect 310532 334762 310560 500126
rect 311176 489914 311204 500126
rect 312188 497894 312216 500126
rect 312176 497888 312228 497894
rect 312176 497830 312228 497836
rect 311900 496188 311952 496194
rect 311900 496130 311952 496136
rect 310624 489886 311204 489914
rect 310624 338774 310652 489886
rect 310612 338768 310664 338774
rect 310612 338710 310664 338716
rect 310520 334756 310572 334762
rect 310520 334698 310572 334704
rect 310336 332240 310388 332246
rect 310336 332182 310388 332188
rect 309232 332104 309284 332110
rect 309232 332046 309284 332052
rect 309140 331968 309192 331974
rect 309140 331910 309192 331916
rect 309048 331764 309100 331770
rect 309048 331706 309100 331712
rect 307760 331424 307812 331430
rect 307760 331366 307812 331372
rect 307772 329868 307800 331366
rect 309060 329868 309088 331706
rect 310348 329868 310376 332182
rect 311912 329882 311940 496130
rect 312648 489914 312676 500126
rect 312004 489886 312676 489914
rect 312004 341630 312032 489886
rect 313384 351286 313412 500126
rect 314718 499882 314746 500140
rect 314672 499854 314746 499882
rect 315132 500126 315468 500154
rect 316052 500126 316204 500154
rect 316604 500126 316940 500154
rect 317432 500126 317676 500154
rect 314672 497554 314700 499854
rect 315132 497826 315160 500126
rect 315120 497820 315172 497826
rect 315120 497762 315172 497768
rect 316052 497758 316080 500126
rect 316040 497752 316092 497758
rect 316040 497694 316092 497700
rect 316604 497622 316632 500126
rect 316592 497616 316644 497622
rect 316592 497558 316644 497564
rect 314660 497548 314712 497554
rect 314660 497490 314712 497496
rect 317432 497486 317460 500126
rect 317420 497480 317472 497486
rect 317420 497422 317472 497428
rect 317420 389224 317472 389230
rect 317420 389166 317472 389172
rect 313372 351280 313424 351286
rect 313372 351222 313424 351228
rect 314660 345704 314712 345710
rect 314660 345646 314712 345652
rect 311992 341624 312044 341630
rect 311992 341566 312044 341572
rect 313556 331628 313608 331634
rect 313556 331570 313608 331576
rect 311912 329854 312294 329882
rect 313568 329868 313596 331570
rect 314672 329882 314700 345646
rect 317432 345014 317460 389166
rect 317432 344986 317736 345014
rect 316130 331392 316186 331401
rect 316130 331327 316186 331336
rect 314672 329854 314870 329882
rect 316144 329868 316172 331327
rect 317708 329882 317736 344986
rect 318812 338842 318840 508150
rect 318892 506524 318944 506530
rect 318892 506466 318944 506472
rect 318904 340270 318932 506466
rect 318984 506388 319036 506394
rect 318984 506330 319036 506336
rect 318996 487830 319024 506330
rect 319088 494766 319116 510614
rect 319350 508328 319406 508337
rect 319350 508263 319352 508272
rect 319404 508263 319406 508272
rect 319352 508234 319404 508240
rect 319364 507890 319392 508234
rect 319352 507884 319404 507890
rect 319352 507826 319404 507832
rect 319350 506560 319406 506569
rect 319350 506495 319352 506504
rect 319404 506495 319406 506504
rect 319352 506466 319404 506472
rect 320088 506388 320140 506394
rect 320088 506330 320140 506336
rect 320100 506093 320128 506330
rect 320086 506084 320142 506093
rect 320086 506019 320142 506028
rect 319076 494760 319128 494766
rect 319076 494702 319128 494708
rect 318984 487824 319036 487830
rect 318984 487766 319036 487772
rect 320192 351218 320220 537299
rect 320364 510604 320416 510610
rect 320364 510546 320416 510552
rect 320376 509493 320404 510546
rect 320362 509484 320418 509493
rect 320362 509419 320418 509428
rect 320272 508156 320324 508162
rect 320270 508124 320272 508133
rect 320324 508124 320326 508133
rect 320270 508059 320326 508068
rect 320272 507816 320324 507822
rect 320272 507758 320324 507764
rect 320284 507453 320312 507758
rect 320270 507444 320326 507453
rect 320270 507379 320326 507388
rect 320272 506456 320324 506462
rect 320272 506398 320324 506404
rect 320284 505413 320312 506398
rect 320270 505404 320326 505413
rect 320270 505339 320326 505348
rect 320272 503872 320324 503878
rect 320272 503814 320324 503820
rect 320284 486470 320312 503814
rect 320376 496126 320404 509419
rect 320640 508156 320692 508162
rect 320640 508098 320692 508104
rect 320548 507816 320600 507822
rect 320548 507758 320600 507764
rect 320454 505336 320510 505345
rect 320454 505271 320510 505280
rect 320364 496120 320416 496126
rect 320364 496062 320416 496068
rect 320468 493338 320496 505271
rect 320560 503878 320588 507758
rect 320548 503872 320600 503878
rect 320548 503814 320600 503820
rect 320652 498846 320680 508098
rect 320640 498840 320692 498846
rect 320640 498782 320692 498788
rect 320456 493332 320508 493338
rect 320456 493274 320508 493280
rect 320272 486464 320324 486470
rect 320272 486406 320324 486412
rect 320836 365702 320864 640290
rect 320916 598460 320968 598466
rect 320916 598402 320968 598408
rect 320928 498778 320956 598402
rect 321020 560998 321048 641922
rect 321100 641776 321152 641782
rect 321100 641718 321152 641724
rect 321112 562426 321140 641718
rect 321204 577522 321232 642262
rect 322296 642116 322348 642122
rect 322296 642058 322348 642064
rect 322204 639192 322256 639198
rect 322204 639134 322256 639140
rect 321192 577516 321244 577522
rect 321192 577458 321244 577464
rect 321100 562420 321152 562426
rect 321100 562362 321152 562368
rect 321008 560992 321060 560998
rect 321008 560934 321060 560940
rect 322112 535356 322164 535362
rect 322112 535298 322164 535304
rect 322124 534993 322152 535298
rect 322110 534984 322166 534993
rect 322110 534919 322166 534928
rect 321652 532704 321704 532710
rect 321652 532646 321704 532652
rect 321664 532273 321692 532646
rect 321650 532264 321706 532273
rect 321650 532199 321706 532208
rect 322112 528556 322164 528562
rect 322112 528498 322164 528504
rect 322124 528193 322152 528498
rect 322110 528184 322166 528193
rect 322110 528119 322166 528128
rect 322216 527134 322244 639134
rect 322308 554130 322336 642058
rect 322388 640416 322440 640422
rect 322388 640358 322440 640364
rect 322400 578202 322428 640358
rect 324964 639328 325016 639334
rect 324964 639270 325016 639276
rect 323676 598188 323728 598194
rect 323676 598130 323728 598136
rect 323584 597984 323636 597990
rect 323584 597926 323636 597932
rect 322480 592748 322532 592754
rect 322480 592690 322532 592696
rect 322388 578196 322440 578202
rect 322388 578138 322440 578144
rect 322296 554124 322348 554130
rect 322296 554066 322348 554072
rect 322388 551608 322440 551614
rect 322388 551550 322440 551556
rect 322296 548616 322348 548622
rect 322296 548558 322348 548564
rect 322204 527128 322256 527134
rect 322204 527070 322256 527076
rect 322308 525745 322336 548558
rect 322294 525736 322350 525745
rect 322294 525671 322350 525680
rect 322110 524648 322166 524657
rect 322110 524583 322166 524592
rect 322124 521966 322152 524583
rect 322294 524512 322350 524521
rect 322294 524447 322350 524456
rect 322202 522336 322258 522345
rect 322202 522271 322258 522280
rect 322112 521960 322164 521966
rect 322112 521902 322164 521908
rect 322216 520946 322244 522271
rect 322204 520940 322256 520946
rect 322204 520882 322256 520888
rect 322204 520804 322256 520810
rect 322204 520746 322256 520752
rect 322018 520704 322074 520713
rect 322018 520639 322074 520648
rect 322032 520334 322060 520639
rect 322216 520350 322244 520746
rect 322308 520418 322336 524447
rect 322400 520810 322428 551550
rect 322492 546446 322520 592690
rect 322480 546440 322532 546446
rect 322480 546382 322532 546388
rect 322940 537600 322992 537606
rect 322940 537542 322992 537548
rect 322570 536208 322626 536217
rect 322570 536143 322626 536152
rect 322478 535256 322534 535265
rect 322478 535191 322480 535200
rect 322532 535191 322534 535200
rect 322480 535162 322532 535168
rect 322584 534750 322612 536143
rect 322572 534744 322624 534750
rect 322572 534686 322624 534692
rect 322846 534032 322902 534041
rect 322952 534018 322980 537542
rect 322902 533990 322980 534018
rect 322846 533967 322902 533976
rect 322480 533452 322532 533458
rect 322480 533394 322532 533400
rect 322492 533361 322520 533394
rect 322848 533384 322900 533390
rect 322478 533352 322534 533361
rect 322848 533326 322900 533332
rect 322478 533287 322534 533296
rect 322754 532400 322810 532409
rect 322754 532335 322810 532344
rect 322478 531312 322534 531321
rect 322478 531247 322480 531256
rect 322532 531247 322534 531256
rect 322480 531218 322532 531224
rect 322664 530596 322716 530602
rect 322664 530538 322716 530544
rect 322570 530224 322626 530233
rect 322570 530159 322626 530168
rect 322584 529990 322612 530159
rect 322572 529984 322624 529990
rect 322572 529926 322624 529932
rect 322480 529916 322532 529922
rect 322480 529858 322532 529864
rect 322492 529825 322520 529858
rect 322478 529816 322534 529825
rect 322478 529751 322534 529760
rect 322480 529712 322532 529718
rect 322480 529654 322532 529660
rect 322492 528465 322520 529654
rect 322676 529530 322704 530538
rect 322584 529502 322704 529530
rect 322478 528456 322534 528465
rect 322478 528391 322534 528400
rect 322584 527202 322612 529502
rect 322768 528554 322796 532335
rect 322860 529718 322888 533326
rect 322848 529712 322900 529718
rect 322848 529654 322900 529660
rect 322846 528864 322902 528873
rect 322846 528799 322902 528808
rect 322676 528526 322796 528554
rect 322572 527196 322624 527202
rect 322572 527138 322624 527144
rect 322570 527096 322626 527105
rect 322480 527060 322532 527066
rect 322570 527031 322626 527040
rect 322480 527002 322532 527008
rect 322492 526833 322520 527002
rect 322584 526998 322612 527031
rect 322572 526992 322624 526998
rect 322572 526934 322624 526940
rect 322478 526824 322534 526833
rect 322478 526759 322534 526768
rect 322676 523734 322704 528526
rect 322756 527196 322808 527202
rect 322756 527138 322808 527144
rect 322664 523728 322716 523734
rect 322664 523670 322716 523676
rect 322662 523288 322718 523297
rect 322662 523223 322718 523232
rect 322478 523152 322534 523161
rect 322478 523087 322534 523096
rect 322492 522306 322520 523087
rect 322572 522980 322624 522986
rect 322572 522922 322624 522928
rect 322480 522300 322532 522306
rect 322480 522242 322532 522248
rect 322584 522209 322612 522922
rect 322570 522200 322626 522209
rect 322570 522135 322626 522144
rect 322676 522050 322704 523223
rect 322584 522022 322704 522050
rect 322480 521620 322532 521626
rect 322480 521562 322532 521568
rect 322388 520804 322440 520810
rect 322388 520746 322440 520752
rect 322492 520577 322520 521562
rect 322478 520568 322534 520577
rect 322478 520503 322534 520512
rect 322308 520390 322520 520418
rect 322020 520328 322072 520334
rect 322216 520322 322428 520350
rect 322020 520270 322072 520276
rect 321652 520260 321704 520266
rect 321652 520202 321704 520208
rect 321664 519489 321692 520202
rect 322202 519616 322258 519625
rect 322202 519551 322258 519560
rect 321650 519480 321706 519489
rect 321650 519415 321706 519424
rect 322216 519314 322244 519551
rect 322204 519308 322256 519314
rect 322204 519250 322256 519256
rect 321744 518084 321796 518090
rect 321744 518026 321796 518032
rect 321756 517857 321784 518026
rect 322294 517984 322350 517993
rect 322294 517919 322350 517928
rect 321742 517848 321798 517857
rect 321742 517783 321798 517792
rect 322308 517614 322336 517919
rect 322296 517608 322348 517614
rect 322296 517550 322348 517556
rect 322296 516112 322348 516118
rect 322296 516054 322348 516060
rect 322308 515409 322336 516054
rect 322294 515400 322350 515409
rect 322294 515335 322350 515344
rect 322294 513496 322350 513505
rect 322294 513431 322296 513440
rect 322348 513431 322350 513440
rect 322296 513402 322348 513408
rect 321742 512680 321798 512689
rect 321742 512615 321798 512624
rect 322202 512680 322258 512689
rect 322202 512615 322204 512624
rect 321558 511320 321614 511329
rect 321558 511255 321560 511264
rect 321612 511255 321614 511264
rect 321560 511226 321612 511232
rect 321572 506070 321600 511226
rect 321650 509688 321706 509697
rect 321650 509623 321706 509632
rect 321664 508638 321692 509623
rect 321652 508632 321704 508638
rect 321652 508574 321704 508580
rect 321572 506042 321692 506070
rect 321558 504656 321614 504665
rect 321558 504591 321614 504600
rect 321572 503742 321600 504591
rect 321560 503736 321612 503742
rect 321560 503678 321612 503684
rect 320916 498772 320968 498778
rect 320916 498714 320968 498720
rect 320824 365696 320876 365702
rect 320824 365638 320876 365644
rect 320180 351212 320232 351218
rect 320180 351154 320232 351160
rect 318892 340264 318944 340270
rect 318892 340206 318944 340212
rect 318800 338836 318852 338842
rect 318800 338778 318852 338784
rect 319352 336048 319404 336054
rect 319352 335990 319404 335996
rect 317708 329854 318090 329882
rect 319364 329868 319392 335990
rect 321572 334626 321600 503678
rect 321664 349761 321692 506042
rect 321756 500274 321784 512615
rect 322256 512615 322258 512624
rect 322204 512586 322256 512592
rect 322202 512136 322258 512145
rect 322202 512071 322258 512080
rect 322216 511970 322244 512071
rect 322204 511964 322256 511970
rect 322204 511906 322256 511912
rect 321744 500268 321796 500274
rect 321744 500210 321796 500216
rect 321650 349752 321706 349761
rect 321650 349687 321706 349696
rect 322216 336025 322244 511906
rect 322296 509244 322348 509250
rect 322296 509186 322348 509192
rect 322308 508638 322336 509186
rect 322296 508632 322348 508638
rect 322296 508574 322348 508580
rect 322308 337482 322336 508574
rect 322400 506841 322428 520322
rect 322386 506832 322442 506841
rect 322386 506767 322442 506776
rect 322492 505186 322520 520390
rect 322584 505306 322612 522022
rect 322664 521960 322716 521966
rect 322664 521902 322716 521908
rect 322572 505300 322624 505306
rect 322572 505242 322624 505248
rect 322492 505158 322612 505186
rect 322480 505096 322532 505102
rect 322480 505038 322532 505044
rect 322492 504529 322520 505038
rect 322478 504520 322534 504529
rect 322478 504455 322534 504464
rect 322480 503668 322532 503674
rect 322480 503610 322532 503616
rect 322492 503577 322520 503610
rect 322478 503568 322534 503577
rect 322478 503503 322534 503512
rect 322478 502480 322534 502489
rect 322478 502415 322534 502424
rect 322492 500342 322520 502415
rect 322584 500954 322612 505158
rect 322676 502994 322704 521902
rect 322768 517449 322796 527138
rect 322860 525094 322888 528799
rect 322848 525088 322900 525094
rect 322848 525030 322900 525036
rect 322848 517472 322900 517478
rect 322754 517440 322810 517449
rect 322848 517414 322900 517420
rect 322754 517375 322810 517384
rect 322860 516769 322888 517414
rect 322846 516760 322902 516769
rect 322846 516695 322902 516704
rect 322846 515536 322902 515545
rect 322846 515471 322902 515480
rect 322860 515438 322888 515471
rect 322848 515432 322900 515438
rect 322848 515374 322900 515380
rect 322754 514176 322810 514185
rect 322754 514111 322810 514120
rect 322768 514078 322796 514111
rect 322756 514072 322808 514078
rect 322756 514014 322808 514020
rect 322940 514072 322992 514078
rect 322940 514014 322992 514020
rect 322756 505300 322808 505306
rect 322756 505242 322808 505248
rect 322664 502988 322716 502994
rect 322664 502930 322716 502936
rect 322572 500948 322624 500954
rect 322572 500890 322624 500896
rect 322480 500336 322532 500342
rect 322480 500278 322532 500284
rect 322768 500274 322796 505242
rect 322952 500410 322980 514014
rect 322940 500404 322992 500410
rect 322940 500346 322992 500352
rect 322756 500268 322808 500274
rect 322756 500210 322808 500216
rect 323596 499322 323624 597926
rect 323688 499390 323716 598130
rect 324228 549432 324280 549438
rect 324228 549374 324280 549380
rect 324240 518945 324268 549374
rect 324226 518936 324282 518945
rect 324226 518871 324282 518880
rect 324240 518090 324268 518871
rect 324228 518084 324280 518090
rect 324228 518026 324280 518032
rect 324320 517676 324372 517682
rect 324320 517618 324372 517624
rect 324332 517478 324360 517618
rect 324320 517472 324372 517478
rect 324320 517414 324372 517420
rect 324228 515432 324280 515438
rect 324228 515374 324280 515380
rect 324240 509930 324268 515374
rect 324228 509924 324280 509930
rect 324228 509866 324280 509872
rect 323676 499384 323728 499390
rect 323676 499326 323728 499332
rect 323584 499316 323636 499322
rect 323584 499258 323636 499264
rect 323584 423700 323636 423706
rect 323584 423642 323636 423648
rect 322296 337476 322348 337482
rect 322296 337418 322348 337424
rect 322202 336016 322258 336025
rect 322202 335951 322258 335960
rect 321560 334620 321612 334626
rect 321560 334562 321612 334568
rect 323596 332382 323624 423642
rect 324976 419490 325004 639270
rect 327736 599282 327764 642466
rect 331864 642252 331916 642258
rect 331864 642194 331916 642200
rect 329104 642184 329156 642190
rect 329104 642126 329156 642132
rect 327816 641912 327868 641918
rect 327816 641854 327868 641860
rect 327724 599276 327776 599282
rect 327724 599218 327776 599224
rect 325608 596828 325660 596834
rect 325608 596770 325660 596776
rect 325620 596154 325648 596770
rect 325608 596148 325660 596154
rect 325608 596090 325660 596096
rect 327724 594176 327776 594182
rect 327724 594118 327776 594124
rect 325516 549296 325568 549302
rect 325516 549238 325568 549244
rect 325056 519308 325108 519314
rect 325056 519250 325108 519256
rect 325068 498846 325096 519250
rect 325528 517682 325556 549238
rect 326344 543108 326396 543114
rect 326344 543050 326396 543056
rect 326356 526998 326384 543050
rect 326344 526992 326396 526998
rect 326344 526934 326396 526940
rect 325516 517676 325568 517682
rect 325516 517618 325568 517624
rect 327736 509182 327764 594118
rect 327828 574870 327856 641854
rect 329116 578950 329144 642126
rect 329748 590028 329800 590034
rect 329748 589970 329800 589976
rect 329104 578944 329156 578950
rect 329104 578886 329156 578892
rect 327816 574864 327868 574870
rect 327816 574806 327868 574812
rect 327816 549364 327868 549370
rect 327816 549306 327868 549312
rect 327724 509176 327776 509182
rect 327724 509118 327776 509124
rect 327828 508162 327856 549306
rect 329102 547088 329158 547097
rect 329102 547023 329158 547032
rect 329116 514078 329144 547023
rect 329564 533452 329616 533458
rect 329564 533394 329616 533400
rect 329576 532030 329604 533394
rect 329564 532024 329616 532030
rect 329564 531966 329616 531972
rect 329196 517540 329248 517546
rect 329196 517482 329248 517488
rect 329104 514072 329156 514078
rect 329104 514014 329156 514020
rect 327816 508156 327868 508162
rect 327816 508098 327868 508104
rect 329208 505102 329236 517482
rect 329760 506394 329788 589970
rect 331218 516760 331274 516769
rect 331218 516695 331274 516704
rect 331232 512650 331260 516695
rect 331876 513330 331904 642194
rect 331954 641880 332010 641889
rect 331954 641815 332010 641824
rect 331968 599214 331996 641815
rect 331956 599208 332008 599214
rect 331956 599150 332008 599156
rect 334624 591388 334676 591394
rect 334624 591330 334676 591336
rect 336096 591388 336148 591394
rect 336096 591330 336148 591336
rect 333888 587240 333940 587246
rect 333888 587182 333940 587188
rect 331956 585812 332008 585818
rect 331956 585754 332008 585760
rect 331968 515438 331996 585754
rect 332600 545760 332652 545766
rect 332600 545702 332652 545708
rect 332612 539578 332640 545702
rect 332600 539572 332652 539578
rect 332600 539514 332652 539520
rect 331956 515432 332008 515438
rect 331956 515374 332008 515380
rect 331864 513324 331916 513330
rect 331864 513266 331916 513272
rect 331220 512644 331272 512650
rect 331220 512586 331272 512592
rect 333900 511290 333928 587182
rect 334636 524414 334664 591330
rect 336004 577584 336056 577590
rect 336004 577526 336056 577532
rect 334624 524408 334676 524414
rect 334624 524350 334676 524356
rect 333888 511284 333940 511290
rect 333888 511226 333940 511232
rect 336016 507754 336044 577526
rect 336108 532030 336136 591330
rect 336096 532024 336148 532030
rect 336096 531966 336148 531972
rect 336004 507748 336056 507754
rect 336004 507690 336056 507696
rect 329748 506388 329800 506394
rect 329748 506330 329800 506336
rect 329760 505782 329788 506330
rect 329748 505776 329800 505782
rect 329748 505718 329800 505724
rect 329196 505096 329248 505102
rect 329196 505038 329248 505044
rect 337396 502314 337424 697546
rect 403716 670744 403768 670750
rect 403716 670686 403768 670692
rect 352840 663808 352892 663814
rect 352840 663750 352892 663756
rect 352656 662924 352708 662930
rect 352656 662866 352708 662872
rect 349804 662856 349856 662862
rect 349804 662798 349856 662804
rect 338764 640688 338816 640694
rect 338764 640630 338816 640636
rect 337476 596964 337528 596970
rect 337476 596906 337528 596912
rect 337488 535294 337516 596906
rect 337476 535288 337528 535294
rect 337476 535230 337528 535236
rect 337936 534744 337988 534750
rect 337936 534686 337988 534692
rect 337948 530641 337976 534686
rect 338028 533452 338080 533458
rect 338028 533394 338080 533400
rect 338040 531282 338068 533394
rect 338028 531276 338080 531282
rect 338028 531218 338080 531224
rect 337934 530632 337990 530641
rect 337934 530567 337990 530576
rect 337384 502308 337436 502314
rect 337384 502250 337436 502256
rect 325056 498840 325108 498846
rect 325056 498782 325108 498788
rect 332600 482316 332652 482322
rect 332600 482258 332652 482264
rect 324964 419484 325016 419490
rect 324964 419426 325016 419432
rect 332612 345014 332640 482258
rect 338776 471986 338804 640630
rect 347688 596964 347740 596970
rect 347688 596906 347740 596912
rect 341524 595536 341576 595542
rect 341524 595478 341576 595484
rect 338856 588668 338908 588674
rect 338856 588610 338908 588616
rect 338868 529854 338896 588610
rect 340144 585880 340196 585886
rect 340144 585822 340196 585828
rect 338856 529848 338908 529854
rect 338856 529790 338908 529796
rect 340156 517478 340184 585822
rect 340144 517472 340196 517478
rect 340144 517414 340196 517420
rect 341536 505102 341564 595478
rect 343548 594176 343600 594182
rect 343548 594118 343600 594124
rect 342168 588668 342220 588674
rect 342168 588610 342220 588616
rect 342180 550730 342208 588610
rect 342904 587172 342956 587178
rect 342904 587114 342956 587120
rect 341616 550724 341668 550730
rect 341616 550666 341668 550672
rect 342168 550724 342220 550730
rect 342168 550666 342220 550672
rect 341628 510610 341656 550666
rect 342260 516112 342312 516118
rect 342260 516054 342312 516060
rect 342272 515438 342300 516054
rect 342260 515432 342312 515438
rect 342260 515374 342312 515380
rect 342916 514758 342944 587114
rect 342996 532024 343048 532030
rect 342996 531966 343048 531972
rect 342904 514752 342956 514758
rect 342904 514694 342956 514700
rect 343008 510610 343036 531966
rect 343560 515438 343588 594118
rect 345664 594108 345716 594114
rect 345664 594050 345716 594056
rect 343548 515432 343600 515438
rect 343548 515374 343600 515380
rect 341616 510604 341668 510610
rect 341616 510546 341668 510552
rect 342996 510604 343048 510610
rect 342996 510546 343048 510552
rect 345676 509114 345704 594050
rect 347044 592680 347096 592686
rect 347044 592622 347096 592628
rect 345756 584452 345808 584458
rect 345756 584394 345808 584400
rect 345768 532642 345796 584394
rect 345846 541104 345902 541113
rect 345846 541039 345902 541048
rect 345756 532636 345808 532642
rect 345756 532578 345808 532584
rect 345860 511902 345888 541039
rect 347056 536790 347084 592622
rect 347136 552832 347188 552838
rect 347136 552774 347188 552780
rect 347044 536784 347096 536790
rect 347044 536726 347096 536732
rect 347044 520328 347096 520334
rect 347044 520270 347096 520276
rect 345848 511896 345900 511902
rect 345848 511838 345900 511844
rect 345664 509108 345716 509114
rect 345664 509050 345716 509056
rect 341524 505096 341576 505102
rect 341524 505038 341576 505044
rect 347056 500886 347084 520270
rect 347148 503674 347176 552774
rect 347228 540320 347280 540326
rect 347228 540262 347280 540268
rect 347240 511902 347268 540262
rect 347700 520198 347728 596906
rect 348424 552084 348476 552090
rect 348424 552026 348476 552032
rect 348436 522986 348464 552026
rect 348516 525088 348568 525094
rect 348516 525030 348568 525036
rect 348424 522980 348476 522986
rect 348424 522922 348476 522928
rect 347688 520192 347740 520198
rect 347688 520134 347740 520140
rect 347228 511896 347280 511902
rect 347228 511838 347280 511844
rect 347136 503668 347188 503674
rect 347136 503610 347188 503616
rect 347044 500880 347096 500886
rect 347044 500822 347096 500828
rect 348528 497185 348556 525030
rect 349068 504212 349120 504218
rect 349068 504154 349120 504160
rect 349080 503742 349108 504154
rect 349068 503736 349120 503742
rect 349068 503678 349120 503684
rect 349080 497622 349108 503678
rect 349068 497616 349120 497622
rect 349068 497558 349120 497564
rect 349816 497282 349844 662798
rect 352564 662584 352616 662590
rect 352564 662526 352616 662532
rect 349896 642388 349948 642394
rect 349896 642330 349948 642336
rect 349908 497418 349936 642330
rect 349988 641776 350040 641782
rect 349988 641718 350040 641724
rect 350000 599010 350028 641718
rect 349988 599004 350040 599010
rect 349988 598946 350040 598952
rect 349988 595536 350040 595542
rect 349988 595478 350040 595484
rect 350000 504218 350028 595478
rect 350080 588600 350132 588606
rect 350080 588542 350132 588548
rect 350092 518906 350120 588542
rect 350448 565276 350500 565282
rect 350448 565218 350500 565224
rect 350172 541680 350224 541686
rect 350172 541622 350224 541628
rect 350080 518900 350132 518906
rect 350080 518842 350132 518848
rect 350080 509924 350132 509930
rect 350080 509866 350132 509872
rect 349988 504212 350040 504218
rect 349988 504154 350040 504160
rect 350092 497486 350120 509866
rect 350184 506394 350212 541622
rect 350460 531298 350488 565218
rect 351276 550860 351328 550866
rect 351276 550802 351328 550808
rect 351184 550656 351236 550662
rect 351184 550598 351236 550604
rect 350460 531270 350580 531298
rect 350552 530602 350580 531270
rect 350540 530596 350592 530602
rect 350540 530538 350592 530544
rect 350172 506388 350224 506394
rect 350172 506330 350224 506336
rect 350080 497480 350132 497486
rect 350080 497422 350132 497428
rect 349896 497412 349948 497418
rect 349896 497354 349948 497360
rect 349804 497276 349856 497282
rect 349804 497218 349856 497224
rect 348514 497176 348570 497185
rect 348514 497111 348570 497120
rect 350092 496913 350120 497422
rect 350078 496904 350134 496913
rect 350078 496839 350134 496848
rect 349712 487892 349764 487898
rect 349712 487834 349764 487840
rect 338764 471980 338816 471986
rect 338764 471922 338816 471928
rect 346492 347812 346544 347818
rect 346492 347754 346544 347760
rect 332612 344986 333192 345014
rect 332232 335368 332284 335374
rect 332232 335310 332284 335316
rect 323584 332376 323636 332382
rect 323584 332318 323636 332324
rect 325148 332376 325200 332382
rect 325148 332318 325200 332324
rect 320640 332036 320692 332042
rect 320640 331978 320692 331984
rect 320652 329868 320680 331978
rect 321928 331832 321980 331838
rect 321928 331774 321980 331780
rect 321940 329868 321968 331774
rect 323216 331492 323268 331498
rect 323216 331434 323268 331440
rect 323228 329868 323256 331434
rect 325160 329868 325188 332318
rect 330944 331560 330996 331566
rect 330944 331502 330996 331508
rect 327724 331424 327776 331430
rect 327724 331366 327776 331372
rect 326436 330200 326488 330206
rect 326436 330142 326488 330148
rect 326448 329868 326476 330142
rect 327736 329868 327764 331366
rect 329012 330132 329064 330138
rect 329012 330074 329064 330080
rect 329024 329868 329052 330074
rect 330956 329868 330984 331502
rect 332244 329868 332272 335310
rect 333164 329882 333192 344986
rect 341892 331696 341944 331702
rect 341892 331638 341944 331644
rect 339316 331560 339368 331566
rect 339316 331502 339368 331508
rect 336096 331492 336148 331498
rect 336096 331434 336148 331440
rect 334532 330064 334584 330070
rect 334532 330006 334584 330012
rect 334544 329882 334572 330006
rect 333164 329854 333546 329882
rect 334544 329854 334834 329882
rect 336108 329868 336136 331434
rect 338028 331356 338080 331362
rect 338028 331298 338080 331304
rect 338040 329868 338068 331298
rect 339328 329868 339356 331502
rect 340236 329996 340288 330002
rect 340236 329938 340288 329944
rect 340248 329882 340276 329938
rect 340248 329854 340630 329882
rect 341904 329868 341932 331638
rect 345112 331288 345164 331294
rect 345112 331230 345164 331236
rect 343640 329928 343692 329934
rect 343692 329876 343850 329882
rect 343640 329870 343850 329876
rect 343652 329854 343850 329870
rect 345124 329868 345152 331230
rect 346504 329882 346532 347754
rect 347688 332308 347740 332314
rect 347688 332250 347740 332256
rect 346426 329854 346532 329882
rect 347700 329868 347728 332250
rect 348974 331528 349030 331537
rect 348974 331463 349030 331472
rect 348988 329868 349016 331463
rect 349724 316010 349752 487834
rect 349988 411324 350040 411330
rect 349988 411266 350040 411272
rect 349804 341556 349856 341562
rect 349804 341498 349856 341504
rect 349816 318782 349844 341498
rect 349896 331288 349948 331294
rect 349896 331230 349948 331236
rect 349908 318794 349936 331230
rect 350000 321554 350028 411266
rect 350080 349852 350132 349858
rect 350080 349794 350132 349800
rect 350092 327729 350120 349794
rect 350264 338768 350316 338774
rect 350264 338710 350316 338716
rect 350172 333260 350224 333266
rect 350172 333202 350224 333208
rect 350078 327720 350134 327729
rect 350078 327655 350134 327664
rect 350184 325694 350212 333202
rect 350276 329089 350304 338710
rect 350262 329080 350318 329089
rect 350262 329015 350318 329024
rect 350184 325666 350396 325694
rect 350000 321526 350304 321554
rect 349804 318776 349856 318782
rect 349908 318766 350212 318794
rect 349804 318718 349856 318724
rect 349988 318708 350040 318714
rect 349988 318650 350040 318656
rect 349802 316024 349858 316033
rect 349724 315982 349802 316010
rect 349802 315959 349858 315968
rect 349802 312216 349858 312225
rect 349724 312174 349802 312202
rect 299848 295180 299900 295186
rect 299848 295122 299900 295128
rect 299756 278384 299808 278390
rect 299756 278326 299808 278332
rect 299664 276140 299716 276146
rect 299664 276082 299716 276088
rect 299572 271176 299624 271182
rect 299572 271118 299624 271124
rect 299860 223038 299888 295122
rect 300124 280628 300176 280634
rect 300124 280570 300176 280576
rect 300044 277642 300072 280092
rect 300032 277636 300084 277642
rect 300032 277578 300084 277584
rect 300136 277394 300164 280570
rect 301332 278730 301360 280092
rect 302252 280078 302634 280106
rect 301320 278724 301372 278730
rect 301320 278666 301372 278672
rect 299952 277366 300164 277394
rect 299952 223514 299980 277366
rect 301504 258732 301556 258738
rect 301504 258674 301556 258680
rect 299940 223508 299992 223514
rect 299940 223450 299992 223456
rect 299848 223032 299900 223038
rect 299848 222974 299900 222980
rect 301516 222290 301544 258674
rect 302252 223242 302280 280078
rect 303804 279948 303856 279954
rect 303804 279890 303856 279896
rect 303712 278180 303764 278186
rect 303712 278122 303764 278128
rect 302332 257372 302384 257378
rect 302332 257314 302384 257320
rect 302344 229094 302372 257314
rect 302344 229066 302464 229094
rect 302240 223236 302292 223242
rect 302240 223178 302292 223184
rect 301504 222284 301556 222290
rect 301504 222226 301556 222232
rect 299480 222148 299532 222154
rect 299480 222090 299532 222096
rect 300768 222148 300820 222154
rect 300768 222090 300820 222096
rect 300780 220862 300808 222090
rect 300768 220856 300820 220862
rect 300768 220798 300820 220804
rect 299388 220312 299440 220318
rect 299388 220254 299440 220260
rect 299294 101008 299350 101017
rect 299294 100943 299350 100952
rect 298834 93528 298890 93537
rect 298834 93463 298890 93472
rect 298006 90536 298062 90545
rect 298006 90471 298062 90480
rect 297364 90364 297416 90370
rect 297364 90306 297416 90312
rect 296812 89004 296864 89010
rect 296812 88946 296864 88952
rect 296824 84561 296852 88946
rect 297180 86964 297232 86970
rect 297180 86906 297232 86912
rect 297192 86057 297220 86906
rect 297178 86048 297234 86057
rect 297178 85983 297234 85992
rect 296810 84552 296866 84561
rect 296810 84487 296866 84496
rect 297180 77240 297232 77246
rect 297180 77182 297232 77188
rect 297192 77081 297220 77182
rect 297178 77072 297234 77081
rect 297178 77007 297234 77016
rect 296812 73160 296864 73166
rect 296812 73102 296864 73108
rect 296824 72593 296852 73102
rect 296810 72584 296866 72593
rect 296810 72519 296866 72528
rect 297180 69012 297232 69018
rect 297180 68954 297232 68960
rect 297192 68105 297220 68954
rect 297178 68096 297234 68105
rect 297178 68031 297234 68040
rect 297376 65113 297404 90306
rect 299400 89049 299428 220254
rect 300780 219980 300808 220798
rect 301516 219994 301544 222226
rect 302436 219994 302464 229066
rect 303724 219994 303752 278122
rect 303816 229094 303844 279890
rect 303908 278322 303936 280092
rect 305196 278662 305224 280092
rect 306668 280078 307142 280106
rect 305184 278656 305236 278662
rect 305184 278598 305236 278604
rect 303896 278316 303948 278322
rect 303896 278258 303948 278264
rect 305644 277636 305696 277642
rect 305644 277578 305696 277584
rect 305000 276140 305052 276146
rect 305000 276082 305052 276088
rect 305012 229094 305040 276082
rect 303816 229066 304488 229094
rect 305012 229066 305408 229094
rect 304460 219994 304488 229066
rect 305380 219994 305408 229066
rect 305656 223582 305684 277578
rect 306668 258074 306696 280078
rect 308416 278730 308444 280092
rect 309244 280078 309718 280106
rect 310624 280078 311006 280106
rect 311912 280078 312294 280106
rect 313292 280078 314226 280106
rect 308404 278724 308456 278730
rect 308404 278666 308456 278672
rect 309140 276820 309192 276826
rect 309140 276762 309192 276768
rect 306392 258046 306696 258074
rect 305644 223576 305696 223582
rect 305644 223518 305696 223524
rect 306392 220318 306420 258046
rect 308864 225616 308916 225622
rect 308864 225558 308916 225564
rect 307852 223576 307904 223582
rect 307852 223518 307904 223524
rect 306840 223508 306892 223514
rect 306840 223450 306892 223456
rect 306380 220312 306432 220318
rect 306380 220254 306432 220260
rect 301516 219966 301806 219994
rect 302436 219966 302818 219994
rect 303724 219966 303830 219994
rect 304460 219966 304842 219994
rect 305380 219966 305854 219994
rect 306852 219980 306880 223450
rect 307864 219980 307892 223518
rect 308876 219980 308904 225558
rect 309152 220130 309180 276762
rect 309244 223174 309272 280078
rect 310520 279472 310572 279478
rect 310520 279414 310572 279420
rect 309232 223168 309284 223174
rect 309232 223110 309284 223116
rect 309152 220102 309456 220130
rect 309428 219994 309456 220102
rect 310532 219994 310560 279414
rect 310624 233918 310652 280078
rect 311164 275392 311216 275398
rect 311164 275334 311216 275340
rect 310612 233912 310664 233918
rect 310612 233854 310664 233860
rect 311176 222902 311204 275334
rect 311912 235278 311940 280078
rect 311900 235272 311952 235278
rect 311900 235214 311952 235220
rect 311164 222896 311216 222902
rect 311164 222838 311216 222844
rect 312912 222896 312964 222902
rect 312912 222838 312964 222844
rect 311900 222828 311952 222834
rect 311900 222770 311952 222776
rect 309428 219966 309902 219994
rect 310532 219966 310914 219994
rect 311912 219980 311940 222770
rect 312924 219980 312952 222838
rect 313292 220250 313320 280078
rect 315500 279070 315528 280092
rect 315488 279064 315540 279070
rect 315488 279006 315540 279012
rect 316788 278730 316816 280092
rect 313372 278724 313424 278730
rect 313372 278666 313424 278672
rect 316776 278724 316828 278730
rect 316776 278666 316828 278672
rect 313384 229094 313412 278666
rect 318076 278390 318104 280092
rect 320008 278526 320036 280092
rect 321296 279002 321324 280092
rect 321652 279472 321704 279478
rect 321652 279414 321704 279420
rect 321284 278996 321336 279002
rect 321284 278938 321336 278944
rect 319996 278520 320048 278526
rect 319996 278462 320048 278468
rect 318064 278384 318116 278390
rect 318064 278326 318116 278332
rect 317420 278044 317472 278050
rect 317420 277986 317472 277992
rect 314752 276820 314804 276826
rect 314752 276762 314804 276768
rect 314764 229094 314792 276762
rect 317432 229094 317460 277986
rect 318800 271176 318852 271182
rect 318800 271118 318852 271124
rect 313384 229066 313504 229094
rect 314764 229066 315528 229094
rect 317432 229066 317552 229094
rect 313280 220244 313332 220250
rect 313280 220186 313332 220192
rect 313476 219994 313504 229066
rect 314936 223236 314988 223242
rect 314936 223178 314988 223184
rect 313476 219966 313950 219994
rect 314948 219980 314976 223178
rect 315500 219994 315528 229066
rect 316960 222896 317012 222902
rect 316960 222838 317012 222844
rect 315500 219966 315974 219994
rect 316972 219980 317000 222838
rect 317524 219994 317552 229066
rect 318812 224330 318840 271118
rect 318892 260160 318944 260166
rect 318892 260102 318944 260108
rect 318800 224324 318852 224330
rect 318800 224266 318852 224272
rect 318904 219994 318932 260102
rect 319628 224324 319680 224330
rect 319628 224266 319680 224272
rect 319640 219994 319668 224266
rect 321008 223032 321060 223038
rect 321008 222974 321060 222980
rect 317524 219966 317998 219994
rect 318904 219966 319010 219994
rect 319640 219966 320022 219994
rect 321020 219980 321048 222974
rect 321664 219994 321692 279414
rect 322584 278458 322612 280092
rect 323124 278724 323176 278730
rect 323124 278666 323176 278672
rect 322572 278452 322624 278458
rect 322572 278394 322624 278400
rect 323136 229094 323164 278666
rect 323872 277574 323900 280092
rect 324700 280078 325174 280106
rect 323860 277568 323912 277574
rect 323860 277510 323912 277516
rect 324320 277432 324372 277438
rect 324320 277374 324372 277380
rect 323136 229066 323624 229094
rect 323032 223168 323084 223174
rect 323032 223110 323084 223116
rect 321664 219966 322046 219994
rect 323044 219980 323072 223110
rect 323596 219994 323624 229066
rect 324332 220130 324360 277374
rect 324700 258074 324728 280078
rect 326344 277568 326396 277574
rect 326344 277510 326396 277516
rect 324424 258046 324728 258074
rect 324424 228410 324452 258046
rect 324412 228404 324464 228410
rect 324412 228346 324464 228352
rect 326068 228404 326120 228410
rect 326068 228346 326120 228352
rect 324332 220102 324728 220130
rect 324700 219994 324728 220102
rect 323596 219966 324070 219994
rect 324700 219966 325082 219994
rect 326080 219980 326108 228346
rect 326356 223106 326384 277510
rect 327092 277438 327120 280092
rect 328012 280078 328394 280106
rect 329300 280078 329682 280106
rect 327080 277432 327132 277438
rect 327080 277374 327132 277380
rect 328012 258074 328040 280078
rect 329300 258074 329328 280078
rect 330956 278934 330984 280092
rect 332612 280078 332902 280106
rect 330944 278928 330996 278934
rect 330944 278870 330996 278876
rect 327276 258046 328040 258074
rect 328472 258046 329328 258074
rect 326344 223100 326396 223106
rect 326344 223042 326396 223048
rect 327276 219994 327304 258046
rect 328092 223168 328144 223174
rect 328092 223110 328144 223116
rect 327106 219966 327304 219994
rect 328104 219980 328132 223110
rect 328472 220182 328500 258046
rect 332612 225622 332640 280078
rect 334176 278118 334204 280092
rect 335464 278594 335492 280092
rect 336766 280078 336964 280106
rect 335452 278588 335504 278594
rect 335452 278530 335504 278536
rect 334164 278112 334216 278118
rect 334164 278054 334216 278060
rect 335360 274032 335412 274038
rect 335360 273974 335412 273980
rect 333980 272672 334032 272678
rect 333980 272614 334032 272620
rect 333992 229094 334020 272614
rect 335372 229094 335400 273974
rect 333992 229066 334848 229094
rect 335372 229066 335768 229094
rect 332600 225616 332652 225622
rect 332600 225558 332652 225564
rect 329104 223236 329156 223242
rect 329104 223178 329156 223184
rect 328460 220176 328512 220182
rect 328460 220118 328512 220124
rect 329116 219980 329144 223178
rect 333152 223100 333204 223106
rect 333152 223042 333204 223048
rect 334164 223100 334216 223106
rect 334164 223042 334216 223048
rect 331128 223032 331180 223038
rect 331128 222974 331180 222980
rect 330116 222964 330168 222970
rect 330116 222906 330168 222912
rect 330128 219980 330156 222906
rect 331140 219980 331168 222974
rect 332140 222964 332192 222970
rect 332140 222906 332192 222912
rect 332152 219980 332180 222906
rect 333164 219980 333192 223042
rect 334176 219980 334204 223042
rect 334820 219994 334848 229066
rect 335740 219994 335768 229066
rect 336936 221610 336964 280078
rect 337384 278384 337436 278390
rect 337384 278326 337436 278332
rect 337200 223236 337252 223242
rect 337200 223178 337252 223184
rect 336924 221604 336976 221610
rect 336924 221546 336976 221552
rect 334820 219966 335202 219994
rect 335740 219966 336214 219994
rect 337212 219980 337240 223178
rect 337396 221542 337424 278326
rect 338040 278254 338068 280092
rect 339972 278662 340000 280092
rect 339960 278656 340012 278662
rect 339960 278598 340012 278604
rect 341260 278390 341288 280092
rect 342548 278866 342576 280092
rect 342536 278860 342588 278866
rect 342536 278802 342588 278808
rect 341248 278384 341300 278390
rect 341248 278326 341300 278332
rect 338028 278248 338080 278254
rect 338028 278190 338080 278196
rect 338212 278112 338264 278118
rect 338212 278054 338264 278060
rect 337384 221536 337436 221542
rect 337384 221478 337436 221484
rect 338224 219980 338252 278054
rect 343836 278050 343864 280092
rect 343824 278044 343876 278050
rect 343824 277986 343876 277992
rect 345768 277982 345796 280092
rect 347056 278730 347084 280092
rect 347884 280078 348358 280106
rect 347044 278724 347096 278730
rect 347044 278666 347096 278672
rect 345756 277976 345808 277982
rect 345756 277918 345808 277924
rect 347884 258074 347912 280078
rect 349632 278798 349660 280092
rect 349620 278792 349672 278798
rect 349620 278734 349672 278740
rect 347792 258046 347912 258074
rect 347792 253230 347820 258046
rect 347780 253224 347832 253230
rect 347780 253166 347832 253172
rect 349724 228410 349752 312174
rect 350000 312186 350028 318650
rect 349802 312151 349858 312160
rect 349988 312180 350040 312186
rect 349988 312122 350040 312128
rect 349804 312112 349856 312118
rect 350184 312066 350212 318766
rect 349804 312054 349856 312060
rect 349816 290873 349844 312054
rect 349908 312038 350212 312066
rect 349802 290864 349858 290873
rect 349802 290799 349858 290808
rect 349802 286376 349858 286385
rect 349802 286311 349858 286320
rect 349816 272678 349844 286311
rect 349804 272672 349856 272678
rect 349804 272614 349856 272620
rect 349712 228404 349764 228410
rect 349712 228346 349764 228352
rect 349908 223106 349936 312038
rect 350078 310856 350134 310865
rect 350078 310791 350134 310800
rect 350092 223242 350120 310791
rect 350276 309126 350304 321526
rect 350264 309120 350316 309126
rect 350264 309062 350316 309068
rect 350368 303929 350396 325666
rect 350354 303920 350410 303929
rect 350354 303855 350410 303864
rect 350080 223236 350132 223242
rect 350080 223178 350132 223184
rect 349896 223100 349948 223106
rect 349896 223042 349948 223048
rect 339224 222216 339276 222222
rect 339224 222158 339276 222164
rect 339236 219980 339264 222158
rect 341062 147520 341118 147529
rect 341062 147455 341118 147464
rect 340142 145344 340198 145353
rect 340142 145279 340198 145288
rect 340050 129976 340106 129985
rect 340050 129911 340106 129920
rect 299386 89040 299442 89049
rect 299386 88975 299442 88984
rect 298008 88324 298060 88330
rect 298008 88266 298060 88272
rect 298020 87553 298048 88266
rect 298006 87544 298062 87553
rect 298006 87479 298062 87488
rect 297916 84176 297968 84182
rect 297916 84118 297968 84124
rect 297928 83065 297956 84118
rect 297914 83056 297970 83065
rect 297914 82991 297970 83000
rect 297916 82816 297968 82822
rect 297916 82758 297968 82764
rect 297928 81569 297956 82758
rect 297914 81560 297970 81569
rect 297914 81495 297970 81504
rect 298006 80064 298062 80073
rect 298006 79999 298008 80008
rect 298060 79999 298062 80008
rect 298008 79970 298060 79976
rect 297548 78668 297600 78674
rect 297548 78610 297600 78616
rect 297560 78577 297588 78610
rect 297546 78568 297602 78577
rect 297546 78503 297602 78512
rect 298008 75880 298060 75886
rect 298008 75822 298060 75828
rect 298020 75585 298048 75822
rect 298006 75576 298062 75585
rect 298006 75511 298062 75520
rect 298008 74520 298060 74526
rect 298008 74462 298060 74468
rect 298020 74089 298048 74462
rect 298006 74080 298062 74089
rect 298006 74015 298062 74024
rect 297732 71732 297784 71738
rect 297732 71674 297784 71680
rect 297744 71097 297772 71674
rect 297730 71088 297786 71097
rect 297730 71023 297786 71032
rect 298008 70372 298060 70378
rect 298008 70314 298060 70320
rect 298020 69601 298048 70314
rect 298006 69592 298062 69601
rect 298006 69527 298062 69536
rect 297548 67584 297600 67590
rect 297548 67526 297600 67532
rect 297560 66609 297588 67526
rect 297546 66600 297602 66609
rect 297546 66535 297602 66544
rect 297362 65104 297418 65113
rect 297362 65039 297418 65048
rect 297916 64864 297968 64870
rect 297916 64806 297968 64812
rect 297928 63617 297956 64806
rect 297914 63608 297970 63617
rect 297914 63543 297970 63552
rect 298006 62112 298062 62121
rect 298006 62047 298008 62056
rect 298060 62047 298062 62056
rect 298008 62018 298060 62024
rect 296628 60376 296680 60382
rect 296628 60318 296680 60324
rect 303620 60376 303672 60382
rect 303620 60318 303672 60324
rect 295248 60308 295300 60314
rect 295248 60250 295300 60256
rect 303632 16574 303660 60318
rect 310520 60308 310572 60314
rect 310520 60250 310572 60256
rect 314660 60308 314712 60314
rect 314660 60250 314712 60256
rect 310532 16574 310560 60250
rect 292592 16546 293264 16574
rect 303632 16546 303936 16574
rect 310532 16546 311480 16574
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 297270 3632 297326 3641
rect 297270 3567 297326 3576
rect 300766 3632 300822 3641
rect 300766 3567 300822 3576
rect 297284 480 297312 3567
rect 300780 480 300808 3567
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 354 303936 16546
rect 307944 3868 307996 3874
rect 307944 3810 307996 3816
rect 307956 480 307984 3810
rect 311452 480 311480 16546
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 60250
rect 317418 60072 317474 60081
rect 317418 60007 317474 60016
rect 317432 16574 317460 60007
rect 340064 42226 340092 129911
rect 340156 58886 340184 145279
rect 340878 140992 340934 141001
rect 340878 140927 340934 140936
rect 340234 138816 340290 138825
rect 340234 138751 340290 138760
rect 340144 58880 340196 58886
rect 340144 58822 340196 58828
rect 340248 55962 340276 138751
rect 340326 119232 340382 119241
rect 340326 119167 340382 119176
rect 340236 55956 340288 55962
rect 340236 55898 340288 55904
rect 340340 44878 340368 119167
rect 340418 110528 340474 110537
rect 340418 110463 340474 110472
rect 340432 55894 340460 110463
rect 340510 75712 340566 75721
rect 340510 75647 340566 75656
rect 340524 60042 340552 75647
rect 340512 60036 340564 60042
rect 340512 59978 340564 59984
rect 340420 55888 340472 55894
rect 340420 55830 340472 55836
rect 340328 44872 340380 44878
rect 340328 44814 340380 44820
rect 340052 42220 340104 42226
rect 340052 42162 340104 42168
rect 317432 16546 318104 16574
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 340892 10334 340920 140927
rect 340970 121408 341026 121417
rect 340970 121343 341026 121352
rect 340880 10328 340932 10334
rect 340880 10270 340932 10276
rect 340984 4894 341012 121343
rect 341076 51746 341104 147455
rect 343086 143168 343142 143177
rect 343086 143103 343142 143112
rect 342442 136640 342498 136649
rect 342442 136575 342498 136584
rect 342258 134464 342314 134473
rect 342258 134399 342314 134408
rect 341154 132288 341210 132297
rect 341154 132223 341210 132232
rect 341168 53106 341196 132223
rect 341338 114880 341394 114889
rect 341338 114815 341394 114824
rect 341246 112704 341302 112713
rect 341246 112639 341302 112648
rect 341156 53100 341208 53106
rect 341156 53042 341208 53048
rect 341064 51740 341116 51746
rect 341064 51682 341116 51688
rect 341260 42158 341288 112639
rect 341352 60178 341380 114815
rect 341430 104000 341486 104009
rect 341430 103935 341486 103944
rect 341340 60172 341392 60178
rect 341340 60114 341392 60120
rect 341444 57322 341472 103935
rect 341522 101824 341578 101833
rect 341522 101759 341578 101768
rect 341432 57316 341484 57322
rect 341432 57258 341484 57264
rect 341536 57254 341564 101759
rect 341614 99648 341670 99657
rect 341614 99583 341670 99592
rect 341628 58818 341656 99583
rect 341706 97472 341762 97481
rect 341706 97407 341762 97416
rect 341720 60110 341748 97407
rect 341708 60104 341760 60110
rect 341708 60046 341760 60052
rect 341616 58812 341668 58818
rect 341616 58754 341668 58760
rect 341524 57248 341576 57254
rect 341524 57190 341576 57196
rect 341248 42152 341300 42158
rect 341248 42094 341300 42100
rect 342272 7682 342300 134399
rect 342352 117292 342404 117298
rect 342352 117234 342404 117240
rect 342364 117065 342392 117234
rect 342350 117056 342406 117065
rect 342350 116991 342406 117000
rect 342352 108996 342404 109002
rect 342352 108938 342404 108944
rect 342364 108361 342392 108938
rect 342350 108352 342406 108361
rect 342350 108287 342406 108296
rect 342352 106276 342404 106282
rect 342352 106218 342404 106224
rect 342364 106185 342392 106218
rect 342350 106176 342406 106185
rect 342350 106111 342406 106120
rect 342350 93120 342406 93129
rect 342350 93055 342406 93064
rect 342364 79393 342392 93055
rect 342350 79384 342406 79393
rect 342350 79319 342406 79328
rect 342350 79248 342406 79257
rect 342350 79183 342406 79192
rect 342364 62778 342392 79183
rect 342456 62898 342484 136575
rect 342534 127936 342590 127945
rect 342534 127871 342590 127880
rect 342444 62892 342496 62898
rect 342444 62834 342496 62840
rect 342364 62750 342484 62778
rect 342350 62656 342406 62665
rect 342350 62591 342406 62600
rect 342364 62150 342392 62591
rect 342352 62144 342404 62150
rect 342352 62086 342404 62092
rect 342456 58682 342484 62750
rect 342444 58676 342496 58682
rect 342444 58618 342496 58624
rect 342548 54534 342576 127871
rect 342626 125760 342682 125769
rect 342626 125695 342682 125704
rect 342640 61538 342668 125695
rect 342718 123584 342774 123593
rect 342718 123519 342774 123528
rect 342628 61532 342680 61538
rect 342628 61474 342680 61480
rect 342732 60246 342760 123519
rect 342810 90944 342866 90953
rect 342810 90879 342866 90888
rect 342824 61470 342852 90879
rect 342902 88768 342958 88777
rect 342902 88703 342958 88712
rect 342812 61464 342864 61470
rect 342812 61406 342864 61412
rect 342916 61402 342944 88703
rect 342994 69184 343050 69193
rect 342994 69119 343050 69128
rect 343008 69086 343036 69119
rect 342996 69080 343048 69086
rect 342996 69022 343048 69028
rect 342994 67008 343050 67017
rect 342994 66943 343050 66952
rect 343008 66298 343036 66943
rect 342996 66292 343048 66298
rect 342996 66234 343048 66240
rect 342994 64832 343050 64841
rect 342994 64767 343050 64776
rect 343008 63578 343036 64767
rect 342996 63572 343048 63578
rect 342996 63514 343048 63520
rect 342996 62892 343048 62898
rect 342996 62834 343048 62840
rect 342904 61396 342956 61402
rect 342904 61338 342956 61344
rect 342720 60240 342772 60246
rect 342720 60182 342772 60188
rect 343008 57390 343036 62834
rect 342996 57384 343048 57390
rect 342996 57326 343048 57332
rect 342536 54528 342588 54534
rect 342536 54470 342588 54476
rect 343100 46238 343128 143103
rect 343178 86592 343234 86601
rect 343178 86527 343234 86536
rect 343192 58750 343220 86527
rect 343180 58744 343232 58750
rect 343180 58686 343232 58692
rect 343088 46232 343140 46238
rect 343088 46174 343140 46180
rect 349160 28348 349212 28354
rect 349160 28290 349212 28296
rect 346400 22772 346452 22778
rect 346400 22714 346452 22720
rect 346412 16574 346440 22714
rect 346412 16546 346992 16574
rect 342260 7676 342312 7682
rect 342260 7618 342312 7624
rect 340972 4888 341024 4894
rect 340972 4830 341024 4836
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 325608 4004 325660 4010
rect 325608 3946 325660 3952
rect 322112 3936 322164 3942
rect 322112 3878 322164 3884
rect 322124 480 322152 3878
rect 325620 480 325648 3946
rect 329194 3632 329250 3641
rect 329194 3567 329250 3576
rect 329208 480 329236 3567
rect 332704 480 332732 4082
rect 336280 4072 336332 4078
rect 336280 4014 336332 4020
rect 336292 480 336320 4014
rect 339868 3392 339920 3398
rect 339868 3334 339920 3340
rect 339880 480 339908 3334
rect 343364 3256 343416 3262
rect 343364 3198 343416 3204
rect 343376 480 343404 3198
rect 346964 480 346992 16546
rect 349172 3398 349200 28290
rect 350552 4010 350580 530538
rect 350724 517676 350776 517682
rect 350724 517618 350776 517624
rect 350632 517608 350684 517614
rect 350632 517550 350684 517556
rect 350644 4146 350672 517550
rect 350632 4140 350684 4146
rect 350632 4082 350684 4088
rect 350540 4004 350592 4010
rect 350540 3946 350592 3952
rect 350736 3942 350764 517618
rect 351196 506462 351224 550598
rect 351288 529922 351316 550802
rect 352380 549908 352432 549914
rect 352380 549850 352432 549856
rect 352392 535362 352420 549850
rect 352472 549568 352524 549574
rect 352472 549510 352524 549516
rect 352380 535356 352432 535362
rect 352380 535298 352432 535304
rect 352484 532710 352512 549510
rect 352472 532704 352524 532710
rect 352472 532646 352524 532652
rect 351276 529916 351328 529922
rect 351276 529858 351328 529864
rect 352472 522300 352524 522306
rect 352472 522242 352524 522248
rect 351276 520940 351328 520946
rect 351276 520882 351328 520888
rect 351184 506456 351236 506462
rect 351184 506398 351236 506404
rect 351288 497321 351316 520882
rect 352484 497826 352512 522242
rect 352576 497894 352604 662526
rect 352564 497888 352616 497894
rect 352564 497830 352616 497836
rect 352472 497820 352524 497826
rect 352472 497762 352524 497768
rect 352668 497350 352696 662866
rect 352748 662652 352800 662658
rect 352748 662594 352800 662600
rect 352760 497554 352788 662594
rect 352852 499254 352880 663750
rect 353024 662992 353076 662998
rect 353024 662934 353076 662940
rect 352932 641844 352984 641850
rect 352932 641786 352984 641792
rect 352944 499526 352972 641786
rect 353036 520266 353064 662934
rect 355416 662788 355468 662794
rect 355416 662730 355468 662736
rect 355324 662720 355376 662726
rect 355324 662662 355376 662668
rect 353116 642048 353168 642054
rect 353116 641990 353168 641996
rect 353128 599146 353156 641990
rect 354036 640552 354088 640558
rect 354036 640494 354088 640500
rect 354128 640552 354180 640558
rect 354128 640494 354180 640500
rect 353944 639124 353996 639130
rect 353944 639066 353996 639072
rect 353116 599140 353168 599146
rect 353116 599082 353168 599088
rect 353116 572076 353168 572082
rect 353116 572018 353168 572024
rect 353024 520260 353076 520266
rect 353024 520202 353076 520208
rect 353128 506462 353156 572018
rect 353208 550044 353260 550050
rect 353208 549986 353260 549992
rect 353220 521642 353248 549986
rect 353300 540252 353352 540258
rect 353300 540194 353352 540200
rect 353312 532710 353340 540194
rect 353300 532704 353352 532710
rect 353300 532646 353352 532652
rect 353298 530632 353354 530641
rect 353298 530567 353354 530576
rect 353312 529961 353340 530567
rect 353298 529952 353354 529961
rect 353298 529887 353354 529896
rect 353574 529952 353630 529961
rect 353574 529887 353630 529896
rect 353220 521626 353432 521642
rect 353208 521620 353432 521626
rect 353260 521614 353432 521620
rect 353208 521562 353260 521568
rect 353220 521531 353248 521562
rect 353116 506456 353168 506462
rect 353116 506398 353168 506404
rect 352932 499520 352984 499526
rect 352932 499462 352984 499468
rect 352840 499248 352892 499254
rect 352840 499190 352892 499196
rect 352748 497548 352800 497554
rect 352748 497490 352800 497496
rect 352656 497344 352708 497350
rect 351274 497312 351330 497321
rect 352656 497286 352708 497292
rect 351274 497247 351330 497256
rect 351920 491972 351972 491978
rect 351920 491914 351972 491920
rect 353300 491972 353352 491978
rect 353300 491914 353352 491920
rect 350908 429208 350960 429214
rect 350908 429150 350960 429156
rect 350816 400240 350868 400246
rect 350816 400182 350868 400188
rect 350828 280809 350856 400182
rect 350920 314129 350948 429150
rect 351092 376780 351144 376786
rect 351092 376722 351144 376728
rect 350998 325000 351054 325009
rect 350998 324935 351054 324944
rect 350906 314120 350962 314129
rect 350906 314055 350962 314064
rect 350906 291680 350962 291689
rect 350906 291615 350962 291624
rect 350814 280800 350870 280809
rect 350814 280735 350870 280744
rect 350920 258738 350948 291615
rect 351012 260166 351040 324935
rect 351104 317529 351132 376722
rect 351368 342916 351420 342922
rect 351368 342858 351420 342864
rect 351276 334688 351328 334694
rect 351276 334630 351328 334636
rect 351090 317520 351146 317529
rect 351090 317455 351146 317464
rect 351184 310616 351236 310622
rect 351184 310558 351236 310564
rect 351090 308000 351146 308009
rect 351090 307935 351146 307944
rect 351104 276826 351132 307935
rect 351092 276820 351144 276826
rect 351092 276762 351144 276768
rect 351000 260160 351052 260166
rect 351000 260102 351052 260108
rect 350908 258732 350960 258738
rect 350908 258674 350960 258680
rect 351196 222902 351224 310558
rect 351288 288289 351316 334630
rect 351380 299169 351408 342858
rect 351460 329860 351512 329866
rect 351460 329802 351512 329808
rect 351472 305289 351500 329802
rect 351932 326369 351960 491914
rect 352196 354000 352248 354006
rect 352196 353942 352248 353948
rect 352012 344344 352064 344350
rect 352012 344286 352064 344292
rect 351918 326360 351974 326369
rect 351918 326295 351974 326304
rect 351918 321600 351974 321609
rect 351918 321535 351974 321544
rect 351932 310622 351960 321535
rect 352024 318889 352052 344286
rect 352104 337408 352156 337414
rect 352104 337350 352156 337356
rect 352010 318880 352066 318889
rect 352010 318815 352066 318824
rect 351920 310616 351972 310622
rect 351920 310558 351972 310564
rect 351920 309120 351972 309126
rect 351920 309062 351972 309068
rect 351458 305280 351514 305289
rect 351458 305215 351514 305224
rect 351932 301889 351960 309062
rect 351918 301880 351974 301889
rect 351918 301815 351974 301824
rect 351918 300520 351974 300529
rect 351918 300455 351974 300464
rect 351366 299160 351422 299169
rect 351366 299095 351422 299104
rect 351368 291712 351420 291718
rect 351366 291680 351368 291689
rect 351420 291680 351422 291689
rect 351366 291615 351422 291624
rect 351274 288280 351330 288289
rect 351274 288215 351330 288224
rect 351932 280022 351960 300455
rect 352116 297809 352144 337350
rect 352102 297800 352158 297809
rect 352102 297735 352158 297744
rect 352010 294400 352066 294409
rect 352010 294335 352066 294344
rect 352024 281314 352052 294335
rect 352102 285560 352158 285569
rect 352102 285495 352158 285504
rect 352012 281308 352064 281314
rect 352012 281250 352064 281256
rect 351920 280016 351972 280022
rect 351920 279958 351972 279964
rect 352116 276758 352144 285495
rect 352208 282849 352236 353942
rect 352288 340196 352340 340202
rect 352288 340138 352340 340144
rect 352300 296449 352328 340138
rect 352564 334756 352616 334762
rect 352564 334698 352616 334704
rect 352472 333328 352524 333334
rect 352472 333270 352524 333276
rect 352378 323640 352434 323649
rect 352378 323575 352434 323584
rect 352286 296440 352342 296449
rect 352286 296375 352342 296384
rect 352286 293040 352342 293049
rect 352286 292975 352342 292984
rect 352194 282840 352250 282849
rect 352194 282775 352250 282784
rect 352104 276752 352156 276758
rect 352104 276694 352156 276700
rect 352300 236706 352328 292975
rect 352392 272610 352420 323575
rect 352484 284209 352512 333270
rect 352576 306649 352604 334698
rect 352656 331492 352708 331498
rect 352656 331434 352708 331440
rect 352562 306640 352618 306649
rect 352562 306575 352618 306584
rect 352470 284200 352526 284209
rect 352470 284135 352526 284144
rect 352380 272604 352432 272610
rect 352380 272546 352432 272552
rect 352288 236700 352340 236706
rect 352288 236642 352340 236648
rect 352668 223174 352696 331434
rect 352748 331424 352800 331430
rect 352748 331366 352800 331372
rect 352656 223168 352708 223174
rect 352656 223110 352708 223116
rect 352760 222970 352788 331366
rect 352838 310040 352894 310049
rect 352838 309975 352894 309984
rect 352748 222964 352800 222970
rect 352748 222906 352800 222912
rect 351184 222896 351236 222902
rect 351184 222838 351236 222844
rect 352852 221474 352880 309975
rect 352840 221468 352892 221474
rect 352840 221410 352892 221416
rect 350724 3936 350776 3942
rect 350724 3878 350776 3884
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 353312 354 353340 491914
rect 353404 3262 353432 521614
rect 353484 498840 353536 498846
rect 353484 498782 353536 498788
rect 353496 3330 353524 498782
rect 353588 291718 353616 529887
rect 353760 331968 353812 331974
rect 353760 331910 353812 331916
rect 353668 331356 353720 331362
rect 353668 331298 353720 331304
rect 353576 291712 353628 291718
rect 353576 291654 353628 291660
rect 353680 223038 353708 331298
rect 353772 278662 353800 331910
rect 353852 331900 353904 331906
rect 353852 331842 353904 331848
rect 353864 278730 353892 331842
rect 353852 278724 353904 278730
rect 353852 278666 353904 278672
rect 353760 278656 353812 278662
rect 353760 278598 353812 278604
rect 353668 223032 353720 223038
rect 353668 222974 353720 222980
rect 353956 60722 353984 639066
rect 354048 139398 354076 640494
rect 354140 598534 354168 640494
rect 354128 598528 354180 598534
rect 354128 598470 354180 598476
rect 354220 576224 354272 576230
rect 354220 576166 354272 576172
rect 354128 543040 354180 543046
rect 354128 542982 354180 542988
rect 354140 497758 354168 542982
rect 354232 535430 354260 576166
rect 354312 565140 354364 565146
rect 354312 565082 354364 565088
rect 354220 535424 354272 535430
rect 354220 535366 354272 535372
rect 354324 535362 354352 565082
rect 355232 552356 355284 552362
rect 355232 552298 355284 552304
rect 354404 552220 354456 552226
rect 354404 552162 354456 552168
rect 354312 535356 354364 535362
rect 354312 535298 354364 535304
rect 354416 527066 354444 552162
rect 355140 551676 355192 551682
rect 355140 551618 355192 551624
rect 355152 535226 355180 551618
rect 355140 535220 355192 535226
rect 355140 535162 355192 535168
rect 355244 528562 355272 552298
rect 355232 528556 355284 528562
rect 355232 528498 355284 528504
rect 355336 527066 355364 662662
rect 355428 536722 355456 662730
rect 403256 662516 403308 662522
rect 403256 662458 403308 662464
rect 356704 661496 356756 661502
rect 356704 661438 356756 661444
rect 355968 641980 356020 641986
rect 355968 641922 356020 641928
rect 355508 640824 355560 640830
rect 355508 640766 355560 640772
rect 355520 598398 355548 640766
rect 355508 598392 355560 598398
rect 355508 598334 355560 598340
rect 355600 554260 355652 554266
rect 355600 554202 355652 554208
rect 355508 544400 355560 544406
rect 355508 544342 355560 544348
rect 355416 536716 355468 536722
rect 355416 536658 355468 536664
rect 354404 527060 354456 527066
rect 354404 527002 354456 527008
rect 355324 527060 355376 527066
rect 355324 527002 355376 527008
rect 355232 523728 355284 523734
rect 355232 523670 355284 523676
rect 354220 520192 354272 520198
rect 354220 520134 354272 520140
rect 354232 498234 354260 520134
rect 354220 498228 354272 498234
rect 354220 498170 354272 498176
rect 354128 497752 354180 497758
rect 354128 497694 354180 497700
rect 355244 497593 355272 523670
rect 355416 515432 355468 515438
rect 355416 515374 355468 515380
rect 355324 513460 355376 513466
rect 355324 513402 355376 513408
rect 355336 497690 355364 513402
rect 355428 499118 355456 515374
rect 355416 499112 355468 499118
rect 355416 499054 355468 499060
rect 355428 498234 355456 499054
rect 355416 498228 355468 498234
rect 355416 498170 355468 498176
rect 355416 498092 355468 498098
rect 355416 498034 355468 498040
rect 355324 497684 355376 497690
rect 355324 497626 355376 497632
rect 355230 497584 355286 497593
rect 355230 497519 355286 497528
rect 354128 331560 354180 331566
rect 354128 331502 354180 331508
rect 354140 279478 354168 331502
rect 354128 279472 354180 279478
rect 354128 279414 354180 279420
rect 354036 139392 354088 139398
rect 354036 139334 354088 139340
rect 353944 60716 353996 60722
rect 353944 60658 353996 60664
rect 355336 3874 355364 497626
rect 355428 4078 355456 498034
rect 355520 497962 355548 544342
rect 355612 509250 355640 554202
rect 355784 554192 355836 554198
rect 355784 554134 355836 554140
rect 355692 549976 355744 549982
rect 355692 549918 355744 549924
rect 355600 509244 355652 509250
rect 355600 509186 355652 509192
rect 355704 507822 355732 549918
rect 355796 511970 355824 554134
rect 355876 550044 355928 550050
rect 355876 549986 355928 549992
rect 355888 517614 355916 549986
rect 355876 517608 355928 517614
rect 355876 517550 355928 517556
rect 355784 511964 355836 511970
rect 355784 511906 355836 511912
rect 355692 507816 355744 507822
rect 355692 507758 355744 507764
rect 355600 498228 355652 498234
rect 355600 498170 355652 498176
rect 355508 497956 355560 497962
rect 355508 497898 355560 497904
rect 355508 487824 355560 487830
rect 355508 487766 355560 487772
rect 355520 45558 355548 487766
rect 355612 60314 355640 498170
rect 355980 498030 356008 641922
rect 356716 552770 356744 661438
rect 358820 661428 358872 661434
rect 358820 661370 358872 661376
rect 358832 661337 358860 661370
rect 401600 661360 401652 661366
rect 358818 661328 358874 661337
rect 358818 661263 358874 661272
rect 401598 661328 401600 661337
rect 401652 661328 401654 661337
rect 401598 661263 401654 661272
rect 360936 642728 360988 642734
rect 360936 642670 360988 642676
rect 379428 642728 379480 642734
rect 379428 642670 379480 642676
rect 359556 642592 359608 642598
rect 359556 642534 359608 642540
rect 359464 642320 359516 642326
rect 359464 642262 359516 642268
rect 358820 642252 358872 642258
rect 358820 642194 358872 642200
rect 357348 642116 357400 642122
rect 357348 642058 357400 642064
rect 357072 640756 357124 640762
rect 357072 640698 357124 640704
rect 356980 640620 357032 640626
rect 356980 640562 357032 640568
rect 356796 640484 356848 640490
rect 356796 640426 356848 640432
rect 356704 552764 356756 552770
rect 356704 552706 356756 552712
rect 356612 552288 356664 552294
rect 356612 552230 356664 552236
rect 356624 548622 356652 552230
rect 356612 548616 356664 548622
rect 356612 548558 356664 548564
rect 356704 537532 356756 537538
rect 356704 537474 356756 537480
rect 356612 507884 356664 507890
rect 356612 507826 356664 507832
rect 356624 499497 356652 507826
rect 356716 503305 356744 537474
rect 356702 503296 356758 503305
rect 356702 503231 356758 503240
rect 356610 499488 356666 499497
rect 356610 499423 356666 499432
rect 355968 498024 356020 498030
rect 355968 497966 356020 497972
rect 355600 60308 355652 60314
rect 355600 60250 355652 60256
rect 355508 45552 355560 45558
rect 355508 45494 355560 45500
rect 356808 20602 356836 640426
rect 356888 639056 356940 639062
rect 356888 638998 356940 639004
rect 356900 179382 356928 638998
rect 356992 313274 357020 640562
rect 357084 598670 357112 640698
rect 357164 640620 357216 640626
rect 357164 640562 357216 640568
rect 357072 598664 357124 598670
rect 357072 598606 357124 598612
rect 357176 598602 357204 640562
rect 357164 598596 357216 598602
rect 357164 598538 357216 598544
rect 357072 569220 357124 569226
rect 357072 569162 357124 569168
rect 357084 550361 357112 569162
rect 357164 552152 357216 552158
rect 357164 552094 357216 552100
rect 357070 550352 357126 550361
rect 357070 550287 357126 550296
rect 357072 548548 357124 548554
rect 357072 548490 357124 548496
rect 357084 498166 357112 548490
rect 357176 533390 357204 552094
rect 357164 533384 357216 533390
rect 357164 533326 357216 533332
rect 357164 529984 357216 529990
rect 357164 529926 357216 529932
rect 357176 499186 357204 529926
rect 357256 511284 357308 511290
rect 357256 511226 357308 511232
rect 357164 499180 357216 499186
rect 357164 499122 357216 499128
rect 357268 499050 357296 511226
rect 357256 499044 357308 499050
rect 357256 498986 357308 498992
rect 357360 498914 357388 642058
rect 358636 639804 358688 639810
rect 358636 639746 358688 639752
rect 358452 639736 358504 639742
rect 358452 639678 358504 639684
rect 357808 639600 357860 639606
rect 357808 639542 357860 639548
rect 357530 548992 357586 549001
rect 357530 548927 357586 548936
rect 357440 547868 357492 547874
rect 357440 547810 357492 547816
rect 357452 547777 357480 547810
rect 357438 547768 357494 547777
rect 357438 547703 357494 547712
rect 357440 546440 357492 546446
rect 357440 546382 357492 546388
rect 357452 546281 357480 546382
rect 357438 546272 357494 546281
rect 357438 546207 357494 546216
rect 357440 545080 357492 545086
rect 357440 545022 357492 545028
rect 357452 544785 357480 545022
rect 357438 544776 357494 544785
rect 357438 544711 357494 544720
rect 357440 539572 357492 539578
rect 357440 539514 357492 539520
rect 357452 539209 357480 539514
rect 357438 539200 357494 539209
rect 357438 539135 357494 539144
rect 357440 536784 357492 536790
rect 357438 536752 357440 536761
rect 357492 536752 357494 536761
rect 357438 536687 357494 536696
rect 357544 535566 357572 548927
rect 357624 543788 357676 543794
rect 357624 543730 357676 543736
rect 357532 535560 357584 535566
rect 357532 535502 357584 535508
rect 357532 535424 357584 535430
rect 357438 535392 357494 535401
rect 357532 535366 357584 535372
rect 357438 535327 357494 535336
rect 357452 535294 357480 535327
rect 357440 535288 357492 535294
rect 357544 535265 357572 535366
rect 357440 535230 357492 535236
rect 357530 535256 357586 535265
rect 357530 535191 357586 535200
rect 357530 533488 357586 533497
rect 357530 533423 357532 533432
rect 357584 533423 357586 533432
rect 357532 533394 357584 533400
rect 357532 532704 357584 532710
rect 357532 532646 357584 532652
rect 357440 532636 357492 532642
rect 357440 532578 357492 532584
rect 357452 532409 357480 532578
rect 357438 532400 357494 532409
rect 357438 532335 357494 532344
rect 357544 531865 357572 532646
rect 357530 531856 357586 531865
rect 357530 531791 357586 531800
rect 357440 529848 357492 529854
rect 357440 529790 357492 529796
rect 357452 529553 357480 529790
rect 357438 529544 357494 529553
rect 357438 529479 357494 529488
rect 357440 527128 357492 527134
rect 357438 527096 357440 527105
rect 357492 527096 357494 527105
rect 357438 527031 357494 527040
rect 357532 527060 357584 527066
rect 357532 527002 357584 527008
rect 357544 526425 357572 527002
rect 357530 526416 357586 526425
rect 357530 526351 357586 526360
rect 357440 524408 357492 524414
rect 357440 524350 357492 524356
rect 357452 523705 357480 524350
rect 357438 523696 357494 523705
rect 357438 523631 357494 523640
rect 357636 521665 357664 543730
rect 357714 543552 357770 543561
rect 357714 543487 357770 543496
rect 357728 543114 357756 543487
rect 357716 543108 357768 543114
rect 357716 543050 357768 543056
rect 357714 539336 357770 539345
rect 357714 539271 357770 539280
rect 357622 521656 357678 521665
rect 357622 521591 357678 521600
rect 357440 520260 357492 520266
rect 357440 520202 357492 520208
rect 357452 519625 357480 520202
rect 357438 519616 357494 519625
rect 357438 519551 357494 519560
rect 357440 518900 357492 518906
rect 357440 518842 357492 518848
rect 357452 518809 357480 518842
rect 357438 518800 357494 518809
rect 357438 518735 357494 518744
rect 357530 517576 357586 517585
rect 357530 517511 357532 517520
rect 357584 517511 357586 517520
rect 357532 517482 357584 517488
rect 357440 517472 357492 517478
rect 357438 517440 357440 517449
rect 357492 517440 357494 517449
rect 357438 517375 357494 517384
rect 357440 514752 357492 514758
rect 357438 514720 357440 514729
rect 357492 514720 357494 514729
rect 357438 514655 357494 514664
rect 357530 513496 357586 513505
rect 357530 513431 357586 513440
rect 357440 513324 357492 513330
rect 357440 513266 357492 513272
rect 357452 512825 357480 513266
rect 357438 512816 357494 512825
rect 357438 512751 357494 512760
rect 357440 511896 357492 511902
rect 357440 511838 357492 511844
rect 357452 511465 357480 511838
rect 357438 511456 357494 511465
rect 357438 511391 357494 511400
rect 357440 510604 357492 510610
rect 357440 510546 357492 510552
rect 357452 510513 357480 510546
rect 357438 510504 357494 510513
rect 357438 510439 357494 510448
rect 357440 509108 357492 509114
rect 357440 509050 357492 509056
rect 357452 509017 357480 509050
rect 357438 509008 357494 509017
rect 357438 508943 357494 508952
rect 357440 507748 357492 507754
rect 357440 507690 357492 507696
rect 357452 507385 357480 507690
rect 357438 507376 357494 507385
rect 357438 507311 357494 507320
rect 357440 506456 357492 506462
rect 357438 506424 357440 506433
rect 357492 506424 357494 506433
rect 357438 506359 357494 506368
rect 357440 505096 357492 505102
rect 357440 505038 357492 505044
rect 357452 504665 357480 505038
rect 357438 504656 357494 504665
rect 357438 504591 357494 504600
rect 357440 502308 357492 502314
rect 357440 502250 357492 502256
rect 357452 501945 357480 502250
rect 357438 501936 357494 501945
rect 357438 501871 357494 501880
rect 357348 498908 357400 498914
rect 357348 498850 357400 498856
rect 357072 498160 357124 498166
rect 357072 498102 357124 498108
rect 357544 496398 357572 513431
rect 357624 506388 357676 506394
rect 357624 506330 357676 506336
rect 357636 505889 357664 506330
rect 357622 505880 357678 505889
rect 357622 505815 357678 505824
rect 357624 504416 357676 504422
rect 357624 504358 357676 504364
rect 357532 496392 357584 496398
rect 357532 496334 357584 496340
rect 356980 313268 357032 313274
rect 356980 313210 357032 313216
rect 356888 179376 356940 179382
rect 356888 179318 356940 179324
rect 357636 177410 357664 504358
rect 357624 177404 357676 177410
rect 357624 177346 357676 177352
rect 357728 109750 357756 539271
rect 357820 524657 357848 639542
rect 358268 565140 358320 565146
rect 358268 565082 358320 565088
rect 357900 556912 357952 556918
rect 357900 556854 357952 556860
rect 357912 545057 357940 556854
rect 358084 551744 358136 551750
rect 358084 551686 358136 551692
rect 357898 545048 357954 545057
rect 357898 544983 357954 544992
rect 358096 543561 358124 551686
rect 358176 551268 358228 551274
rect 358176 551210 358228 551216
rect 358082 543552 358138 543561
rect 358082 543487 358138 543496
rect 357900 536716 357952 536722
rect 357900 536658 357952 536664
rect 357912 536625 357940 536658
rect 357898 536616 357954 536625
rect 357898 536551 357954 536560
rect 357900 535356 357952 535362
rect 357900 535298 357952 535304
rect 357912 534585 357940 535298
rect 357898 534576 357954 534585
rect 357898 534511 357954 534520
rect 358188 528329 358216 551210
rect 358280 538121 358308 565082
rect 358360 563780 358412 563786
rect 358360 563722 358412 563728
rect 358266 538112 358322 538121
rect 358266 538047 358322 538056
rect 358280 537606 358308 538047
rect 358268 537600 358320 537606
rect 358268 537542 358320 537548
rect 358280 536926 358308 537542
rect 358268 536920 358320 536926
rect 358268 536862 358320 536868
rect 358372 533497 358400 563722
rect 358464 542337 358492 639678
rect 358544 639396 358596 639402
rect 358544 639338 358596 639344
rect 358450 542328 358506 542337
rect 358450 542263 358506 542272
rect 358556 540977 358584 639338
rect 358542 540968 358598 540977
rect 358542 540903 358598 540912
rect 358648 537985 358676 639746
rect 358728 550792 358780 550798
rect 358728 550734 358780 550740
rect 358740 548865 358768 550734
rect 358726 548856 358782 548865
rect 358726 548791 358782 548800
rect 358634 537976 358690 537985
rect 358634 537911 358690 537920
rect 358452 536852 358504 536858
rect 358452 536794 358504 536800
rect 358358 533488 358414 533497
rect 358358 533423 358414 533432
rect 358358 528592 358414 528601
rect 358358 528527 358414 528536
rect 358174 528320 358230 528329
rect 358174 528255 358230 528264
rect 358268 525836 358320 525842
rect 358268 525778 358320 525784
rect 357806 524648 357862 524657
rect 357806 524583 357862 524592
rect 357806 523832 357862 523841
rect 357806 523767 357862 523776
rect 357716 109744 357768 109750
rect 357716 109686 357768 109692
rect 357820 89010 357848 523767
rect 358082 519752 358138 519761
rect 358082 519687 358138 519696
rect 358096 511970 358124 519687
rect 358174 515128 358230 515137
rect 358174 515063 358230 515072
rect 358084 511964 358136 511970
rect 358084 511906 358136 511912
rect 357898 511592 357954 511601
rect 357898 511527 357954 511536
rect 357912 504422 357940 511527
rect 357992 509176 358044 509182
rect 357992 509118 358044 509124
rect 358004 508745 358032 509118
rect 357990 508736 358046 508745
rect 357990 508671 358046 508680
rect 357900 504416 357952 504422
rect 357900 504358 357952 504364
rect 358188 496194 358216 515063
rect 358280 503713 358308 525778
rect 358266 503704 358322 503713
rect 358266 503639 358322 503648
rect 358176 496188 358228 496194
rect 358176 496130 358228 496136
rect 358372 494766 358400 528527
rect 358464 507793 358492 536794
rect 358634 532808 358690 532817
rect 358634 532743 358690 532752
rect 358542 522472 358598 522481
rect 358542 522407 358598 522416
rect 358450 507784 358506 507793
rect 358450 507719 358506 507728
rect 358360 494760 358412 494766
rect 358360 494702 358412 494708
rect 358556 175982 358584 522407
rect 358648 514350 358676 532743
rect 358636 514344 358688 514350
rect 358636 514286 358688 514292
rect 358832 510105 358860 642194
rect 358912 641844 358964 641850
rect 358912 641786 358964 641792
rect 358924 543425 358952 641786
rect 359096 563848 359148 563854
rect 359096 563790 359148 563796
rect 359004 558272 359056 558278
rect 359004 558214 359056 558220
rect 358910 543416 358966 543425
rect 358910 543351 358966 543360
rect 358912 536920 358964 536926
rect 358912 536862 358964 536868
rect 358818 510096 358874 510105
rect 358818 510031 358874 510040
rect 358924 499458 358952 536862
rect 359016 513369 359044 558214
rect 359108 522345 359136 563790
rect 359188 555552 359240 555558
rect 359188 555494 359240 555500
rect 359094 522336 359150 522345
rect 359094 522271 359150 522280
rect 359200 520985 359228 555494
rect 359476 525842 359504 642262
rect 359568 536858 359596 642534
rect 360844 642388 360896 642394
rect 360844 642330 360896 642336
rect 359740 642184 359792 642190
rect 359740 642126 359792 642132
rect 359648 598596 359700 598602
rect 359648 598538 359700 598544
rect 359660 543794 359688 598538
rect 359648 543788 359700 543794
rect 359648 543730 359700 543736
rect 359556 536852 359608 536858
rect 359556 536794 359608 536800
rect 359648 535424 359700 535430
rect 359648 535366 359700 535372
rect 359464 525836 359516 525842
rect 359464 525778 359516 525784
rect 359554 524784 359610 524793
rect 359554 524719 359610 524728
rect 359186 520976 359242 520985
rect 359186 520911 359242 520920
rect 359002 513360 359058 513369
rect 359002 513295 359058 513304
rect 359464 511964 359516 511970
rect 359464 511906 359516 511912
rect 359280 505776 359332 505782
rect 359280 505718 359332 505724
rect 359292 500818 359320 505718
rect 359372 502988 359424 502994
rect 359372 502930 359424 502936
rect 359280 500812 359332 500818
rect 359280 500754 359332 500760
rect 358912 499452 358964 499458
rect 358912 499394 358964 499400
rect 359384 497865 359412 502930
rect 359370 497856 359426 497865
rect 359370 497791 359426 497800
rect 358544 175976 358596 175982
rect 358544 175918 358596 175924
rect 357808 89004 357860 89010
rect 357808 88946 357860 88952
rect 356796 20596 356848 20602
rect 356796 20538 356848 20544
rect 359476 6866 359504 511906
rect 359568 46918 359596 524719
rect 359660 245614 359688 535366
rect 359752 500857 359780 642126
rect 360016 641912 360068 641918
rect 360016 641854 360068 641860
rect 359832 640892 359884 640898
rect 359832 640834 359884 640840
rect 359844 598806 359872 640834
rect 360028 599593 360056 641854
rect 360108 639464 360160 639470
rect 360108 639406 360160 639412
rect 360014 599584 360070 599593
rect 360014 599519 360070 599528
rect 359832 598800 359884 598806
rect 359832 598742 359884 598748
rect 360120 552974 360148 639406
rect 360108 552968 360160 552974
rect 360108 552910 360160 552916
rect 360660 552696 360712 552702
rect 360660 552638 360712 552644
rect 360014 552120 360070 552129
rect 360014 552055 360070 552064
rect 360028 549916 360056 552055
rect 360672 549916 360700 552638
rect 360856 550798 360884 642330
rect 360948 599078 360976 642670
rect 370044 642660 370096 642666
rect 370044 642602 370096 642608
rect 368938 642152 368994 642161
rect 368938 642087 368994 642096
rect 366732 641844 366784 641850
rect 366732 641786 366784 641792
rect 363420 641776 363472 641782
rect 363420 641718 363472 641724
rect 361212 640416 361264 640422
rect 361212 640358 361264 640364
rect 361120 640348 361172 640354
rect 361120 640290 361172 640296
rect 360936 599072 360988 599078
rect 360936 599014 360988 599020
rect 361132 598738 361160 640290
rect 361224 598874 361252 640358
rect 363432 639948 363460 641718
rect 364524 640484 364576 640490
rect 364524 640426 364576 640432
rect 364536 639948 364564 640426
rect 365272 639946 365654 639962
rect 366744 639948 366772 641786
rect 367008 641776 367060 641782
rect 367008 641718 367060 641724
rect 364984 639940 365036 639946
rect 364984 639882 365036 639888
rect 365260 639940 365654 639946
rect 365312 639934 365654 639940
rect 365260 639882 365312 639888
rect 362224 639736 362276 639742
rect 362224 639678 362276 639684
rect 361488 639532 361540 639538
rect 361488 639474 361540 639480
rect 361212 598868 361264 598874
rect 361212 598810 361264 598816
rect 361120 598732 361172 598738
rect 361120 598674 361172 598680
rect 361028 598664 361080 598670
rect 361028 598606 361080 598612
rect 360936 598528 360988 598534
rect 360936 598470 360988 598476
rect 360948 551750 360976 598470
rect 360936 551744 360988 551750
rect 360936 551686 360988 551692
rect 361040 551274 361068 598606
rect 361120 585880 361172 585886
rect 361120 585822 361172 585828
rect 361132 552362 361160 585822
rect 361500 552702 361528 639474
rect 361946 639432 362002 639441
rect 361592 639390 361946 639418
rect 361592 638994 361620 639390
rect 362236 639402 362264 639678
rect 362498 639568 362554 639577
rect 362342 639526 362498 639554
rect 362498 639503 362554 639512
rect 362590 639432 362646 639441
rect 361946 639367 362002 639376
rect 362224 639396 362276 639402
rect 364062 639432 364118 639441
rect 362646 639390 362894 639418
rect 363998 639390 364062 639418
rect 362590 639367 362646 639376
rect 364996 639402 365024 639882
rect 367020 639878 367048 641718
rect 368952 639948 368980 642087
rect 369490 641744 369546 641753
rect 369490 641679 369546 641688
rect 369504 639948 369532 641679
rect 370056 639948 370084 642602
rect 376116 642592 376168 642598
rect 376116 642534 376168 642540
rect 371148 642456 371200 642462
rect 371148 642398 371200 642404
rect 371160 639948 371188 642398
rect 373356 642320 373408 642326
rect 373356 642262 373408 642268
rect 373908 642320 373960 642326
rect 373908 642262 373960 642268
rect 371700 641912 371752 641918
rect 371700 641854 371752 641860
rect 371712 639948 371740 641854
rect 372252 641776 372304 641782
rect 372252 641718 372304 641724
rect 372264 639948 372292 641718
rect 372804 640688 372856 640694
rect 372804 640630 372856 640636
rect 372816 639948 372844 640630
rect 373368 639948 373396 642262
rect 373920 639948 373948 642262
rect 375288 641912 375340 641918
rect 375288 641854 375340 641860
rect 367008 639872 367060 639878
rect 367008 639814 367060 639820
rect 375300 639810 375328 641854
rect 376128 639948 376156 642534
rect 377772 642524 377824 642530
rect 377772 642466 377824 642472
rect 377784 639948 377812 642466
rect 378048 641776 378100 641782
rect 378048 641718 378100 641724
rect 378060 641073 378088 641718
rect 378046 641064 378102 641073
rect 378046 640999 378102 641008
rect 378324 640824 378376 640830
rect 378324 640766 378376 640772
rect 378336 639948 378364 640766
rect 378874 640384 378930 640393
rect 378874 640319 378930 640328
rect 378888 639948 378916 640319
rect 379440 639948 379468 642670
rect 392676 642592 392728 642598
rect 392676 642534 392728 642540
rect 400772 642592 400824 642598
rect 400772 642534 400824 642540
rect 389916 642524 389968 642530
rect 389916 642466 389968 642472
rect 388260 642252 388312 642258
rect 388260 642194 388312 642200
rect 386604 642048 386656 642054
rect 386604 641990 386656 641996
rect 387708 642048 387760 642054
rect 387708 641990 387760 641996
rect 382186 641880 382242 641889
rect 379520 641844 379572 641850
rect 382186 641815 382242 641824
rect 386052 641844 386104 641850
rect 379520 641786 379572 641792
rect 379532 640937 379560 641786
rect 379518 640928 379574 640937
rect 379518 640863 379574 640872
rect 381636 640892 381688 640898
rect 381636 640834 381688 640840
rect 379980 640416 380032 640422
rect 379980 640358 380032 640364
rect 379992 639948 380020 640358
rect 381648 639948 381676 640834
rect 382200 639948 382228 641815
rect 386052 641786 386104 641792
rect 384396 641776 384448 641782
rect 384396 641718 384448 641724
rect 383844 640552 383896 640558
rect 383844 640494 383896 640500
rect 382740 640348 382792 640354
rect 382740 640290 382792 640296
rect 382752 639948 382780 640290
rect 383856 639948 383884 640494
rect 384408 639948 384436 641718
rect 384948 640756 385000 640762
rect 384948 640698 385000 640704
rect 384960 639948 384988 640698
rect 385500 640620 385552 640626
rect 385500 640562 385552 640568
rect 385512 639948 385540 640562
rect 386064 639948 386092 641786
rect 386616 639948 386644 641990
rect 387156 640552 387208 640558
rect 387156 640494 387208 640500
rect 387168 639948 387196 640494
rect 387720 639948 387748 641990
rect 388272 639948 388300 642194
rect 388812 642116 388864 642122
rect 388812 642058 388864 642064
rect 388824 639948 388852 642058
rect 389364 641912 389416 641918
rect 389364 641854 389416 641860
rect 389376 639948 389404 641854
rect 389928 639948 389956 642466
rect 390468 642184 390520 642190
rect 390468 642126 390520 642132
rect 390480 639948 390508 642126
rect 392124 642116 392176 642122
rect 392124 642058 392176 642064
rect 391020 641980 391072 641986
rect 391020 641922 391072 641928
rect 391032 639948 391060 641922
rect 392136 639948 392164 642058
rect 392688 639948 392716 642534
rect 399484 642524 399536 642530
rect 399484 642466 399536 642472
rect 396540 642388 396592 642394
rect 396540 642330 396592 642336
rect 394332 642252 394384 642258
rect 394332 642194 394384 642200
rect 393228 642184 393280 642190
rect 393228 642126 393280 642132
rect 393240 639948 393268 642126
rect 393780 641844 393832 641850
rect 393780 641786 393832 641792
rect 393792 639948 393820 641786
rect 394344 639948 394372 642194
rect 394884 641912 394936 641918
rect 394884 641854 394936 641860
rect 394896 639948 394924 641854
rect 395436 641776 395488 641782
rect 395436 641718 395488 641724
rect 395448 639948 395476 641718
rect 396552 639948 396580 642330
rect 398194 642288 398250 642297
rect 398194 642223 398250 642232
rect 397090 642016 397146 642025
rect 397090 641951 397146 641960
rect 397104 639948 397132 641951
rect 398208 641753 398236 642223
rect 399300 641844 399352 641850
rect 399300 641786 399352 641792
rect 398194 641744 398250 641753
rect 398194 641679 398250 641688
rect 399206 641744 399262 641753
rect 399206 641679 399262 641688
rect 398208 639948 398236 641679
rect 375288 639804 375340 639810
rect 375288 639746 375340 639752
rect 374644 639736 374696 639742
rect 367310 639674 367600 639690
rect 380162 639704 380218 639713
rect 374696 639684 375038 639690
rect 374644 639678 375038 639684
rect 367310 639668 367612 639674
rect 367310 639662 367560 639668
rect 367560 639610 367612 639616
rect 372528 639668 372580 639674
rect 374656 639662 375038 639678
rect 380218 639662 380558 639690
rect 399116 639668 399168 639674
rect 380162 639639 380218 639648
rect 372528 639610 372580 639616
rect 399116 639610 399168 639616
rect 370240 639538 370622 639554
rect 370228 639532 370622 639538
rect 370280 639526 370622 639532
rect 370228 639474 370280 639480
rect 368204 639464 368256 639470
rect 368110 639432 368166 639441
rect 365102 639402 365392 639418
rect 366206 639402 366496 639418
rect 364062 639367 364118 639376
rect 364984 639396 365036 639402
rect 362224 639338 362276 639344
rect 365102 639396 365404 639402
rect 365102 639390 365352 639396
rect 364984 639338 365036 639344
rect 366206 639396 366508 639402
rect 366206 639390 366456 639396
rect 365352 639338 365404 639344
rect 367862 639390 368110 639418
rect 369674 639432 369730 639441
rect 368256 639412 368414 639418
rect 368204 639406 368414 639412
rect 368216 639390 368414 639406
rect 372540 639402 372568 639610
rect 376300 639600 376352 639606
rect 396172 639600 396224 639606
rect 382922 639568 382978 639577
rect 376352 639548 376694 639554
rect 376300 639542 376694 639548
rect 376312 639526 376694 639542
rect 382978 639526 383318 639554
rect 396014 639548 396172 639554
rect 396014 639542 396224 639548
rect 399024 639600 399076 639606
rect 399024 639542 399076 639548
rect 391204 639532 391256 639538
rect 382922 639503 382978 639512
rect 396014 639526 396212 639542
rect 391204 639474 391256 639480
rect 374736 639464 374788 639470
rect 374486 639412 374736 639418
rect 377496 639464 377548 639470
rect 374486 639406 374788 639412
rect 368110 639367 368166 639376
rect 369674 639367 369676 639376
rect 366456 639338 366508 639344
rect 369728 639367 369730 639376
rect 372528 639396 372580 639402
rect 369676 639338 369728 639344
rect 374486 639390 374776 639406
rect 375590 639402 375880 639418
rect 377246 639412 377496 639418
rect 377246 639406 377548 639412
rect 380898 639432 380954 639441
rect 375590 639396 375892 639402
rect 375590 639390 375840 639396
rect 372528 639338 372580 639344
rect 377246 639390 377536 639406
rect 380954 639390 381110 639418
rect 391216 639402 391244 639474
rect 397920 639464 397972 639470
rect 391294 639432 391350 639441
rect 391204 639396 391256 639402
rect 380898 639367 380954 639376
rect 375840 639338 375892 639344
rect 391350 639390 391598 639418
rect 397670 639412 397920 639418
rect 397670 639406 397972 639412
rect 398932 639464 398984 639470
rect 398932 639406 398984 639412
rect 397670 639390 397960 639406
rect 391294 639367 391350 639376
rect 391204 639338 391256 639344
rect 361580 638988 361632 638994
rect 361580 638930 361632 638936
rect 398380 600296 398432 600302
rect 398380 600238 398432 600244
rect 398392 600114 398420 600238
rect 361776 599078 361804 600100
rect 361764 599072 361816 599078
rect 361764 599014 361816 599020
rect 361578 593192 361634 593201
rect 361578 593127 361634 593136
rect 361488 552696 361540 552702
rect 361488 552638 361540 552644
rect 361120 552356 361172 552362
rect 361120 552298 361172 552304
rect 361028 551268 361080 551274
rect 361028 551210 361080 551216
rect 360844 550792 360896 550798
rect 360844 550734 360896 550740
rect 361132 549930 361160 552298
rect 361592 549930 361620 593127
rect 361776 592034 361804 599014
rect 362328 593337 362356 600100
rect 362880 597582 362908 600100
rect 363432 598398 363460 600100
rect 363420 598392 363472 598398
rect 363420 598334 363472 598340
rect 362868 597576 362920 597582
rect 362868 597518 362920 597524
rect 363984 595542 364012 600100
rect 364352 600086 364550 600114
rect 364720 600086 365102 600114
rect 365272 600086 365654 600114
rect 363972 595536 364024 595542
rect 363972 595478 364024 595484
rect 362314 593328 362370 593337
rect 362314 593263 362370 593272
rect 361776 592006 361896 592034
rect 361868 551993 361896 592006
rect 362960 563712 363012 563718
rect 362960 563654 363012 563660
rect 362972 557534 363000 563654
rect 363236 559700 363288 559706
rect 363236 559642 363288 559648
rect 362972 557506 363184 557534
rect 362592 556844 362644 556850
rect 362592 556786 362644 556792
rect 361854 551984 361910 551993
rect 361854 551919 361910 551928
rect 362604 549930 362632 556786
rect 363156 551274 363184 557506
rect 363144 551268 363196 551274
rect 363144 551210 363196 551216
rect 362960 550044 363012 550050
rect 362960 549986 363012 549992
rect 361132 549902 361330 549930
rect 361592 549902 361974 549930
rect 362328 549916 362632 549930
rect 362972 549930 363000 549986
rect 363248 549930 363276 559642
rect 363604 551268 363656 551274
rect 363604 551210 363656 551216
rect 362972 549916 363276 549930
rect 363616 549930 363644 551210
rect 364352 551138 364380 600086
rect 364432 596080 364484 596086
rect 364432 596022 364484 596028
rect 364444 559638 364472 596022
rect 364720 590034 364748 600086
rect 365272 596086 365300 600086
rect 365720 599616 365772 599622
rect 365720 599558 365772 599564
rect 365260 596080 365312 596086
rect 365260 596022 365312 596028
rect 364708 590028 364760 590034
rect 364708 589970 364760 589976
rect 364522 581632 364578 581641
rect 364522 581567 364578 581576
rect 364432 559632 364484 559638
rect 364432 559574 364484 559580
rect 364340 551132 364392 551138
rect 364340 551074 364392 551080
rect 364352 550662 364380 551074
rect 364340 550656 364392 550662
rect 364340 550598 364392 550604
rect 362328 549902 362618 549916
rect 362972 549902 363262 549916
rect 363616 549902 363906 549930
rect 364536 549916 364564 581567
rect 365168 551132 365220 551138
rect 365168 551074 365220 551080
rect 365180 549916 365208 551074
rect 365732 549930 365760 599558
rect 366192 598466 366220 600100
rect 366284 600086 366758 600114
rect 366180 598460 366232 598466
rect 366180 598402 366232 598408
rect 366284 586514 366312 600086
rect 367296 596426 367324 600100
rect 367388 600086 367862 600114
rect 368032 600086 368414 600114
rect 368492 600086 368966 600114
rect 369044 600086 369518 600114
rect 369964 600086 370070 600114
rect 370240 600086 370622 600114
rect 370792 600086 371174 600114
rect 371252 600086 371726 600114
rect 371804 600086 372278 600114
rect 367284 596420 367336 596426
rect 367284 596362 367336 596368
rect 367284 596216 367336 596222
rect 367284 596158 367336 596164
rect 367100 596080 367152 596086
rect 367100 596022 367152 596028
rect 365824 586486 366312 586514
rect 365824 556238 365852 586486
rect 365904 565208 365956 565214
rect 365904 565150 365956 565156
rect 365916 557534 365944 565150
rect 365916 557506 366128 557534
rect 365812 556232 365864 556238
rect 365812 556174 365864 556180
rect 366100 549930 366128 557506
rect 367112 554810 367140 596022
rect 367192 589484 367244 589490
rect 367192 589426 367244 589432
rect 367204 588674 367232 589426
rect 367192 588668 367244 588674
rect 367192 588610 367244 588616
rect 367192 581664 367244 581670
rect 367192 581606 367244 581612
rect 367204 557534 367232 581606
rect 367296 568585 367324 596158
rect 367388 589490 367416 600086
rect 368032 596086 368060 600086
rect 368020 596080 368072 596086
rect 368020 596022 368072 596028
rect 367376 589484 367428 589490
rect 367376 589426 367428 589432
rect 367376 573436 367428 573442
rect 367376 573378 367428 573384
rect 367282 568576 367338 568585
rect 367282 568511 367338 568520
rect 367388 557534 367416 573378
rect 367204 557506 367324 557534
rect 367388 557506 367968 557534
rect 367100 554804 367152 554810
rect 367100 554746 367152 554752
rect 367112 554266 367140 554746
rect 367100 554260 367152 554266
rect 367100 554202 367152 554208
rect 367296 553394 367324 557506
rect 367296 553366 367416 553394
rect 367100 550792 367152 550798
rect 367100 550734 367152 550740
rect 365732 549902 365838 549930
rect 366100 549902 366482 549930
rect 367112 549916 367140 550734
rect 367388 549930 367416 553366
rect 367940 549930 367968 557506
rect 368492 551721 368520 600086
rect 369044 597666 369072 600086
rect 369860 598188 369912 598194
rect 369860 598130 369912 598136
rect 368584 597638 369072 597666
rect 368584 587246 368612 597638
rect 368664 597576 368716 597582
rect 368664 597518 368716 597524
rect 368572 587240 368624 587246
rect 368572 587182 368624 587188
rect 368572 567928 368624 567934
rect 368572 567870 368624 567876
rect 368478 551712 368534 551721
rect 368478 551647 368534 551656
rect 368584 551018 368612 567870
rect 368676 552906 368704 597518
rect 369872 554169 369900 598130
rect 369964 554878 369992 600086
rect 370240 598194 370268 600086
rect 370228 598188 370280 598194
rect 370228 598130 370280 598136
rect 370792 586514 370820 600086
rect 370056 586486 370820 586514
rect 370056 563145 370084 586486
rect 370134 565040 370190 565049
rect 370134 564975 370190 564984
rect 370042 563136 370098 563145
rect 370042 563071 370098 563080
rect 370148 563054 370176 564975
rect 370148 563026 370544 563054
rect 369952 554872 370004 554878
rect 369952 554814 370004 554820
rect 369964 554198 369992 554814
rect 369952 554192 370004 554198
rect 369858 554160 369914 554169
rect 369952 554134 370004 554140
rect 369858 554095 369914 554104
rect 368664 552900 368716 552906
rect 368664 552842 368716 552848
rect 368584 550990 369256 551018
rect 369032 550656 369084 550662
rect 369032 550598 369084 550604
rect 367388 549902 367770 549930
rect 367940 549902 368414 549930
rect 369044 549916 369072 550598
rect 369228 549930 369256 550990
rect 370516 549930 370544 563026
rect 371252 555529 371280 600086
rect 371804 594182 371832 600086
rect 372620 599684 372672 599690
rect 372620 599626 372672 599632
rect 371792 594176 371844 594182
rect 371792 594118 371844 594124
rect 371884 594108 371936 594114
rect 371884 594050 371936 594056
rect 371332 556232 371384 556238
rect 371332 556174 371384 556180
rect 371238 555520 371294 555529
rect 371238 555455 371294 555464
rect 371344 549930 371372 556174
rect 371896 552158 371924 594050
rect 371884 552152 371936 552158
rect 371884 552094 371936 552100
rect 371896 549930 371924 552094
rect 372632 549930 372660 599626
rect 372712 598188 372764 598194
rect 372712 598130 372764 598136
rect 372724 565894 372752 598130
rect 372816 585818 372844 600100
rect 372908 600086 373382 600114
rect 373552 600086 373934 600114
rect 374012 600086 374486 600114
rect 374656 600086 375038 600114
rect 372908 595542 372936 600086
rect 373552 598194 373580 600086
rect 373540 598188 373592 598194
rect 373540 598130 373592 598136
rect 372896 595536 372948 595542
rect 372896 595478 372948 595484
rect 372804 585812 372856 585818
rect 372804 585754 372856 585760
rect 372712 565888 372764 565894
rect 372712 565830 372764 565836
rect 372724 565282 372752 565830
rect 372712 565276 372764 565282
rect 372712 565218 372764 565224
rect 374012 556850 374040 600086
rect 374656 586514 374684 600086
rect 375576 596970 375604 600100
rect 376128 597689 376156 600100
rect 376220 600086 376694 600114
rect 376772 600086 377246 600114
rect 377416 600086 377798 600114
rect 378244 600086 378350 600114
rect 378428 600086 378902 600114
rect 379072 600086 379454 600114
rect 379624 600086 380006 600114
rect 376114 597680 376170 597689
rect 376114 597615 376170 597624
rect 375564 596964 375616 596970
rect 375564 596906 375616 596912
rect 376220 586514 376248 600086
rect 374104 586486 374684 586514
rect 375668 586486 376248 586514
rect 374104 559706 374132 586486
rect 374276 570716 374328 570722
rect 374276 570658 374328 570664
rect 374288 563054 374316 570658
rect 374288 563026 374408 563054
rect 374092 559700 374144 559706
rect 374092 559642 374144 559648
rect 374000 556844 374052 556850
rect 374000 556786 374052 556792
rect 374184 552696 374236 552702
rect 374184 552638 374236 552644
rect 373540 552152 373592 552158
rect 373540 552094 373592 552100
rect 369228 549902 369702 549930
rect 370516 549902 370990 549930
rect 371344 549902 371634 549930
rect 371896 549902 372278 549930
rect 372632 549902 372922 549930
rect 373552 549916 373580 552094
rect 374196 549916 374224 552638
rect 374380 549930 374408 563026
rect 375472 558204 375524 558210
rect 375472 558146 375524 558152
rect 375012 551948 375064 551954
rect 375012 551890 375064 551896
rect 375024 550118 375052 551890
rect 375012 550112 375064 550118
rect 375012 550054 375064 550060
rect 374380 549902 374854 549930
rect 375484 549916 375512 558146
rect 375668 552362 375696 586486
rect 376668 559632 376720 559638
rect 376668 559574 376720 559580
rect 376116 552696 376168 552702
rect 376116 552638 376168 552644
rect 375656 552356 375708 552362
rect 375656 552298 375708 552304
rect 375668 551954 375696 552298
rect 375656 551948 375708 551954
rect 375656 551890 375708 551896
rect 376128 549916 376156 552638
rect 376680 551614 376708 559574
rect 376772 558210 376800 600086
rect 377416 586514 377444 600086
rect 376956 586486 377444 586514
rect 376852 566500 376904 566506
rect 376852 566442 376904 566448
rect 376864 563054 376892 566442
rect 376956 565865 376984 586486
rect 376942 565856 376998 565865
rect 376942 565791 376998 565800
rect 376864 563026 376984 563054
rect 376760 558204 376812 558210
rect 376760 558146 376812 558152
rect 376758 552664 376814 552673
rect 376758 552599 376814 552608
rect 376668 551608 376720 551614
rect 376668 551550 376720 551556
rect 376772 549916 376800 552599
rect 376956 549930 376984 563026
rect 378244 558385 378272 600086
rect 378428 598346 378456 600086
rect 378508 599752 378560 599758
rect 378508 599694 378560 599700
rect 378336 598318 378456 598346
rect 378336 562465 378364 598318
rect 378416 598188 378468 598194
rect 378416 598130 378468 598136
rect 378428 571985 378456 598130
rect 378414 571976 378470 571985
rect 378414 571911 378470 571920
rect 378520 563054 378548 599694
rect 379072 598194 379100 600086
rect 379060 598188 379112 598194
rect 379060 598130 379112 598136
rect 379624 577561 379652 600086
rect 380544 598670 380572 600100
rect 381110 600086 381216 600114
rect 380532 598664 380584 598670
rect 380532 598606 380584 598612
rect 380992 598188 381044 598194
rect 380992 598130 381044 598136
rect 379610 577552 379666 577561
rect 379520 577516 379572 577522
rect 379610 577487 379666 577496
rect 379520 577458 379572 577464
rect 378520 563026 379008 563054
rect 378322 562456 378378 562465
rect 378322 562391 378378 562400
rect 378230 558376 378286 558385
rect 378230 558311 378286 558320
rect 377128 558204 377180 558210
rect 377128 558146 377180 558152
rect 377140 551682 377168 558146
rect 378048 556844 378100 556850
rect 378048 556786 378100 556792
rect 377128 551676 377180 551682
rect 377128 551618 377180 551624
rect 376956 549902 377430 549930
rect 378060 549916 378088 556786
rect 378692 552968 378744 552974
rect 378692 552910 378744 552916
rect 378704 549916 378732 552910
rect 378784 549976 378836 549982
rect 378784 549918 378836 549924
rect 378980 549930 379008 563026
rect 379532 557534 379560 577458
rect 381004 558278 381032 598130
rect 381084 562352 381136 562358
rect 381084 562294 381136 562300
rect 380992 558272 381044 558278
rect 380992 558214 381044 558220
rect 379532 557506 380296 557534
rect 379980 552832 380032 552838
rect 379980 552774 380032 552780
rect 362328 549846 362356 549902
rect 371344 549846 371372 549902
rect 378796 549846 378824 549918
rect 378980 549902 379362 549930
rect 379992 549916 380020 552774
rect 380164 550112 380216 550118
rect 380164 550054 380216 550060
rect 380176 549914 380204 550054
rect 380268 549930 380296 557506
rect 380992 549976 381044 549982
rect 380164 549908 380216 549914
rect 380268 549902 380650 549930
rect 380992 549918 381044 549924
rect 381096 549930 381124 562294
rect 381188 556918 381216 600086
rect 381280 600086 381662 600114
rect 381280 598194 381308 600086
rect 382200 598602 382228 600100
rect 382384 600086 382766 600114
rect 382280 599820 382332 599826
rect 382280 599762 382332 599768
rect 382188 598596 382240 598602
rect 382188 598538 382240 598544
rect 381268 598188 381320 598194
rect 381268 598130 381320 598136
rect 381544 590028 381596 590034
rect 381544 589970 381596 589976
rect 381176 556912 381228 556918
rect 381176 556854 381228 556860
rect 381556 552090 381584 589970
rect 381544 552084 381596 552090
rect 381544 552026 381596 552032
rect 381556 549930 381584 552026
rect 382292 551274 382320 599762
rect 382384 563689 382412 600086
rect 383304 598233 383332 600100
rect 383764 600086 383870 600114
rect 383948 600086 384422 600114
rect 384592 600086 384974 600114
rect 385052 600086 385526 600114
rect 385604 600086 386078 600114
rect 386524 600086 386630 600114
rect 383290 598224 383346 598233
rect 383290 598159 383346 598168
rect 383660 597236 383712 597242
rect 383660 597178 383712 597184
rect 382464 578944 382516 578950
rect 382464 578886 382516 578892
rect 382370 563680 382426 563689
rect 382370 563615 382426 563624
rect 382280 551268 382332 551274
rect 382280 551210 382332 551216
rect 382476 549930 382504 578886
rect 383672 551614 383700 597178
rect 383764 552974 383792 600086
rect 383844 595536 383896 595542
rect 383844 595478 383896 595484
rect 383752 552968 383804 552974
rect 383752 552910 383804 552916
rect 383660 551608 383712 551614
rect 383660 551550 383712 551556
rect 382924 551268 382976 551274
rect 382924 551210 382976 551216
rect 382936 549930 382964 551210
rect 383856 549930 383884 595478
rect 383948 595270 383976 600086
rect 384592 597242 384620 600086
rect 384580 597236 384632 597242
rect 384580 597178 384632 597184
rect 383936 595264 383988 595270
rect 383936 595206 383988 595212
rect 384304 560788 384356 560794
rect 384304 560730 384356 560736
rect 384316 552226 384344 560730
rect 385052 553314 385080 600086
rect 385604 586514 385632 600086
rect 386420 598868 386472 598874
rect 386420 598810 386472 598816
rect 385684 592068 385736 592074
rect 385684 592010 385736 592016
rect 385144 586486 385632 586514
rect 385144 555558 385172 586486
rect 385132 555552 385184 555558
rect 385132 555494 385184 555500
rect 385040 553308 385092 553314
rect 385040 553250 385092 553256
rect 385696 552294 385724 592010
rect 386432 590034 386460 598810
rect 386420 590028 386472 590034
rect 386420 589970 386472 589976
rect 386524 563854 386552 600086
rect 386604 599004 386656 599010
rect 386604 598946 386656 598952
rect 386616 581641 386644 598946
rect 387168 598874 387196 600100
rect 387720 599146 387748 600100
rect 387708 599140 387760 599146
rect 387708 599082 387760 599088
rect 387720 599010 387748 599082
rect 387708 599004 387760 599010
rect 387708 598946 387760 598952
rect 388272 598942 388300 600100
rect 388456 600086 388838 600114
rect 389390 600086 389496 600114
rect 388260 598936 388312 598942
rect 388260 598878 388312 598884
rect 387156 598868 387208 598874
rect 387156 598810 387208 598816
rect 388272 598602 388300 598878
rect 388456 598806 388484 600086
rect 388444 598800 388496 598806
rect 388444 598742 388496 598748
rect 388260 598596 388312 598602
rect 388260 598538 388312 598544
rect 386788 589960 386840 589966
rect 386788 589902 386840 589908
rect 386602 581632 386658 581641
rect 386602 581567 386658 581576
rect 386604 570648 386656 570654
rect 386604 570590 386656 570596
rect 386512 563848 386564 563854
rect 386512 563790 386564 563796
rect 385684 552288 385736 552294
rect 385684 552230 385736 552236
rect 384304 552220 384356 552226
rect 384304 552162 384356 552168
rect 383936 550112 383988 550118
rect 383936 550054 383988 550060
rect 380164 549850 380216 549856
rect 381004 549846 381032 549918
rect 381096 549902 381294 549930
rect 381556 549902 381938 549930
rect 382476 549902 382582 549930
rect 382936 549902 383226 549930
rect 383580 549916 383884 549930
rect 383580 549914 383870 549916
rect 383948 549914 383976 550054
rect 384316 549930 384344 552162
rect 385696 549930 385724 552230
rect 386616 550594 386644 570590
rect 386696 567860 386748 567866
rect 386696 567802 386748 567808
rect 386604 550588 386656 550594
rect 386604 550530 386656 550536
rect 386708 549930 386736 567802
rect 386800 557534 386828 589902
rect 388456 564505 388484 598742
rect 388536 598596 388588 598602
rect 388536 598538 388588 598544
rect 388548 569401 388576 598538
rect 389272 598188 389324 598194
rect 389272 598130 389324 598136
rect 389180 598120 389232 598126
rect 389180 598062 389232 598068
rect 389192 592074 389220 598062
rect 389180 592068 389232 592074
rect 389180 592010 389232 592016
rect 389284 579601 389312 598130
rect 389270 579592 389326 579601
rect 389270 579527 389326 579536
rect 389272 576156 389324 576162
rect 389272 576098 389324 576104
rect 388534 569392 388590 569401
rect 388534 569327 388590 569336
rect 388536 567248 388588 567254
rect 388536 567190 388588 567196
rect 388442 564496 388498 564505
rect 388442 564431 388498 564440
rect 386800 557506 387288 557534
rect 387064 550588 387116 550594
rect 387064 550530 387116 550536
rect 383568 549908 383870 549914
rect 383620 549902 383870 549908
rect 383936 549908 383988 549914
rect 383568 549850 383620 549856
rect 384316 549902 384514 549930
rect 385696 549902 385802 549930
rect 386446 549902 386736 549930
rect 387076 549916 387104 550530
rect 387260 549930 387288 557506
rect 388352 552900 388404 552906
rect 388352 552842 388404 552848
rect 387260 549902 387734 549930
rect 388364 549916 388392 552842
rect 388548 550866 388576 567190
rect 389284 557534 389312 576098
rect 389284 557506 389404 557534
rect 389272 553104 389324 553110
rect 389272 553046 389324 553052
rect 388536 550860 388588 550866
rect 388536 550802 388588 550808
rect 388996 550860 389048 550866
rect 388996 550802 389048 550808
rect 389008 549916 389036 550802
rect 389284 549930 389312 553046
rect 389376 550066 389404 557506
rect 389468 551750 389496 600086
rect 389560 600086 389942 600114
rect 390112 600086 390494 600114
rect 390756 600086 391046 600114
rect 389560 598194 389588 600086
rect 389548 598188 389600 598194
rect 389548 598130 389600 598136
rect 390112 598126 390140 600086
rect 390100 598120 390152 598126
rect 390100 598062 390152 598068
rect 390652 573368 390704 573374
rect 390652 573310 390704 573316
rect 389456 551744 389508 551750
rect 389456 551686 389508 551692
rect 389376 550038 389864 550066
rect 389836 549930 389864 550038
rect 390664 549930 390692 573310
rect 390756 560794 390784 600086
rect 391584 598534 391612 600100
rect 392044 600086 392150 600114
rect 392320 600086 392702 600114
rect 392872 600086 393254 600114
rect 393424 600086 393806 600114
rect 393976 600086 394358 600114
rect 394712 600086 394910 600114
rect 391940 600024 391992 600030
rect 391940 599966 391992 599972
rect 391572 598528 391624 598534
rect 391572 598470 391624 598476
rect 391202 595504 391258 595513
rect 391202 595439 391258 595448
rect 390744 560788 390796 560794
rect 390744 560730 390796 560736
rect 391216 552090 391244 595439
rect 391952 594114 391980 599966
rect 392044 598210 392072 600086
rect 392320 600030 392348 600086
rect 392308 600024 392360 600030
rect 392308 599966 392360 599972
rect 392308 599888 392360 599894
rect 392308 599830 392360 599836
rect 392044 598182 392164 598210
rect 392032 598120 392084 598126
rect 392032 598062 392084 598068
rect 391940 594108 391992 594114
rect 391940 594050 391992 594056
rect 392044 563689 392072 598062
rect 392136 585886 392164 598182
rect 392124 585880 392176 585886
rect 392124 585822 392176 585828
rect 392030 563680 392086 563689
rect 392030 563615 392086 563624
rect 392320 557534 392348 599830
rect 392872 598126 392900 600086
rect 393320 598188 393372 598194
rect 393320 598130 393372 598136
rect 392860 598120 392912 598126
rect 392860 598062 392912 598068
rect 392584 595264 392636 595270
rect 392584 595206 392636 595212
rect 392320 557506 392440 557534
rect 392216 553308 392268 553314
rect 392216 553250 392268 553256
rect 391204 552084 391256 552090
rect 391204 552026 391256 552032
rect 391572 552084 391624 552090
rect 391572 552026 391624 552032
rect 389284 549902 389666 549930
rect 389836 549902 390310 549930
rect 390664 549902 390954 549930
rect 391584 549916 391612 552026
rect 392228 549916 392256 553250
rect 392412 549930 392440 557506
rect 392596 553382 392624 595206
rect 392584 553376 392636 553382
rect 392584 553318 392636 553324
rect 393332 550526 393360 598130
rect 393424 567254 393452 600086
rect 393976 598194 394004 600086
rect 393964 598188 394016 598194
rect 393964 598130 394016 598136
rect 393412 567248 393464 567254
rect 393412 567190 393464 567196
rect 394712 563786 394740 600086
rect 395448 597854 395476 600100
rect 395540 600086 396014 600114
rect 396184 600086 396566 600114
rect 396736 600086 397118 600114
rect 397564 600086 397670 600114
rect 398222 600100 398420 600114
rect 398208 600086 398420 600100
rect 395436 597848 395488 597854
rect 395436 597790 395488 597796
rect 395540 586514 395568 600086
rect 396080 598188 396132 598194
rect 396080 598130 396132 598136
rect 394804 586486 395568 586514
rect 394804 575521 394832 586486
rect 394790 575512 394846 575521
rect 394790 575447 394846 575456
rect 394884 574796 394936 574802
rect 394884 574738 394936 574744
rect 394700 563780 394752 563786
rect 394700 563722 394752 563728
rect 394896 557534 394924 574738
rect 396092 565146 396120 598130
rect 396184 591394 396212 600086
rect 396736 598194 396764 600086
rect 396724 598188 396776 598194
rect 396724 598130 396776 598136
rect 396172 591388 396224 591394
rect 396172 591330 396224 591336
rect 397458 581768 397514 581777
rect 397458 581703 397514 581712
rect 396172 574864 396224 574870
rect 396172 574806 396224 574812
rect 396080 565140 396132 565146
rect 396080 565082 396132 565088
rect 396080 559632 396132 559638
rect 396080 559574 396132 559580
rect 394896 557506 395016 557534
rect 394148 553376 394200 553382
rect 394148 553318 394200 553324
rect 393504 552560 393556 552566
rect 393504 552502 393556 552508
rect 393320 550520 393372 550526
rect 393320 550462 393372 550468
rect 392412 549902 392886 549930
rect 393516 549916 393544 552502
rect 394160 549916 394188 553318
rect 394792 552220 394844 552226
rect 394792 552162 394844 552168
rect 394804 549916 394832 552162
rect 394988 549930 395016 557506
rect 394988 549902 395462 549930
rect 396092 549916 396120 559574
rect 396184 557534 396212 574806
rect 396184 557506 397040 557534
rect 396724 552764 396776 552770
rect 396724 552706 396776 552712
rect 396736 549916 396764 552706
rect 397012 549930 397040 557506
rect 397472 549930 397500 581703
rect 397564 550050 397592 600086
rect 397736 598460 397788 598466
rect 397736 598402 397788 598408
rect 397748 557534 397776 598402
rect 398104 598392 398156 598398
rect 398104 598334 398156 598340
rect 397656 557506 397776 557534
rect 397656 550118 397684 557506
rect 398116 552022 398144 598334
rect 398208 596834 398236 600086
rect 398196 596828 398248 596834
rect 398196 596770 398248 596776
rect 398656 552288 398708 552294
rect 398656 552230 398708 552236
rect 398104 552016 398156 552022
rect 398104 551958 398156 551964
rect 397644 550112 397696 550118
rect 397642 550080 397644 550089
rect 397696 550080 397698 550089
rect 397552 550044 397604 550050
rect 397642 550015 397698 550024
rect 397552 549986 397604 549992
rect 397012 549902 397394 549930
rect 397472 549902 398038 549930
rect 398668 549916 398696 552230
rect 398944 549930 398972 639406
rect 399036 552702 399064 639542
rect 399128 553110 399156 639610
rect 399220 599894 399248 641679
rect 399208 599888 399260 599894
rect 399208 599830 399260 599836
rect 399312 599690 399340 641786
rect 399300 599684 399352 599690
rect 399300 599626 399352 599632
rect 399116 553104 399168 553110
rect 399116 553046 399168 553052
rect 399496 552702 399524 642466
rect 400680 642184 400732 642190
rect 400680 642126 400732 642132
rect 400404 642116 400456 642122
rect 400404 642058 400456 642064
rect 399576 642048 399628 642054
rect 399576 641990 399628 641996
rect 399024 552696 399076 552702
rect 399024 552638 399076 552644
rect 399484 552696 399536 552702
rect 399484 552638 399536 552644
rect 399484 551608 399536 551614
rect 399484 551550 399536 551556
rect 398944 549902 399326 549930
rect 383936 549850 383988 549856
rect 359924 549840 359976 549846
rect 359924 549782 359976 549788
rect 362316 549840 362368 549846
rect 362316 549782 362368 549788
rect 371332 549840 371384 549846
rect 371332 549782 371384 549788
rect 378784 549840 378836 549846
rect 378784 549782 378836 549788
rect 380992 549840 381044 549846
rect 380992 549782 381044 549788
rect 359832 549704 359884 549710
rect 359832 549646 359884 549652
rect 359844 549370 359872 549646
rect 359936 549438 359964 549782
rect 359924 549432 359976 549438
rect 359924 549374 359976 549380
rect 359832 549364 359884 549370
rect 359832 549306 359884 549312
rect 359832 514344 359884 514350
rect 359832 514286 359884 514292
rect 359738 500848 359794 500857
rect 359738 500783 359794 500792
rect 359740 500336 359792 500342
rect 359740 500278 359792 500284
rect 359752 499934 359780 500278
rect 359740 499928 359792 499934
rect 359740 499870 359792 499876
rect 359844 458182 359872 514286
rect 399496 507385 399524 551550
rect 399588 546514 399616 641990
rect 399668 641776 399720 641782
rect 399668 641718 399720 641724
rect 399680 550594 399708 641718
rect 400312 640688 400364 640694
rect 400312 640630 400364 640636
rect 400220 640484 400272 640490
rect 400220 640426 400272 640432
rect 399944 639260 399996 639266
rect 399944 639202 399996 639208
rect 399852 555484 399904 555490
rect 399852 555426 399904 555432
rect 399760 551744 399812 551750
rect 399760 551686 399812 551692
rect 399668 550588 399720 550594
rect 399668 550530 399720 550536
rect 399576 546508 399628 546514
rect 399576 546450 399628 546456
rect 399772 537033 399800 551686
rect 399758 537024 399814 537033
rect 399758 536959 399814 536968
rect 399864 536625 399892 555426
rect 399850 536616 399906 536625
rect 399850 536551 399906 536560
rect 399574 536344 399630 536353
rect 399574 536279 399630 536288
rect 399482 507376 399538 507385
rect 399482 507311 399538 507320
rect 399482 501664 399538 501673
rect 399482 501599 399538 501608
rect 359924 500812 359976 500818
rect 359924 500754 359976 500760
rect 359936 498982 359964 500754
rect 360028 499769 360056 500140
rect 360476 499996 360528 500002
rect 360476 499938 360528 499944
rect 360014 499760 360070 499769
rect 360014 499695 360070 499704
rect 359924 498976 359976 498982
rect 359924 498918 359976 498924
rect 360488 497729 360516 499938
rect 360672 499905 360700 500140
rect 360658 499896 360714 499905
rect 360658 499831 360714 499840
rect 361316 498098 361344 500140
rect 361960 498166 361988 500140
rect 361948 498160 362000 498166
rect 361948 498102 362000 498108
rect 361304 498092 361356 498098
rect 361304 498034 361356 498040
rect 360474 497720 360530 497729
rect 360474 497655 360530 497664
rect 362604 497457 362632 500140
rect 362960 499928 363012 499934
rect 362958 499896 362960 499905
rect 363012 499896 363014 499905
rect 362958 499831 363014 499840
rect 362590 497448 362646 497457
rect 362590 497383 362646 497392
rect 363248 497282 363276 500140
rect 363892 499934 363920 500140
rect 363880 499928 363932 499934
rect 363880 499870 363932 499876
rect 364536 498030 364564 500140
rect 365180 499905 365208 500140
rect 365166 499896 365222 499905
rect 365166 499831 365222 499840
rect 365824 499497 365852 500140
rect 365810 499488 365866 499497
rect 365810 499423 365866 499432
rect 364524 498024 364576 498030
rect 364524 497966 364576 497972
rect 366468 497554 366496 500140
rect 367112 498914 367140 500140
rect 367756 499497 367784 500140
rect 368400 499905 368428 500140
rect 368386 499896 368442 499905
rect 368386 499831 368442 499840
rect 367742 499488 367798 499497
rect 367742 499423 367798 499432
rect 367100 498908 367152 498914
rect 367100 498850 367152 498856
rect 367756 498846 367784 499423
rect 367744 498840 367796 498846
rect 367744 498782 367796 498788
rect 369044 498137 369072 500140
rect 369688 499390 369716 500140
rect 369676 499384 369728 499390
rect 369676 499326 369728 499332
rect 370332 498778 370360 500140
rect 370976 499905 371004 500140
rect 371620 499905 371648 500140
rect 370962 499896 371018 499905
rect 370962 499831 371018 499840
rect 371606 499896 371662 499905
rect 371606 499831 371662 499840
rect 370320 498772 370372 498778
rect 370320 498714 370372 498720
rect 369030 498128 369086 498137
rect 369030 498063 369086 498072
rect 366456 497548 366508 497554
rect 366456 497490 366508 497496
rect 369044 497321 369072 498063
rect 371620 497690 371648 499831
rect 371608 497684 371660 497690
rect 371608 497626 371660 497632
rect 372264 497350 372292 500140
rect 372252 497344 372304 497350
rect 369030 497312 369086 497321
rect 363236 497276 363288 497282
rect 372252 497286 372304 497292
rect 369030 497247 369086 497256
rect 363236 497218 363288 497224
rect 362224 496392 362276 496398
rect 362224 496334 362276 496340
rect 359832 458176 359884 458182
rect 359832 458118 359884 458124
rect 362236 353258 362264 496334
rect 364340 480956 364392 480962
rect 364340 480898 364392 480904
rect 363604 475380 363656 475386
rect 363604 475322 363656 475328
rect 362224 353252 362276 353258
rect 362224 353194 362276 353200
rect 359648 245608 359700 245614
rect 359648 245550 359700 245556
rect 363616 117298 363644 475322
rect 363604 117292 363656 117298
rect 363604 117234 363656 117240
rect 359556 46912 359608 46918
rect 359556 46854 359608 46860
rect 364352 16574 364380 480898
rect 371240 478168 371292 478174
rect 371240 478110 371292 478116
rect 364352 16546 364656 16574
rect 359464 6860 359516 6866
rect 359464 6802 359516 6808
rect 357532 4888 357584 4894
rect 357532 4830 357584 4836
rect 355416 4072 355468 4078
rect 355416 4014 355468 4020
rect 355324 3868 355376 3874
rect 355324 3810 355376 3816
rect 353484 3324 353536 3330
rect 353484 3266 353536 3272
rect 353392 3256 353444 3262
rect 353392 3198 353444 3204
rect 357544 480 357572 4830
rect 361120 3868 361172 3874
rect 361120 3810 361172 3816
rect 361132 480 361160 3810
rect 364628 480 364656 16546
rect 367744 14544 367796 14550
rect 367744 14486 367796 14492
rect 354006 354 354118 480
rect 353312 326 354118 354
rect 354006 -960 354118 326
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 14486
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371252 354 371280 478110
rect 372908 126954 372936 500140
rect 373552 499390 373580 500140
rect 373540 499384 373592 499390
rect 374840 499361 374868 500140
rect 373540 499326 373592 499332
rect 374826 499352 374882 499361
rect 374826 499287 374882 499296
rect 375484 498778 375512 500140
rect 375472 498772 375524 498778
rect 375472 498714 375524 498720
rect 376128 498137 376156 500140
rect 376390 499896 376446 499905
rect 376390 499831 376446 499840
rect 376114 498128 376170 498137
rect 376114 498063 376170 498072
rect 376128 497826 376156 498063
rect 376404 497826 376432 499831
rect 376772 499497 376800 500140
rect 377416 499905 377444 500140
rect 377402 499896 377458 499905
rect 377402 499831 377458 499840
rect 376758 499488 376814 499497
rect 376758 499423 376814 499432
rect 376116 497820 376168 497826
rect 376116 497762 376168 497768
rect 376392 497820 376444 497826
rect 376392 497762 376444 497768
rect 378060 497758 378088 500140
rect 378048 497752 378100 497758
rect 378048 497694 378100 497700
rect 374000 496120 374052 496126
rect 374000 496062 374052 496068
rect 372896 126948 372948 126954
rect 372896 126890 372948 126896
rect 374012 3398 374040 496062
rect 376024 494760 376076 494766
rect 376024 494702 376076 494708
rect 376036 405686 376064 494702
rect 378704 493474 378732 500140
rect 379348 499526 379376 500140
rect 379336 499520 379388 499526
rect 379336 499462 379388 499468
rect 379992 497894 380020 500140
rect 380636 499905 380664 500140
rect 381280 499905 381308 500140
rect 380622 499896 380678 499905
rect 380622 499831 380678 499840
rect 381266 499896 381322 499905
rect 381266 499831 381322 499840
rect 381924 498982 381952 500140
rect 382568 499905 382596 500140
rect 382554 499896 382610 499905
rect 382554 499831 382610 499840
rect 381912 498976 381964 498982
rect 381912 498918 381964 498924
rect 379980 497888 380032 497894
rect 379980 497830 380032 497836
rect 382568 497185 382596 499831
rect 382554 497176 382610 497185
rect 382554 497111 382610 497120
rect 378692 493468 378744 493474
rect 378692 493410 378744 493416
rect 376024 405680 376076 405686
rect 376024 405622 376076 405628
rect 383212 299470 383240 500140
rect 383856 497962 383884 500140
rect 383844 497956 383896 497962
rect 383844 497898 383896 497904
rect 383200 299464 383252 299470
rect 383200 299406 383252 299412
rect 384500 257378 384528 500140
rect 385144 499769 385172 500140
rect 385788 499905 385816 500140
rect 385774 499896 385830 499905
rect 385774 499831 385830 499840
rect 385130 499760 385186 499769
rect 385130 499695 385186 499704
rect 385144 497729 385172 499695
rect 385788 497865 385816 499831
rect 386432 498137 386460 500140
rect 386418 498128 386474 498137
rect 386418 498063 386474 498072
rect 387076 498001 387104 500140
rect 387720 499905 387748 500140
rect 387706 499896 387762 499905
rect 387706 499831 387762 499840
rect 387062 497992 387118 498001
rect 388364 497962 388392 500140
rect 389652 499050 389680 500140
rect 390296 499905 390324 500140
rect 390282 499896 390338 499905
rect 390282 499831 390338 499840
rect 389640 499044 389692 499050
rect 389640 498986 389692 498992
rect 387062 497927 387118 497936
rect 388352 497956 388404 497962
rect 388352 497898 388404 497904
rect 385774 497856 385830 497865
rect 385774 497791 385830 497800
rect 385130 497720 385186 497729
rect 385130 497655 385186 497664
rect 389180 479528 389232 479534
rect 389180 479470 389232 479476
rect 385040 352572 385092 352578
rect 385040 352514 385092 352520
rect 384488 257372 384540 257378
rect 384488 257314 384540 257320
rect 382280 177336 382332 177342
rect 382280 177278 382332 177284
rect 378140 17264 378192 17270
rect 378140 17206 378192 17212
rect 378152 16574 378180 17206
rect 382292 16574 382320 177278
rect 385052 16574 385080 352514
rect 389192 16574 389220 479470
rect 378152 16546 378456 16574
rect 382292 16546 382412 16574
rect 385052 16546 386000 16574
rect 389192 16546 389496 16574
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 371670 354 371782 480
rect 371252 326 371782 354
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378428 354 378456 16546
rect 382384 480 382412 16546
rect 385972 480 386000 16546
rect 389468 480 389496 16546
rect 390940 15978 390968 500140
rect 391584 497593 391612 500140
rect 391570 497584 391626 497593
rect 391570 497519 391626 497528
rect 391940 24132 391992 24138
rect 391940 24074 391992 24080
rect 391952 16574 391980 24074
rect 392228 21486 392256 500140
rect 392872 499905 392900 500140
rect 392858 499896 392914 499905
rect 392858 499831 392914 499840
rect 393516 497826 393544 500140
rect 394160 499526 394188 500140
rect 394148 499520 394200 499526
rect 394148 499462 394200 499468
rect 393504 497820 393556 497826
rect 393504 497762 393556 497768
rect 394804 497418 394832 500140
rect 395448 499905 395476 500140
rect 395434 499896 395490 499905
rect 395434 499831 395490 499840
rect 396092 499574 396120 500140
rect 396092 499546 396212 499574
rect 394792 497412 394844 497418
rect 394792 497354 394844 497360
rect 396080 493332 396132 493338
rect 396080 493274 396132 493280
rect 392216 21480 392268 21486
rect 392216 21422 392268 21428
rect 391952 16546 392624 16574
rect 390928 15972 390980 15978
rect 390928 15914 390980 15920
rect 378846 354 378958 480
rect 378428 326 378958 354
rect 378846 -960 378958 326
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 493274
rect 396184 8294 396212 499546
rect 396736 498098 396764 500140
rect 397380 499322 397408 500140
rect 397368 499316 397420 499322
rect 397368 499258 397420 499264
rect 398024 499118 398052 500140
rect 398012 499112 398064 499118
rect 398012 499054 398064 499060
rect 396724 498092 396776 498098
rect 396724 498034 396776 498040
rect 398668 498001 398696 500140
rect 399312 498166 399340 500140
rect 399496 499254 399524 501599
rect 399588 500954 399616 536279
rect 399956 533225 399984 639202
rect 400036 552968 400088 552974
rect 400036 552910 400088 552916
rect 400048 541566 400076 552910
rect 400126 541580 400182 541589
rect 400048 541538 400126 541566
rect 400126 541515 400182 541524
rect 399942 533216 399998 533225
rect 399942 533151 399998 533160
rect 400232 511669 400260 640426
rect 400324 517789 400352 640630
rect 400416 552838 400444 642058
rect 400588 641912 400640 641918
rect 400588 641854 400640 641860
rect 400496 639192 400548 639198
rect 400496 639134 400548 639140
rect 400404 552832 400456 552838
rect 400404 552774 400456 552780
rect 400508 552566 400536 639134
rect 400600 599826 400628 641854
rect 400588 599820 400640 599826
rect 400588 599762 400640 599768
rect 400692 599622 400720 642126
rect 400784 599758 400812 642534
rect 400864 642320 400916 642326
rect 400864 642262 400916 642268
rect 400772 599752 400824 599758
rect 400772 599694 400824 599700
rect 400680 599616 400732 599622
rect 400680 599558 400732 599564
rect 400588 597848 400640 597854
rect 400588 597790 400640 597796
rect 400496 552560 400548 552566
rect 400496 552502 400548 552508
rect 400496 550520 400548 550526
rect 400496 550462 400548 550468
rect 400402 526620 400458 526629
rect 400402 526555 400458 526564
rect 400416 525842 400444 526555
rect 400404 525836 400456 525842
rect 400404 525778 400456 525784
rect 400310 517780 400366 517789
rect 400310 517715 400366 517724
rect 400508 514865 400536 550462
rect 400600 549778 400628 597790
rect 400772 551676 400824 551682
rect 400772 551618 400824 551624
rect 400680 549908 400732 549914
rect 400680 549850 400732 549856
rect 400588 549772 400640 549778
rect 400588 549714 400640 549720
rect 400600 549574 400628 549714
rect 400588 549568 400640 549574
rect 400588 549510 400640 549516
rect 400692 526697 400720 549850
rect 400784 532545 400812 551618
rect 400876 534138 400904 642262
rect 402336 640552 402388 640558
rect 402336 640494 402388 640500
rect 402152 639056 402204 639062
rect 402152 638998 402204 639004
rect 401784 638988 401836 638994
rect 401784 638930 401836 638936
rect 400956 559564 401008 559570
rect 400956 559506 401008 559512
rect 400968 539345 400996 559506
rect 401232 554056 401284 554062
rect 401232 553998 401284 554004
rect 401138 551576 401194 551585
rect 401138 551511 401194 551520
rect 401048 549772 401100 549778
rect 401048 549714 401100 549720
rect 400954 539336 401010 539345
rect 400954 539271 401010 539280
rect 401060 538121 401088 549714
rect 401046 538112 401102 538121
rect 401046 538047 401102 538056
rect 400864 534132 400916 534138
rect 400864 534074 400916 534080
rect 400770 532536 400826 532545
rect 400770 532471 400826 532480
rect 400678 526688 400734 526697
rect 400678 526623 400734 526632
rect 401152 523025 401180 551511
rect 401138 523016 401194 523025
rect 401138 522951 401194 522960
rect 400494 514856 400550 514865
rect 400494 514791 400550 514800
rect 400864 514820 400916 514826
rect 400864 514762 400916 514768
rect 400218 511660 400274 511669
rect 400218 511595 400274 511604
rect 399576 500948 399628 500954
rect 399576 500890 399628 500896
rect 399484 499248 399536 499254
rect 399484 499190 399536 499196
rect 399300 498160 399352 498166
rect 399300 498102 399352 498108
rect 398654 497992 398710 498001
rect 398654 497927 398710 497936
rect 398840 497548 398892 497554
rect 398840 497490 398892 497496
rect 396172 8288 396224 8294
rect 396172 8230 396224 8236
rect 398852 3398 398880 497490
rect 400876 15910 400904 514762
rect 401244 505073 401272 553998
rect 401600 552016 401652 552022
rect 401600 551958 401652 551964
rect 401612 535401 401640 551958
rect 401692 550588 401744 550594
rect 401692 550530 401744 550536
rect 401598 535392 401654 535401
rect 401598 535327 401654 535336
rect 401600 533928 401652 533934
rect 401600 533870 401652 533876
rect 401612 533633 401640 533870
rect 401598 533624 401654 533633
rect 401598 533559 401654 533568
rect 401600 530256 401652 530262
rect 401600 530198 401652 530204
rect 401612 530097 401640 530198
rect 401598 530088 401654 530097
rect 401598 530023 401654 530032
rect 401600 529168 401652 529174
rect 401600 529110 401652 529116
rect 401612 528873 401640 529110
rect 401598 528864 401654 528873
rect 401598 528799 401654 528808
rect 401600 528488 401652 528494
rect 401600 528430 401652 528436
rect 401612 528193 401640 528430
rect 401598 528184 401654 528193
rect 401598 528119 401654 528128
rect 401600 526448 401652 526454
rect 401600 526390 401652 526396
rect 401612 526153 401640 526390
rect 401598 526144 401654 526153
rect 401598 526079 401654 526088
rect 401600 525768 401652 525774
rect 401600 525710 401652 525716
rect 401612 525473 401640 525710
rect 401598 525464 401654 525473
rect 401598 525399 401654 525408
rect 401600 525292 401652 525298
rect 401600 525234 401652 525240
rect 401612 524929 401640 525234
rect 401598 524920 401654 524929
rect 401598 524855 401654 524864
rect 401600 524408 401652 524414
rect 401600 524350 401652 524356
rect 401612 524113 401640 524350
rect 401598 524104 401654 524113
rect 401598 524039 401654 524048
rect 401598 521792 401654 521801
rect 401598 521727 401654 521736
rect 401612 521694 401640 521727
rect 401600 521688 401652 521694
rect 401600 521630 401652 521636
rect 401600 521076 401652 521082
rect 401600 521018 401652 521024
rect 401612 520849 401640 521018
rect 401598 520840 401654 520849
rect 401598 520775 401654 520784
rect 401600 520192 401652 520198
rect 401600 520134 401652 520140
rect 401612 520033 401640 520134
rect 401598 520024 401654 520033
rect 401598 519959 401654 519968
rect 401704 517449 401732 550530
rect 401796 543590 401824 638930
rect 401968 562420 402020 562426
rect 401968 562362 402020 562368
rect 401876 554124 401928 554130
rect 401876 554066 401928 554072
rect 401784 543584 401836 543590
rect 401784 543526 401836 543532
rect 401784 543448 401836 543454
rect 401784 543390 401836 543396
rect 401796 543153 401824 543390
rect 401782 543144 401838 543153
rect 401782 543079 401838 543088
rect 401782 541784 401838 541793
rect 401782 541719 401838 541728
rect 401796 541006 401824 541719
rect 401784 541000 401836 541006
rect 401784 540942 401836 540948
rect 401782 530360 401838 530369
rect 401782 530295 401838 530304
rect 401796 529990 401824 530295
rect 401784 529984 401836 529990
rect 401784 529926 401836 529932
rect 401782 529000 401838 529009
rect 401782 528935 401838 528944
rect 401796 528698 401824 528935
rect 401784 528692 401836 528698
rect 401784 528634 401836 528640
rect 401782 528592 401838 528601
rect 401782 528527 401838 528536
rect 401690 517440 401746 517449
rect 401690 517375 401746 517384
rect 401598 516352 401654 516361
rect 401598 516287 401654 516296
rect 401612 516186 401640 516287
rect 401600 516180 401652 516186
rect 401600 516122 401652 516128
rect 401692 516112 401744 516118
rect 401692 516054 401744 516060
rect 401704 515953 401732 516054
rect 401690 515944 401746 515953
rect 401690 515879 401746 515888
rect 401690 513904 401746 513913
rect 401690 513839 401746 513848
rect 401600 506456 401652 506462
rect 401598 506424 401600 506433
rect 401652 506424 401654 506433
rect 401598 506359 401654 506368
rect 401230 505064 401286 505073
rect 401230 504999 401286 505008
rect 401600 503668 401652 503674
rect 401600 503610 401652 503616
rect 401612 503305 401640 503610
rect 401598 503296 401654 503305
rect 401598 503231 401654 503240
rect 401598 500304 401654 500313
rect 401598 500239 401654 500248
rect 401612 499594 401640 500239
rect 401600 499588 401652 499594
rect 401600 499530 401652 499536
rect 401704 497622 401732 513839
rect 401796 504665 401824 528527
rect 401888 508337 401916 554066
rect 401980 521665 402008 562362
rect 402060 560992 402112 560998
rect 402060 560934 402112 560940
rect 402072 544785 402100 560934
rect 402058 544776 402114 544785
rect 402058 544711 402114 544720
rect 402060 543584 402112 543590
rect 402060 543526 402112 543532
rect 402072 540977 402100 543526
rect 402058 540968 402114 540977
rect 402058 540903 402114 540912
rect 402060 534132 402112 534138
rect 402060 534074 402112 534080
rect 402072 528601 402100 534074
rect 402058 528592 402114 528601
rect 402058 528527 402114 528536
rect 401966 521656 402022 521665
rect 401966 521591 402022 521600
rect 401966 513496 402022 513505
rect 401966 513431 402022 513440
rect 401874 508328 401930 508337
rect 401874 508263 401930 508272
rect 401782 504656 401838 504665
rect 401782 504591 401838 504600
rect 401980 500886 402008 513431
rect 402164 510513 402192 638998
rect 402242 558240 402298 558249
rect 402242 558175 402298 558184
rect 402256 547777 402284 558175
rect 402242 547768 402298 547777
rect 402242 547703 402298 547712
rect 402348 540705 402376 640494
rect 403164 639328 403216 639334
rect 403164 639270 403216 639276
rect 402980 554872 403032 554878
rect 402980 554814 403032 554820
rect 402428 552696 402480 552702
rect 402428 552638 402480 552644
rect 402440 547505 402468 552638
rect 402426 547496 402482 547505
rect 402426 547431 402482 547440
rect 402520 546508 402572 546514
rect 402520 546450 402572 546456
rect 402334 540696 402390 540705
rect 402334 540631 402390 540640
rect 402532 534721 402560 546450
rect 402886 546408 402942 546417
rect 402992 546394 403020 554814
rect 403072 551540 403124 551546
rect 403072 551482 403124 551488
rect 402942 546366 403020 546394
rect 402886 546343 402942 546352
rect 402886 546136 402942 546145
rect 403084 546122 403112 551482
rect 402942 546094 403112 546122
rect 402886 546071 402942 546080
rect 402980 540048 403032 540054
rect 402980 539990 403032 539996
rect 402518 534712 402574 534721
rect 402518 534647 402574 534656
rect 402334 514856 402390 514865
rect 402334 514791 402390 514800
rect 402150 510504 402206 510513
rect 402150 510439 402206 510448
rect 402058 508464 402114 508473
rect 402058 508399 402114 508408
rect 401968 500880 402020 500886
rect 401968 500822 402020 500828
rect 401692 497616 401744 497622
rect 401692 497558 401744 497564
rect 402072 497486 402100 508399
rect 402348 499186 402376 514791
rect 402428 513120 402480 513126
rect 402428 513062 402480 513068
rect 402440 512825 402468 513062
rect 402426 512816 402482 512825
rect 402426 512751 402482 512760
rect 402886 510776 402942 510785
rect 402886 510711 402942 510720
rect 402900 510678 402928 510711
rect 402888 510672 402940 510678
rect 402888 510614 402940 510620
rect 402886 509416 402942 509425
rect 402886 509351 402942 509360
rect 402900 509318 402928 509351
rect 402888 509312 402940 509318
rect 402888 509254 402940 509260
rect 402336 499180 402388 499186
rect 402336 499122 402388 499128
rect 402060 497480 402112 497486
rect 402060 497422 402112 497428
rect 400864 15904 400916 15910
rect 400864 15846 400916 15852
rect 402520 8288 402572 8294
rect 402520 8230 402572 8236
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 402532 480 402560 8230
rect 402992 6914 403020 539990
rect 403176 498098 403204 639270
rect 403268 526454 403296 662458
rect 403624 634840 403676 634846
rect 403624 634782 403676 634788
rect 403636 600302 403664 634782
rect 403624 600296 403676 600302
rect 403624 600238 403676 600244
rect 403440 552356 403492 552362
rect 403440 552298 403492 552304
rect 403348 551472 403400 551478
rect 403348 551414 403400 551420
rect 403256 526448 403308 526454
rect 403256 526390 403308 526396
rect 403360 506462 403388 551414
rect 403452 521082 403480 552298
rect 403532 551404 403584 551410
rect 403532 551346 403584 551352
rect 403544 530262 403572 551346
rect 403624 541340 403676 541346
rect 403624 541282 403676 541288
rect 403532 530256 403584 530262
rect 403532 530198 403584 530204
rect 403440 521076 403492 521082
rect 403440 521018 403492 521024
rect 403348 506456 403400 506462
rect 403348 506398 403400 506404
rect 403164 498092 403216 498098
rect 403164 498034 403216 498040
rect 403636 16574 403664 541282
rect 403728 499526 403756 670686
rect 403808 642660 403860 642666
rect 403808 642602 403860 642608
rect 403820 529174 403848 642602
rect 404636 639532 404688 639538
rect 404636 639474 404688 639480
rect 403900 639124 403952 639130
rect 403900 639066 403952 639072
rect 403808 529168 403860 529174
rect 403808 529110 403860 529116
rect 403716 499520 403768 499526
rect 403716 499462 403768 499468
rect 403912 498166 403940 639066
rect 404544 554804 404596 554810
rect 404544 554746 404596 554752
rect 404452 551336 404504 551342
rect 404452 551278 404504 551284
rect 404360 550724 404412 550730
rect 404360 550666 404412 550672
rect 404372 525298 404400 550666
rect 404464 528494 404492 551278
rect 404556 543454 404584 554746
rect 404544 543448 404596 543454
rect 404544 543390 404596 543396
rect 404452 528488 404504 528494
rect 404452 528430 404504 528436
rect 404648 525774 404676 639474
rect 404728 598324 404780 598330
rect 404728 598266 404780 598272
rect 404636 525768 404688 525774
rect 404636 525710 404688 525716
rect 404360 525292 404412 525298
rect 404360 525234 404412 525240
rect 404740 516118 404768 598266
rect 404820 598256 404872 598262
rect 404820 598198 404872 598204
rect 404832 524414 404860 598198
rect 404912 565888 404964 565894
rect 404912 565830 404964 565836
rect 404924 533934 404952 565830
rect 405016 559745 405044 700470
rect 406476 700392 406528 700398
rect 406476 700334 406528 700340
rect 405280 662448 405332 662454
rect 405280 662390 405332 662396
rect 405188 642252 405240 642258
rect 405188 642194 405240 642200
rect 405002 559736 405058 559745
rect 405002 559671 405058 559680
rect 405004 539640 405056 539646
rect 405004 539582 405056 539588
rect 404912 533928 404964 533934
rect 404912 533870 404964 533876
rect 404820 524408 404872 524414
rect 404820 524350 404872 524356
rect 404728 516112 404780 516118
rect 404728 516054 404780 516060
rect 403900 498160 403952 498166
rect 403900 498102 403952 498108
rect 403636 16546 403756 16574
rect 402992 6886 403664 6914
rect 403636 480 403664 6886
rect 403728 3670 403756 16546
rect 405016 3874 405044 539582
rect 405096 528692 405148 528698
rect 405096 528634 405148 528640
rect 405108 167006 405136 528634
rect 405200 497962 405228 642194
rect 405292 520198 405320 662390
rect 405372 642456 405424 642462
rect 405372 642398 405424 642404
rect 405280 520192 405332 520198
rect 405280 520134 405332 520140
rect 405384 513126 405412 642398
rect 406384 641776 406436 641782
rect 406384 641718 406436 641724
rect 406396 599146 406424 641718
rect 406384 599140 406436 599146
rect 406384 599082 406436 599088
rect 406384 541408 406436 541414
rect 406384 541350 406436 541356
rect 405740 516180 405792 516186
rect 405740 516122 405792 516128
rect 405372 513120 405424 513126
rect 405372 513062 405424 513068
rect 405188 497956 405240 497962
rect 405188 497898 405240 497904
rect 405096 167000 405148 167006
rect 405096 166942 405148 166948
rect 405752 16574 405780 516122
rect 405752 16546 406056 16574
rect 405004 3868 405056 3874
rect 405004 3810 405056 3816
rect 403716 3664 403768 3670
rect 403716 3606 403768 3612
rect 406028 480 406056 16546
rect 406396 3806 406424 541350
rect 406488 499322 406516 700334
rect 407120 661292 407172 661298
rect 407120 661234 407172 661240
rect 407132 503674 407160 661234
rect 409144 552288 409196 552294
rect 409144 552230 409196 552236
rect 407120 503668 407172 503674
rect 407120 503610 407172 503616
rect 406476 499316 406528 499322
rect 406476 499258 406528 499264
rect 408500 496188 408552 496194
rect 408500 496130 408552 496136
rect 407120 490612 407172 490618
rect 407120 490554 407172 490560
rect 407132 16574 407160 490554
rect 408512 16574 408540 496130
rect 409156 206990 409184 552230
rect 409248 499254 409276 700538
rect 410524 539776 410576 539782
rect 410524 539718 410576 539724
rect 409236 499248 409288 499254
rect 409236 499190 409288 499196
rect 409880 497480 409932 497486
rect 409880 497422 409932 497428
rect 409144 206984 409196 206990
rect 409144 206926 409196 206932
rect 409892 16574 409920 497422
rect 407132 16546 407252 16574
rect 408512 16546 409184 16574
rect 409892 16546 410472 16574
rect 406384 3800 406436 3806
rect 406384 3742 406436 3748
rect 407224 480 407252 16546
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410444 3482 410472 16546
rect 410536 3602 410564 539718
rect 412652 527134 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 458824 698964 458876 698970
rect 458824 698906 458876 698912
rect 427084 694816 427136 694822
rect 427084 694758 427136 694764
rect 419540 550792 419592 550798
rect 419540 550734 419592 550740
rect 416780 543040 416832 543046
rect 416780 542982 416832 542988
rect 412640 527128 412692 527134
rect 412640 527070 412692 527076
rect 414020 518968 414072 518974
rect 414020 518910 414072 518916
rect 413284 513392 413336 513398
rect 413284 513334 413336 513340
rect 413296 22778 413324 513334
rect 413284 22772 413336 22778
rect 413284 22714 413336 22720
rect 412640 21480 412692 21486
rect 412640 21422 412692 21428
rect 410524 3596 410576 3602
rect 410524 3538 410576 3544
rect 410444 3454 410840 3482
rect 410812 480 410840 3454
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 412652 354 412680 21422
rect 414032 16574 414060 518910
rect 415400 89004 415452 89010
rect 415400 88946 415452 88952
rect 414032 16546 414336 16574
rect 414308 480 414336 16546
rect 415412 3602 415440 88946
rect 416792 16574 416820 542982
rect 418804 527196 418856 527202
rect 418804 527138 418856 527144
rect 416792 16546 417464 16574
rect 415400 3596 415452 3602
rect 415400 3538 415452 3544
rect 416688 3596 416740 3602
rect 416688 3538 416740 3544
rect 416700 480 416728 3538
rect 413070 354 413182 480
rect 412652 326 413182 354
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 418816 14550 418844 527138
rect 418896 66292 418948 66298
rect 418896 66234 418948 66240
rect 418804 14544 418856 14550
rect 418804 14486 418856 14492
rect 418908 7682 418936 66234
rect 419552 16574 419580 550734
rect 420920 543108 420972 543114
rect 420920 543050 420972 543056
rect 419552 16546 420224 16574
rect 418896 7676 418948 7682
rect 418896 7618 418948 7624
rect 420196 480 420224 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 543050
rect 423680 542564 423732 542570
rect 423680 542506 423732 542512
rect 423036 533384 423088 533390
rect 423036 533326 423088 533332
rect 422944 524476 422996 524482
rect 422944 524418 422996 524424
rect 422956 21418 422984 524418
rect 423048 241466 423076 533326
rect 423036 241460 423088 241466
rect 423036 241402 423088 241408
rect 422944 21412 422996 21418
rect 422944 21354 422996 21360
rect 423692 3602 423720 542506
rect 423772 521688 423824 521694
rect 423772 521630 423824 521636
rect 423680 3596 423732 3602
rect 423680 3538 423732 3544
rect 423784 480 423812 521630
rect 427096 517478 427124 694758
rect 430580 552220 430632 552226
rect 430580 552162 430632 552168
rect 427820 543176 427872 543182
rect 427820 543118 427872 543124
rect 427084 517472 427136 517478
rect 427084 517414 427136 517420
rect 427728 509924 427780 509930
rect 427728 509866 427780 509872
rect 427740 509318 427768 509866
rect 427728 509312 427780 509318
rect 427728 509254 427780 509260
rect 426440 175976 426492 175982
rect 426440 175918 426492 175924
rect 426452 16574 426480 175918
rect 426452 16546 426848 16574
rect 424968 3596 425020 3602
rect 424968 3538 425020 3544
rect 424980 480 425008 3538
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 426820 354 426848 16546
rect 427740 9110 427768 509254
rect 427832 16574 427860 543118
rect 430592 16574 430620 552162
rect 448520 550656 448572 550662
rect 448520 550598 448572 550604
rect 438860 542700 438912 542706
rect 438860 542642 438912 542648
rect 436836 541136 436888 541142
rect 436836 541078 436888 541084
rect 432604 525836 432656 525842
rect 432604 525778 432656 525784
rect 432616 511970 432644 525778
rect 436744 512032 436796 512038
rect 436744 511974 436796 511980
rect 432604 511964 432656 511970
rect 432604 511906 432656 511912
rect 431960 506524 432012 506530
rect 431960 506466 432012 506472
rect 431972 16574 432000 506466
rect 434720 501016 434772 501022
rect 434720 500958 434772 500964
rect 433340 499588 433392 499594
rect 433340 499530 433392 499536
rect 433352 16574 433380 499530
rect 434732 16574 434760 500958
rect 436756 32434 436784 511974
rect 436848 255270 436876 541078
rect 437480 541000 437532 541006
rect 437480 540942 437532 540948
rect 436836 255264 436888 255270
rect 436836 255206 436888 255212
rect 436744 32428 436796 32434
rect 436744 32370 436796 32376
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 431972 16546 432092 16574
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 427728 9104 427780 9110
rect 427728 9046 427780 9052
rect 428476 480 428504 16546
rect 430868 480 430896 16546
rect 432064 480 432092 16546
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 540942
rect 438872 16574 438900 542642
rect 440884 541204 440936 541210
rect 440884 541146 440936 541152
rect 440896 109002 440924 541146
rect 445760 507884 445812 507890
rect 445760 507826 445812 507832
rect 441620 493400 441672 493406
rect 441620 493342 441672 493348
rect 440884 108996 440936 109002
rect 440884 108938 440936 108944
rect 441632 16574 441660 493342
rect 444378 44840 444434 44849
rect 444378 44775 444434 44784
rect 444392 16574 444420 44775
rect 438872 16546 439176 16574
rect 441632 16546 442672 16574
rect 444392 16546 445064 16574
rect 439148 480 439176 16546
rect 440240 15972 440292 15978
rect 440240 15914 440292 15920
rect 440252 3602 440280 15914
rect 440240 3596 440292 3602
rect 440240 3538 440292 3544
rect 441528 3596 441580 3602
rect 441528 3538 441580 3544
rect 441540 480 441568 3538
rect 442644 480 442672 16546
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 507826
rect 448532 16574 448560 550598
rect 454776 532772 454828 532778
rect 454776 532714 454828 532720
rect 452660 528624 452712 528630
rect 452660 528566 452712 528572
rect 450544 517540 450596 517546
rect 450544 517482 450596 517488
rect 450556 20670 450584 517482
rect 451280 510672 451332 510678
rect 451280 510614 451332 510620
rect 450544 20664 450596 20670
rect 450544 20606 450596 20612
rect 451292 16574 451320 510614
rect 452672 16574 452700 528566
rect 454684 499588 454736 499594
rect 454684 499530 454736 499536
rect 454696 28286 454724 499530
rect 454788 224262 454816 532714
rect 458836 531282 458864 698906
rect 458824 531276 458876 531282
rect 458824 531218 458876 531224
rect 458180 529984 458232 529990
rect 458180 529926 458232 529932
rect 457444 514888 457496 514894
rect 457444 514830 457496 514836
rect 456800 497616 456852 497622
rect 456800 497558 456852 497564
rect 455420 493468 455472 493474
rect 455420 493410 455472 493416
rect 454776 224256 454828 224262
rect 454776 224198 454828 224204
rect 454684 28280 454736 28286
rect 454684 28222 454736 28228
rect 455432 16574 455460 493410
rect 456812 16574 456840 497558
rect 457456 267034 457484 514830
rect 457444 267028 457496 267034
rect 457444 266970 457496 266976
rect 458192 16574 458220 529926
rect 460204 525836 460256 525842
rect 460204 525778 460256 525784
rect 459560 497684 459612 497690
rect 459560 497626 459612 497632
rect 459572 16574 459600 497626
rect 460216 480962 460244 525778
rect 462332 500274 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 472716 700324 472768 700330
rect 472716 700266 472768 700272
rect 468668 596828 468720 596834
rect 468668 596770 468720 596776
rect 466460 542428 466512 542434
rect 466460 542370 466512 542376
rect 463700 531344 463752 531350
rect 463700 531286 463752 531292
rect 462964 502376 463016 502382
rect 462964 502318 463016 502324
rect 462320 500268 462372 500274
rect 462320 500210 462372 500216
rect 460204 480956 460256 480962
rect 460204 480898 460256 480904
rect 462976 17270 463004 502318
rect 462964 17264 463016 17270
rect 462964 17206 463016 17212
rect 463712 16574 463740 531286
rect 466472 16574 466500 542370
rect 468484 517608 468536 517614
rect 468484 517550 468536 517556
rect 468496 24138 468524 517550
rect 468680 509930 468708 596770
rect 470600 542972 470652 542978
rect 470600 542914 470652 542920
rect 468668 509924 468720 509930
rect 468668 509866 468720 509872
rect 468576 509312 468628 509318
rect 468576 509254 468628 509260
rect 468588 280158 468616 509254
rect 468576 280152 468628 280158
rect 468576 280094 468628 280100
rect 468484 24132 468536 24138
rect 468484 24074 468536 24080
rect 448532 16546 448652 16574
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 455432 16546 455736 16574
rect 456812 16546 456932 16574
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 448624 480 448652 16546
rect 449808 3596 449860 3602
rect 449808 3538 449860 3544
rect 449820 480 449848 3538
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 455708 480 455736 16546
rect 456904 480 456932 16546
rect 459204 480 459232 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 463988 480 464016 16546
rect 467484 480 467512 16546
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 542914
rect 472624 542768 472676 542774
rect 472624 542710 472676 542716
rect 472636 26926 472664 542710
rect 472728 499526 472756 700266
rect 476948 665848 477000 665854
rect 476948 665790 477000 665796
rect 475384 641844 475436 641850
rect 475384 641786 475436 641792
rect 475396 599078 475424 641786
rect 475384 599072 475436 599078
rect 475384 599014 475436 599020
rect 472808 598256 472860 598262
rect 472808 598198 472860 598204
rect 472716 499520 472768 499526
rect 472716 499462 472768 499468
rect 472820 499390 472848 598198
rect 475568 580304 475620 580310
rect 475568 580246 475620 580252
rect 473360 542836 473412 542842
rect 473360 542778 473412 542784
rect 472808 499384 472860 499390
rect 472808 499326 472860 499332
rect 472624 26920 472676 26926
rect 472624 26862 472676 26868
rect 473372 3398 473400 542778
rect 475476 542632 475528 542638
rect 475476 542574 475528 542580
rect 475384 541272 475436 541278
rect 475384 541214 475436 541220
rect 473452 177404 473504 177410
rect 473452 177346 473504 177352
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 473464 480 473492 177346
rect 475396 3738 475424 541214
rect 475488 25566 475516 542574
rect 475580 498098 475608 580246
rect 476764 542904 476816 542910
rect 476764 542846 476816 542852
rect 475568 498092 475620 498098
rect 475568 498034 475620 498040
rect 475476 25560 475528 25566
rect 475476 25502 475528 25508
rect 476776 18630 476804 542846
rect 476856 512100 476908 512106
rect 476856 512042 476908 512048
rect 476868 28354 476896 512042
rect 476960 510542 476988 665790
rect 477512 654134 477540 702406
rect 527192 699718 527220 703520
rect 543476 700466 543504 703520
rect 559668 700534 559696 703520
rect 559656 700528 559708 700534
rect 559656 700470 559708 700476
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 526444 699712 526496 699718
rect 526444 699654 526496 699660
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 525064 696992 525116 696998
rect 525064 696934 525116 696940
rect 479524 667208 479576 667214
rect 479524 667150 479576 667156
rect 478328 661224 478380 661230
rect 478328 661166 478380 661172
rect 477512 654106 477632 654134
rect 477040 643748 477092 643754
rect 477040 643690 477092 643696
rect 476948 510536 477000 510542
rect 476948 510478 477000 510484
rect 477052 498030 477080 643690
rect 477604 625154 477632 654106
rect 477682 636168 477738 636177
rect 477682 636103 477738 636112
rect 477696 634846 477724 636103
rect 477684 634840 477736 634846
rect 477684 634782 477736 634788
rect 477512 625126 477632 625154
rect 477512 506818 477540 625126
rect 478142 617808 478198 617817
rect 478142 617743 478198 617752
rect 478156 598806 478184 617743
rect 478144 598800 478196 598806
rect 478144 598742 478196 598748
rect 478236 542496 478288 542502
rect 478236 542438 478288 542444
rect 477590 534304 477646 534313
rect 477590 534239 477646 534248
rect 477604 533390 477632 534239
rect 477592 533384 477644 533390
rect 477592 533326 477644 533332
rect 477590 532808 477646 532817
rect 477590 532743 477592 532752
rect 477644 532743 477646 532752
rect 477592 532714 477644 532720
rect 477590 531448 477646 531457
rect 477590 531383 477646 531392
rect 477604 531350 477632 531383
rect 477592 531344 477644 531350
rect 477592 531286 477644 531292
rect 477590 529000 477646 529009
rect 477590 528935 477646 528944
rect 477604 528630 477632 528935
rect 477592 528624 477644 528630
rect 477592 528566 477644 528572
rect 477590 527232 477646 527241
rect 477590 527167 477592 527176
rect 477644 527167 477646 527176
rect 477592 527138 477644 527144
rect 477684 527128 477736 527134
rect 477684 527070 477736 527076
rect 477696 526833 477724 527070
rect 477682 526824 477738 526833
rect 477682 526759 477738 526768
rect 477590 525872 477646 525881
rect 477590 525807 477592 525816
rect 477644 525807 477646 525816
rect 477592 525778 477644 525784
rect 478142 524920 478198 524929
rect 478142 524855 478198 524864
rect 478156 524482 478184 524855
rect 478144 524476 478196 524482
rect 478144 524418 478196 524424
rect 477866 520296 477922 520305
rect 477866 520231 477922 520240
rect 477590 519344 477646 519353
rect 477590 519279 477646 519288
rect 477604 518974 477632 519279
rect 477592 518968 477644 518974
rect 477592 518910 477644 518916
rect 477590 517984 477646 517993
rect 477590 517919 477646 517928
rect 477604 517614 477632 517919
rect 477682 517712 477738 517721
rect 477682 517647 477738 517656
rect 477592 517608 477644 517614
rect 477592 517550 477644 517556
rect 477696 517546 477724 517647
rect 477684 517540 477736 517546
rect 477684 517482 477736 517488
rect 477592 517472 477644 517478
rect 477592 517414 477644 517420
rect 477604 517313 477632 517414
rect 477590 517304 477646 517313
rect 477590 517239 477646 517248
rect 477682 515264 477738 515273
rect 477682 515199 477738 515208
rect 477590 514992 477646 515001
rect 477590 514927 477646 514936
rect 477604 514894 477632 514927
rect 477592 514888 477644 514894
rect 477592 514830 477644 514836
rect 477696 514826 477724 515199
rect 477684 514820 477736 514826
rect 477684 514762 477736 514768
rect 477590 513904 477646 513913
rect 477590 513839 477646 513848
rect 477604 513398 477632 513839
rect 477592 513392 477644 513398
rect 477592 513334 477644 513340
rect 477682 512544 477738 512553
rect 477682 512479 477738 512488
rect 477696 512038 477724 512479
rect 477684 512032 477736 512038
rect 477684 511974 477736 511980
rect 477592 511964 477644 511970
rect 477592 511906 477644 511912
rect 477604 511873 477632 511906
rect 477590 511864 477646 511873
rect 477590 511799 477646 511808
rect 477590 509416 477646 509425
rect 477590 509351 477646 509360
rect 477604 509318 477632 509351
rect 477592 509312 477644 509318
rect 477592 509254 477644 509260
rect 477512 506790 477724 506818
rect 477498 506696 477554 506705
rect 477498 506631 477554 506640
rect 477512 506530 477540 506631
rect 477500 506524 477552 506530
rect 477500 506466 477552 506472
rect 477498 502888 477554 502897
rect 477498 502823 477554 502832
rect 477512 502382 477540 502823
rect 477500 502376 477552 502382
rect 477500 502318 477552 502324
rect 477590 501664 477646 501673
rect 477590 501599 477646 501608
rect 477498 501256 477554 501265
rect 477498 501191 477554 501200
rect 477512 501022 477540 501191
rect 477500 501016 477552 501022
rect 477500 500958 477552 500964
rect 477408 500268 477460 500274
rect 477408 500210 477460 500216
rect 477040 498024 477092 498030
rect 477040 497966 477092 497972
rect 477420 497962 477448 500210
rect 477498 500168 477554 500177
rect 477498 500103 477554 500112
rect 477512 499594 477540 500103
rect 477500 499588 477552 499594
rect 477500 499530 477552 499536
rect 477604 498817 477632 501599
rect 477696 499390 477724 506790
rect 477684 499384 477736 499390
rect 477684 499326 477736 499332
rect 477590 498808 477646 498817
rect 477590 498743 477646 498752
rect 477408 497956 477460 497962
rect 477408 497898 477460 497904
rect 477880 431934 477908 520231
rect 478142 512136 478198 512145
rect 478142 512071 478144 512080
rect 478196 512071 478198 512080
rect 478144 512042 478196 512048
rect 478144 510536 478196 510542
rect 478142 510504 478144 510513
rect 478196 510504 478198 510513
rect 478142 510439 478198 510448
rect 478142 508464 478198 508473
rect 478142 508399 478198 508408
rect 478156 507890 478184 508399
rect 478144 507884 478196 507890
rect 478144 507826 478196 507832
rect 478142 503840 478198 503849
rect 478142 503775 478198 503784
rect 477868 431928 477920 431934
rect 477868 431870 477920 431876
rect 478156 227050 478184 503775
rect 478248 268394 478276 542438
rect 478340 506433 478368 661166
rect 478420 661156 478472 661162
rect 478420 661098 478472 661104
rect 478432 535401 478460 661098
rect 478972 659932 479024 659938
rect 478972 659874 479024 659880
rect 478788 590708 478840 590714
rect 478788 590650 478840 590656
rect 478602 536208 478658 536217
rect 478602 536143 478658 536152
rect 478418 535392 478474 535401
rect 478418 535327 478474 535336
rect 478616 530482 478644 536143
rect 478800 534177 478828 590650
rect 478984 543590 479012 659874
rect 478972 543584 479024 543590
rect 478972 543526 479024 543532
rect 479062 537704 479118 537713
rect 479062 537639 479118 537648
rect 478786 534168 478842 534177
rect 478786 534103 478842 534112
rect 478696 531276 478748 531282
rect 478696 531218 478748 531224
rect 478708 530641 478736 531218
rect 478694 530632 478750 530641
rect 478694 530567 478750 530576
rect 478616 530454 478736 530482
rect 478602 528592 478658 528601
rect 478602 528527 478658 528536
rect 478418 523424 478474 523433
rect 478418 523359 478474 523368
rect 478326 506424 478382 506433
rect 478326 506359 478382 506368
rect 478432 499458 478460 523359
rect 478510 520704 478566 520713
rect 478510 520639 478566 520648
rect 478420 499452 478472 499458
rect 478420 499394 478472 499400
rect 478524 494766 478552 520639
rect 478512 494760 478564 494766
rect 478512 494702 478564 494708
rect 478616 492046 478644 528527
rect 478604 492040 478656 492046
rect 478604 491982 478656 491988
rect 478708 487898 478736 530454
rect 478970 523152 479026 523161
rect 478970 523087 479026 523096
rect 478786 521928 478842 521937
rect 478786 521863 478842 521872
rect 478800 500954 478828 521863
rect 478788 500948 478840 500954
rect 478788 500890 478840 500896
rect 478984 493542 479012 523087
rect 479076 496806 479104 537639
rect 479338 537024 479394 537033
rect 479338 536959 479394 536968
rect 479246 507104 479302 507113
rect 479246 507039 479302 507048
rect 479154 504384 479210 504393
rect 479154 504319 479210 504328
rect 479064 496800 479116 496806
rect 479064 496742 479116 496748
rect 478972 493536 479024 493542
rect 478972 493478 479024 493484
rect 478696 487892 478748 487898
rect 478696 487834 478748 487840
rect 479168 483682 479196 504319
rect 479260 492114 479288 507039
rect 479248 492108 479300 492114
rect 479248 492050 479300 492056
rect 479352 486470 479380 536959
rect 479536 498166 479564 667150
rect 521844 661768 521896 661774
rect 521844 661710 521896 661716
rect 520740 661700 520792 661706
rect 520740 661642 520792 661648
rect 502340 660476 502392 660482
rect 502340 660418 502392 660424
rect 502352 660249 502380 660418
rect 520464 660408 520516 660414
rect 520464 660350 520516 660356
rect 507860 660340 507912 660346
rect 507860 660282 507912 660288
rect 507872 660249 507900 660282
rect 502338 660240 502394 660249
rect 502338 660175 502394 660184
rect 507858 660240 507914 660249
rect 507858 660175 507914 660184
rect 520372 659864 520424 659870
rect 520372 659806 520424 659812
rect 493232 641844 493284 641850
rect 493232 641786 493284 641792
rect 493244 639962 493272 641786
rect 510620 641776 510672 641782
rect 510620 641718 510672 641724
rect 510632 639962 510660 641718
rect 493244 639934 493580 639962
rect 510632 639934 510968 639962
rect 479720 600086 480056 600114
rect 496464 600086 496800 600114
rect 513852 600086 514188 600114
rect 479720 596834 479748 600086
rect 496464 598262 496492 600086
rect 513852 598874 513880 600086
rect 513840 598868 513892 598874
rect 513840 598810 513892 598816
rect 496452 598256 496504 598262
rect 496452 598198 496504 598204
rect 502340 596896 502392 596902
rect 502340 596838 502392 596844
rect 479708 596828 479760 596834
rect 479708 596770 479760 596776
rect 480260 591320 480312 591326
rect 480260 591262 480312 591268
rect 479708 543584 479760 543590
rect 479708 543526 479760 543532
rect 479720 539866 479748 543526
rect 480272 539866 480300 591262
rect 502352 557534 502380 596838
rect 503720 595468 503772 595474
rect 503720 595410 503772 595416
rect 503732 557534 503760 595410
rect 502352 557506 502840 557534
rect 503732 557506 504128 557534
rect 498844 552152 498896 552158
rect 498844 552094 498896 552100
rect 482192 544400 482244 544406
rect 482192 544342 482244 544348
rect 482204 539866 482232 544342
rect 490746 543688 490802 543697
rect 490746 543623 490802 543632
rect 482284 543040 482336 543046
rect 482284 542982 482336 542988
rect 479720 539838 480056 539866
rect 480272 539838 480700 539866
rect 481988 539838 482232 539866
rect 482296 539866 482324 542982
rect 488172 542496 488224 542502
rect 488172 542438 488224 542444
rect 484860 542428 484912 542434
rect 484860 542370 484912 542376
rect 483020 541204 483072 541210
rect 483020 541146 483072 541152
rect 484768 541204 484820 541210
rect 484768 541146 484820 541152
rect 483032 539866 483060 541146
rect 484780 539866 484808 541146
rect 482296 539838 482632 539866
rect 483032 539838 483276 539866
rect 484564 539838 484808 539866
rect 484872 539866 484900 542370
rect 488080 541000 488132 541006
rect 488080 540942 488132 540948
rect 486976 539912 487028 539918
rect 484872 539838 485208 539866
rect 488092 539866 488120 540942
rect 487028 539860 487140 539866
rect 486976 539854 487140 539860
rect 486988 539838 487140 539854
rect 487784 539838 488120 539866
rect 488184 539866 488212 542438
rect 489828 539980 489880 539986
rect 489828 539922 489880 539928
rect 489840 539866 489868 539922
rect 490760 539866 490788 543623
rect 498856 543046 498884 552094
rect 498844 543040 498896 543046
rect 498844 542982 498896 542988
rect 499028 542972 499080 542978
rect 499028 542914 499080 542920
rect 494060 542700 494112 542706
rect 494060 542642 494112 542648
rect 493232 541408 493284 541414
rect 493232 541350 493284 541356
rect 492588 541068 492640 541074
rect 492588 541010 492640 541016
rect 492600 539866 492628 541010
rect 488184 539838 488428 539866
rect 489716 539838 489868 539866
rect 490360 539850 490696 539866
rect 490360 539844 490708 539850
rect 490360 539838 490656 539844
rect 490760 539838 491004 539866
rect 492292 539838 492628 539866
rect 493244 539866 493272 541350
rect 494072 539866 494100 542642
rect 495440 541340 495492 541346
rect 495440 541282 495492 541288
rect 495452 539866 495480 541282
rect 498382 541104 498438 541113
rect 498382 541039 498438 541048
rect 498396 539866 498424 541039
rect 499040 539866 499068 542914
rect 500316 542564 500368 542570
rect 500316 542506 500368 542512
rect 500328 539866 500356 542506
rect 500960 540048 501012 540054
rect 500960 539990 501012 539996
rect 500972 539866 501000 539990
rect 502812 539866 502840 557506
rect 503996 542564 504048 542570
rect 503996 542506 504048 542512
rect 504008 539866 504036 542506
rect 493244 539838 493580 539866
rect 494072 539838 494224 539866
rect 495452 539838 495512 539866
rect 498396 539838 498732 539866
rect 499040 539838 499376 539866
rect 500328 539838 500664 539866
rect 500972 539838 501308 539866
rect 502812 539838 503240 539866
rect 503884 539838 504036 539866
rect 504100 539866 504128 557506
rect 508318 543552 508374 543561
rect 508318 543487 508374 543496
rect 506112 542904 506164 542910
rect 506112 542846 506164 542852
rect 506124 539866 506152 542846
rect 506754 539880 506810 539889
rect 504100 539838 504528 539866
rect 506124 539838 506460 539866
rect 506810 539838 507104 539866
rect 506754 539815 506810 539824
rect 490656 539786 490708 539792
rect 496452 539776 496504 539782
rect 486146 539744 486202 539753
rect 485852 539702 486146 539730
rect 495806 539744 495862 539753
rect 492936 539714 493272 539730
rect 492936 539708 493284 539714
rect 492936 539702 493232 539708
rect 486146 539679 486202 539688
rect 495862 539702 496156 539730
rect 498200 539776 498252 539782
rect 496504 539724 496800 539730
rect 496452 539718 496800 539724
rect 496464 539702 496800 539718
rect 498088 539724 498200 539730
rect 502154 539744 502210 539753
rect 498088 539718 498252 539724
rect 498088 539702 498240 539718
rect 501952 539702 502154 539730
rect 495806 539679 495862 539688
rect 502154 539679 502210 539688
rect 505558 539744 505614 539753
rect 508332 539730 508360 543487
rect 509424 543176 509476 543182
rect 509424 543118 509476 543124
rect 508688 541136 508740 541142
rect 508688 541078 508740 541084
rect 508700 539866 508728 541078
rect 509436 539866 509464 543118
rect 513380 543108 513432 543114
rect 513380 543050 513432 543056
rect 512000 543040 512052 543046
rect 512000 542982 512052 542988
rect 510620 542836 510672 542842
rect 510620 542778 510672 542784
rect 510632 539866 510660 542778
rect 511264 541272 511316 541278
rect 511264 541214 511316 541220
rect 511276 539866 511304 541214
rect 512012 539866 512040 542982
rect 513392 539866 513420 543050
rect 515772 542768 515824 542774
rect 515772 542710 515824 542716
rect 514760 542632 514812 542638
rect 514760 542574 514812 542580
rect 513838 541104 513894 541113
rect 513838 541039 513894 541048
rect 513852 539866 513880 541039
rect 514772 539866 514800 542574
rect 515784 539866 515812 542710
rect 520280 539980 520332 539986
rect 520280 539922 520332 539928
rect 517058 539880 517114 539889
rect 508700 539838 509036 539866
rect 509436 539838 509680 539866
rect 510632 539838 510968 539866
rect 511276 539838 511612 539866
rect 512012 539838 512256 539866
rect 513392 539838 513544 539866
rect 513852 539838 514188 539866
rect 514772 539838 514832 539866
rect 515784 539838 516120 539866
rect 517114 539838 517408 539866
rect 517058 539815 517114 539824
rect 516414 539744 516470 539753
rect 505614 539702 505816 539730
rect 508332 539702 508392 539730
rect 505558 539679 505614 539688
rect 516470 539702 516764 539730
rect 518360 539702 518696 539730
rect 516414 539679 516470 539688
rect 493232 539650 493284 539656
rect 518360 539646 518388 539702
rect 518348 539640 518400 539646
rect 518348 539582 518400 539588
rect 519340 539578 519676 539594
rect 519340 539572 519688 539578
rect 519340 539566 519636 539572
rect 519636 539514 519688 539520
rect 519634 539064 519690 539073
rect 519634 538999 519690 539008
rect 519450 531176 519506 531185
rect 519450 531111 519506 531120
rect 479720 500126 480056 500154
rect 479524 498160 479576 498166
rect 479524 498102 479576 498108
rect 479720 496126 479748 500126
rect 480686 499882 480714 500140
rect 480640 499854 480714 499882
rect 481330 499882 481358 500140
rect 481974 499882 482002 500140
rect 481330 499854 481404 499882
rect 480640 497554 480668 499854
rect 481376 499458 481404 499854
rect 481928 499854 482002 499882
rect 483262 499882 483290 500140
rect 483906 499882 483934 500140
rect 484550 499882 484578 500140
rect 485838 499882 485866 500140
rect 486482 499882 486510 500140
rect 487126 499882 487154 500140
rect 483262 499854 483336 499882
rect 481364 499452 481416 499458
rect 481364 499394 481416 499400
rect 480628 497548 480680 497554
rect 480628 497490 480680 497496
rect 481640 496800 481692 496806
rect 481640 496742 481692 496748
rect 479708 496120 479760 496126
rect 479708 496062 479760 496068
rect 479340 486464 479392 486470
rect 479340 486406 479392 486412
rect 479156 483676 479208 483682
rect 479156 483618 479208 483624
rect 478236 268388 478288 268394
rect 478236 268330 478288 268336
rect 478144 227044 478196 227050
rect 478144 226986 478196 226992
rect 480260 62144 480312 62150
rect 480260 62086 480312 62092
rect 476856 28348 476908 28354
rect 476856 28290 476908 28296
rect 476764 18624 476816 18630
rect 476764 18566 476816 18572
rect 480272 16574 480300 62086
rect 481652 16574 481680 496742
rect 481928 475386 481956 499854
rect 483308 493474 483336 499854
rect 483860 499854 483934 499882
rect 484504 499854 484578 499882
rect 485792 499854 485866 499882
rect 486436 499854 486510 499882
rect 487080 499854 487154 499882
rect 488414 499882 488442 500140
rect 489058 499882 489086 500140
rect 489702 499882 489730 500140
rect 490990 499882 491018 500140
rect 491634 499882 491662 500140
rect 492278 499882 492306 500140
rect 488414 499854 488488 499882
rect 483860 498166 483888 499854
rect 483848 498160 483900 498166
rect 483848 498102 483900 498108
rect 484504 496913 484532 499854
rect 485792 499526 485820 499854
rect 485780 499520 485832 499526
rect 485780 499462 485832 499468
rect 486436 497690 486464 499854
rect 486424 497684 486476 497690
rect 486424 497626 486476 497632
rect 484490 496904 484546 496913
rect 484490 496839 484546 496848
rect 486424 496868 486476 496874
rect 486424 496810 486476 496816
rect 484400 494828 484452 494834
rect 484400 494770 484452 494776
rect 483296 493468 483348 493474
rect 483296 493410 483348 493416
rect 481916 475380 481968 475386
rect 481916 475322 481968 475328
rect 483020 63572 483072 63578
rect 483020 63514 483072 63520
rect 483032 16574 483060 63514
rect 484412 16574 484440 494770
rect 485778 281480 485834 281489
rect 485778 281415 485780 281424
rect 485832 281415 485834 281424
rect 485780 281386 485832 281392
rect 486436 35222 486464 496810
rect 487080 231130 487108 499854
rect 488460 496398 488488 499854
rect 489012 499854 489086 499882
rect 489656 499854 489730 499882
rect 490944 499854 491018 499882
rect 491588 499854 491662 499882
rect 492232 499854 492306 499882
rect 493566 499882 493594 500140
rect 494210 499882 494238 500140
rect 494854 499882 494882 500140
rect 493566 499854 493640 499882
rect 489012 497622 489040 499854
rect 489656 498030 489684 499854
rect 489644 498024 489696 498030
rect 489644 497966 489696 497972
rect 489000 497616 489052 497622
rect 489000 497558 489052 497564
rect 489184 497616 489236 497622
rect 489184 497558 489236 497564
rect 488448 496392 488500 496398
rect 488448 496334 488500 496340
rect 488540 493536 488592 493542
rect 488540 493478 488592 493484
rect 487068 231124 487120 231130
rect 487068 231066 487120 231072
rect 486424 35216 486476 35222
rect 486424 35158 486476 35164
rect 488552 16574 488580 493478
rect 480272 16546 480576 16574
rect 481652 16546 481772 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 488552 16546 488856 16574
rect 475384 3732 475436 3738
rect 475384 3674 475436 3680
rect 478144 3664 478196 3670
rect 478144 3606 478196 3612
rect 474188 3392 474240 3398
rect 474188 3334 474240 3340
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3334
rect 478156 480 478184 3606
rect 480548 480 480576 16546
rect 481744 480 481772 16546
rect 484044 480 484072 16546
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 487620 7676 487672 7682
rect 487620 7618 487672 7624
rect 487632 480 487660 7618
rect 488828 480 488856 16546
rect 489196 3466 489224 497558
rect 490944 496874 490972 499854
rect 490932 496868 490984 496874
rect 490932 496810 490984 496816
rect 490564 496392 490616 496398
rect 490564 496334 490616 496340
rect 490576 325650 490604 496334
rect 491300 496120 491352 496126
rect 491300 496062 491352 496068
rect 490564 325644 490616 325650
rect 490564 325586 490616 325592
rect 489920 69080 489972 69086
rect 489920 69022 489972 69028
rect 489932 16574 489960 69022
rect 491312 16574 491340 496062
rect 489932 16546 490696 16574
rect 491312 16546 491524 16574
rect 489184 3460 489236 3466
rect 489184 3402 489236 3408
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490668 354 490696 16546
rect 491300 3732 491352 3738
rect 491300 3674 491352 3680
rect 491312 3534 491340 3674
rect 491300 3528 491352 3534
rect 491300 3470 491352 3476
rect 491496 3482 491524 16546
rect 491588 6186 491616 499854
rect 492232 499390 492260 499854
rect 493612 499390 493640 499854
rect 494164 499854 494238 499882
rect 494808 499854 494882 499882
rect 492220 499384 492272 499390
rect 492220 499326 492272 499332
rect 493600 499384 493652 499390
rect 493600 499326 493652 499332
rect 491944 497548 491996 497554
rect 491944 497490 491996 497496
rect 491576 6180 491628 6186
rect 491576 6122 491628 6128
rect 491956 3738 491984 497490
rect 493324 496868 493376 496874
rect 493324 496810 493376 496816
rect 493336 31074 493364 496810
rect 494164 487830 494192 499854
rect 494808 499254 494836 499854
rect 496142 499746 496170 500140
rect 496786 499882 496814 500140
rect 497430 499882 497458 500140
rect 496096 499718 496170 499746
rect 496740 499854 496814 499882
rect 497384 499854 497458 499882
rect 498718 499882 498746 500140
rect 499362 499882 499390 500140
rect 500006 499882 500034 500140
rect 498718 499854 498792 499882
rect 496096 499633 496124 499718
rect 496082 499624 496138 499633
rect 496082 499559 496138 499568
rect 494796 499248 494848 499254
rect 494796 499190 494848 499196
rect 496096 496913 496124 499559
rect 494702 496904 494758 496913
rect 494702 496839 494758 496848
rect 496082 496904 496138 496913
rect 496082 496839 496138 496848
rect 494152 487824 494204 487830
rect 494152 487766 494204 487772
rect 493324 31068 493376 31074
rect 493324 31010 493376 31016
rect 494716 13122 494744 496839
rect 496740 272542 496768 499854
rect 497384 496874 497412 499854
rect 497372 496868 497424 496874
rect 497372 496810 497424 496816
rect 498200 496188 498252 496194
rect 498200 496130 498252 496136
rect 496728 272536 496780 272542
rect 496728 272478 496780 272484
rect 494704 13116 494756 13122
rect 494704 13058 494756 13064
rect 494704 9104 494756 9110
rect 494704 9046 494756 9052
rect 491944 3732 491996 3738
rect 491944 3674 491996 3680
rect 491496 3454 492352 3482
rect 492324 480 492352 3454
rect 494716 480 494744 9046
rect 495898 3360 495954 3369
rect 495898 3295 495954 3304
rect 495912 480 495940 3295
rect 498212 480 498240 496130
rect 498764 354006 498792 499854
rect 499316 499854 499390 499882
rect 499960 499854 500034 499882
rect 501294 499882 501322 500140
rect 501938 499882 501966 500140
rect 502582 499905 502610 500140
rect 501294 499854 501368 499882
rect 499316 498030 499344 499854
rect 498844 498024 498896 498030
rect 498844 497966 498896 497972
rect 499304 498024 499356 498030
rect 499304 497966 499356 497972
rect 498752 354000 498804 354006
rect 498752 353942 498804 353948
rect 498856 47598 498884 497966
rect 499960 273222 499988 499854
rect 501340 496262 501368 499854
rect 501892 499854 501966 499882
rect 502568 499896 502624 499905
rect 501328 496256 501380 496262
rect 501328 496198 501380 496204
rect 500224 493060 500276 493066
rect 500224 493002 500276 493008
rect 499948 273216 500000 273222
rect 499948 273158 500000 273164
rect 498844 47592 498896 47598
rect 498844 47534 498896 47540
rect 500236 4146 500264 493002
rect 501892 275330 501920 499854
rect 503870 499882 503898 500140
rect 504514 499882 504542 500140
rect 505158 499882 505186 500140
rect 505802 499882 505830 500140
rect 503870 499854 503944 499882
rect 502568 499831 502624 499840
rect 503916 478174 503944 499854
rect 504468 499854 504542 499882
rect 505112 499854 505186 499882
rect 505756 499854 505830 499882
rect 507090 499882 507118 500140
rect 507734 499882 507762 500140
rect 508378 499882 508406 500140
rect 507090 499854 507164 499882
rect 503904 478168 503956 478174
rect 503904 478110 503956 478116
rect 501880 275324 501932 275330
rect 501880 275266 501932 275272
rect 499396 4140 499448 4146
rect 499396 4082 499448 4088
rect 500224 4140 500276 4146
rect 500224 4082 500276 4088
rect 499408 480 499436 4082
rect 502982 3496 503038 3505
rect 504468 3466 504496 499854
rect 505112 493066 505140 499854
rect 505756 499322 505784 499854
rect 505744 499316 505796 499322
rect 505744 499258 505796 499264
rect 506480 498840 506532 498846
rect 506480 498782 506532 498788
rect 505100 493060 505152 493066
rect 505100 493002 505152 493008
rect 502982 3431 503038 3440
rect 504456 3460 504508 3466
rect 502996 480 503024 3431
rect 504456 3402 504508 3408
rect 506492 480 506520 498782
rect 507136 229770 507164 499854
rect 507688 499854 507762 499882
rect 508332 499854 508406 499882
rect 509666 499882 509694 500140
rect 510310 499882 510338 500140
rect 510954 499882 510982 500140
rect 512242 499882 512270 500140
rect 512886 499882 512914 500140
rect 513530 499882 513558 500140
rect 514818 499882 514846 500140
rect 515462 499882 515490 500140
rect 516106 499882 516134 500140
rect 517394 499882 517422 500140
rect 518038 499882 518066 500140
rect 518682 499882 518710 500140
rect 509666 499854 509740 499882
rect 510310 499854 510384 499882
rect 507688 280090 507716 499854
rect 507676 280084 507728 280090
rect 507676 280026 507728 280032
rect 507124 229764 507176 229770
rect 507124 229706 507176 229712
rect 508332 4826 508360 499854
rect 509712 40730 509740 499854
rect 510356 497690 510384 499854
rect 510908 499854 510982 499882
rect 512196 499854 512270 499882
rect 512840 499854 512914 499882
rect 513484 499854 513558 499882
rect 514772 499854 514846 499882
rect 515416 499854 515490 499882
rect 516060 499854 516134 499882
rect 517348 499854 517422 499882
rect 517992 499854 518066 499882
rect 518636 499854 518710 499882
rect 510344 497684 510396 497690
rect 510344 497626 510396 497632
rect 509700 40724 509752 40730
rect 509700 40666 509752 40672
rect 510908 33114 510936 499854
rect 512196 498098 512224 499854
rect 512184 498092 512236 498098
rect 512184 498034 512236 498040
rect 512840 497622 512868 499854
rect 513484 498030 513512 499854
rect 513472 498024 513524 498030
rect 513472 497966 513524 497972
rect 512828 497616 512880 497622
rect 512828 497558 512880 497564
rect 514772 497486 514800 499854
rect 514760 497480 514812 497486
rect 514760 497422 514812 497428
rect 515416 479534 515444 499854
rect 516060 497962 516088 499854
rect 516784 498908 516836 498914
rect 516784 498850 516836 498856
rect 516048 497956 516100 497962
rect 516048 497898 516100 497904
rect 516140 492108 516192 492114
rect 516140 492050 516192 492056
rect 515404 479528 515456 479534
rect 515404 479470 515456 479476
rect 510896 33108 510948 33114
rect 510896 33050 510948 33056
rect 516152 16574 516180 492050
rect 516152 16546 516732 16574
rect 508320 4820 508372 4826
rect 508320 4762 508372 4768
rect 510066 4040 510122 4049
rect 510066 3975 510122 3984
rect 510080 480 510108 3975
rect 513562 3496 513618 3505
rect 516704 3482 516732 16546
rect 516796 3602 516824 498850
rect 517348 497554 517376 499854
rect 517336 497548 517388 497554
rect 517336 497490 517388 497496
rect 516876 496256 516928 496262
rect 516876 496198 516928 496204
rect 516888 193186 516916 496198
rect 516876 193180 516928 193186
rect 516876 193122 516928 193128
rect 517992 4894 518020 499854
rect 518256 499044 518308 499050
rect 518256 498986 518308 498992
rect 518164 498976 518216 498982
rect 518164 498918 518216 498924
rect 517980 4888 518032 4894
rect 517980 4830 518032 4836
rect 518176 3670 518204 498918
rect 518268 106282 518296 498986
rect 518636 153202 518664 499854
rect 519464 276690 519492 531111
rect 519542 530088 519598 530097
rect 519542 530023 519598 530032
rect 519556 281518 519584 530023
rect 519648 491978 519676 538999
rect 519726 529000 519782 529009
rect 519726 528935 519782 528944
rect 519740 504370 519768 528935
rect 520094 518460 520150 518469
rect 520094 518395 520150 518404
rect 519910 505200 519966 505209
rect 519910 505135 519966 505144
rect 519740 504342 519860 504370
rect 519728 500948 519780 500954
rect 519728 500890 519780 500896
rect 519740 500585 519768 500890
rect 519726 500576 519782 500585
rect 519726 500511 519782 500520
rect 519832 498846 519860 504342
rect 519820 498840 519872 498846
rect 519820 498782 519872 498788
rect 519636 491972 519688 491978
rect 519636 491914 519688 491920
rect 519544 281512 519596 281518
rect 519544 281454 519596 281460
rect 519452 276684 519504 276690
rect 519452 276626 519504 276632
rect 518624 153196 518676 153202
rect 518624 153138 518676 153144
rect 518256 106276 518308 106282
rect 518256 106218 518308 106224
rect 519924 14482 519952 505135
rect 520002 503840 520058 503849
rect 520002 503775 520058 503784
rect 520016 490618 520044 503775
rect 520108 496194 520136 518395
rect 520096 496188 520148 496194
rect 520096 496130 520148 496136
rect 520004 490612 520056 490618
rect 520004 490554 520056 490560
rect 519912 14476 519964 14482
rect 519912 14418 519964 14424
rect 518164 3664 518216 3670
rect 518164 3606 518216 3612
rect 516784 3596 516836 3602
rect 516784 3538 516836 3544
rect 516704 3454 517192 3482
rect 513562 3431 513618 3440
rect 513576 480 513604 3431
rect 517164 480 517192 3454
rect 491086 354 491198 480
rect 490668 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520292 354 520320 539922
rect 520384 526629 520412 659806
rect 520370 526620 520426 526629
rect 520370 526555 520426 526564
rect 520476 515545 520504 660350
rect 520556 552084 520608 552090
rect 520556 552026 520608 552032
rect 520568 520169 520596 552026
rect 520646 527368 520702 527377
rect 520646 527303 520702 527312
rect 520554 520160 520610 520169
rect 520554 520095 520610 520104
rect 520554 517576 520610 517585
rect 520554 517511 520610 517520
rect 520462 515536 520518 515545
rect 520462 515471 520518 515480
rect 520370 508940 520426 508949
rect 520370 508875 520426 508884
rect 520384 494834 520412 508875
rect 520372 494828 520424 494834
rect 520372 494770 520424 494776
rect 520568 42090 520596 517511
rect 520660 220114 520688 527303
rect 520752 508745 520780 661642
rect 521660 660000 521712 660006
rect 521660 659942 521712 659948
rect 520830 612368 520886 612377
rect 520830 612303 520886 612312
rect 520738 508736 520794 508745
rect 520738 508671 520794 508680
rect 520738 505744 520794 505753
rect 520738 505679 520794 505688
rect 520752 273970 520780 505679
rect 520844 499458 520872 612303
rect 521014 528592 521070 528601
rect 521014 528527 521070 528536
rect 520922 515672 520978 515681
rect 520922 515607 520978 515616
rect 520832 499452 520884 499458
rect 520832 499394 520884 499400
rect 520936 496126 520964 515607
rect 520924 496120 520976 496126
rect 520924 496062 520976 496068
rect 520740 273964 520792 273970
rect 520740 273906 520792 273912
rect 520648 220108 520700 220114
rect 520648 220050 520700 220056
rect 520556 42084 520608 42090
rect 520556 42026 520608 42032
rect 521028 8974 521056 528527
rect 521106 520296 521162 520305
rect 521106 520231 521162 520240
rect 521120 9042 521148 520231
rect 521672 510241 521700 659942
rect 521750 630728 521806 630737
rect 521750 630663 521806 630672
rect 521764 598942 521792 630663
rect 521752 598936 521804 598942
rect 521752 598878 521804 598884
rect 521750 535528 521806 535537
rect 521750 535463 521806 535472
rect 521658 510232 521714 510241
rect 521658 510167 521714 510176
rect 521764 177342 521792 535463
rect 521856 512825 521884 661710
rect 522028 661088 522080 661094
rect 522028 661030 522080 661036
rect 521934 641744 521990 641753
rect 521934 641679 521990 641688
rect 521948 612377 521976 641679
rect 521934 612368 521990 612377
rect 521934 612303 521990 612312
rect 521934 524648 521990 524657
rect 521934 524583 521990 524592
rect 521842 512816 521898 512825
rect 521842 512751 521898 512760
rect 521842 500984 521898 500993
rect 521842 500919 521898 500928
rect 521856 281382 521884 500919
rect 521948 352578 521976 524583
rect 522040 517449 522068 661030
rect 523684 641028 523736 641034
rect 523684 640970 523736 640976
rect 523696 632058 523724 640970
rect 523684 632052 523736 632058
rect 523684 631994 523736 632000
rect 522120 572008 522172 572014
rect 522120 571950 522172 571956
rect 522026 517440 522082 517449
rect 522026 517375 522082 517384
rect 522026 513768 522082 513777
rect 522026 513703 522082 513712
rect 522040 493338 522068 513703
rect 522132 500857 522160 571950
rect 525076 544406 525104 696934
rect 525064 544400 525116 544406
rect 525064 544342 525116 544348
rect 525064 539708 525116 539714
rect 525064 539650 525116 539656
rect 523040 539572 523092 539578
rect 523040 539514 523092 539520
rect 522302 537024 522358 537033
rect 522302 536959 522358 536968
rect 522210 536344 522266 536353
rect 522210 536279 522266 536288
rect 522224 535702 522252 536279
rect 522212 535696 522264 535702
rect 522212 535638 522264 535644
rect 522210 534304 522266 534313
rect 522210 534239 522266 534248
rect 522118 500848 522174 500857
rect 522118 500783 522174 500792
rect 522224 493406 522252 534239
rect 522316 498914 522344 536959
rect 522948 532704 523000 532710
rect 522948 532646 523000 532652
rect 522960 532409 522988 532646
rect 522946 532400 523002 532409
rect 522946 532335 523002 532344
rect 522946 525872 523002 525881
rect 522946 525807 522948 525816
rect 523000 525807 523002 525816
rect 522948 525778 523000 525784
rect 522946 523152 523002 523161
rect 522946 523087 523002 523096
rect 522960 523054 522988 523087
rect 522948 523048 523000 523054
rect 522948 522990 523000 522996
rect 522486 521928 522542 521937
rect 522486 521863 522542 521872
rect 522394 502480 522450 502489
rect 522394 502415 522450 502424
rect 522408 499050 522436 502415
rect 522396 499044 522448 499050
rect 522396 498986 522448 498992
rect 522500 498982 522528 521863
rect 522946 520976 523002 520985
rect 522946 520911 523002 520920
rect 522960 520674 522988 520911
rect 522948 520668 523000 520674
rect 522948 520610 523000 520616
rect 522856 513256 522908 513262
rect 522854 513224 522856 513233
rect 522908 513224 522910 513233
rect 522854 513159 522910 513168
rect 522946 511184 523002 511193
rect 522946 511119 523002 511128
rect 522960 510746 522988 511119
rect 522948 510740 523000 510746
rect 522948 510682 523000 510688
rect 522578 510640 522634 510649
rect 522578 510575 522634 510584
rect 522488 498976 522540 498982
rect 522488 498918 522540 498924
rect 522304 498908 522356 498914
rect 522304 498850 522356 498856
rect 522212 493400 522264 493406
rect 522212 493342 522264 493348
rect 522028 493332 522080 493338
rect 522028 493274 522080 493280
rect 521936 352572 521988 352578
rect 521936 352514 521988 352520
rect 521844 281376 521896 281382
rect 521844 281318 521896 281324
rect 521752 177336 521804 177342
rect 521752 177278 521804 177284
rect 521108 9036 521160 9042
rect 521108 8978 521160 8984
rect 521016 8968 521068 8974
rect 521016 8910 521068 8916
rect 522592 7614 522620 510575
rect 522946 506560 523002 506569
rect 522946 506495 522948 506504
rect 523000 506495 523002 506504
rect 522948 506466 523000 506472
rect 523052 16574 523080 539514
rect 523684 536852 523736 536858
rect 523684 536794 523736 536800
rect 523696 499390 523724 536794
rect 523684 499384 523736 499390
rect 523684 499326 523736 499332
rect 523052 16546 523816 16574
rect 522580 7608 522632 7614
rect 522580 7550 522632 7556
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523788 354 523816 16546
rect 525076 3602 525104 539650
rect 525156 535696 525208 535702
rect 525156 535638 525208 535644
rect 525168 485790 525196 535638
rect 526456 513262 526484 699654
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 534724 643136 534776 643142
rect 534724 643078 534776 643084
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 527824 640960 527876 640966
rect 527824 640902 527876 640908
rect 527836 525774 527864 640902
rect 534736 532710 534764 643078
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 538864 616888 538916 616894
rect 538864 616830 538916 616836
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 538876 556850 538904 616830
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580172 578196 580224 578202
rect 580172 578138 580224 578144
rect 580184 577697 580212 578138
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580262 564360 580318 564369
rect 580262 564295 580318 564304
rect 538864 556844 538916 556850
rect 538864 556786 538916 556792
rect 580276 554033 580304 564295
rect 580262 554024 580318 554033
rect 580262 553959 580318 553968
rect 540244 542564 540296 542570
rect 540244 542506 540296 542512
rect 534724 532704 534776 532710
rect 534724 532646 534776 532652
rect 536104 525836 536156 525842
rect 536104 525778 536156 525784
rect 527824 525768 527876 525774
rect 527824 525710 527876 525716
rect 534724 523048 534776 523054
rect 534724 522990 534776 522996
rect 530584 520668 530636 520674
rect 530584 520610 530636 520616
rect 526444 513256 526496 513262
rect 526444 513198 526496 513204
rect 526444 510672 526496 510678
rect 526444 510614 526496 510620
rect 526456 498778 526484 510614
rect 527824 506524 527876 506530
rect 527824 506466 527876 506472
rect 526444 498772 526496 498778
rect 526444 498714 526496 498720
rect 526444 497684 526496 497690
rect 526444 497626 526496 497632
rect 525156 485784 525208 485790
rect 525156 485726 525208 485732
rect 525064 3596 525116 3602
rect 525064 3538 525116 3544
rect 526456 3534 526484 497626
rect 527836 16574 527864 506466
rect 530596 113150 530624 520610
rect 534080 486464 534132 486470
rect 534080 486406 534132 486412
rect 530584 113144 530636 113150
rect 530584 113086 530636 113092
rect 534092 16574 534120 486406
rect 534736 233238 534764 522990
rect 534724 233232 534776 233238
rect 534724 233174 534776 233180
rect 527836 16546 527956 16574
rect 534092 16546 534488 16574
rect 527928 3534 527956 16546
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 526444 3528 526496 3534
rect 526444 3470 526496 3476
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 527916 3528 527968 3534
rect 527916 3470 527968 3476
rect 527836 480 527864 3470
rect 531332 480 531360 3538
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534460 354 534488 16546
rect 536116 3602 536144 525778
rect 538864 510740 538916 510746
rect 538864 510682 538916 510688
rect 536104 3596 536156 3602
rect 536104 3538 536156 3544
rect 538876 3534 538904 510682
rect 540256 3670 540284 542506
rect 543004 541204 543056 541210
rect 543004 541146 543056 541152
rect 540980 354000 541032 354006
rect 540980 353942 541032 353948
rect 540992 16574 541020 353942
rect 543016 73166 543044 541146
rect 556160 541068 556212 541074
rect 556160 541010 556212 541016
rect 545120 541000 545172 541006
rect 545120 540942 545172 540948
rect 544384 539776 544436 539782
rect 544384 539718 544436 539724
rect 544396 379506 544424 539718
rect 544384 379500 544436 379506
rect 544384 379442 544436 379448
rect 543004 73160 543056 73166
rect 543004 73102 543056 73108
rect 545132 16574 545160 540942
rect 547880 539912 547932 539918
rect 547880 539854 547932 539860
rect 547892 16574 547920 539854
rect 552020 493468 552072 493474
rect 552020 493410 552072 493416
rect 552032 16574 552060 493410
rect 540992 16546 542032 16574
rect 545132 16546 545528 16574
rect 547892 16546 548656 16574
rect 552032 16546 552704 16574
rect 540244 3664 540296 3670
rect 540244 3606 540296 3612
rect 538404 3528 538456 3534
rect 538404 3470 538456 3476
rect 538864 3528 538916 3534
rect 538864 3470 538916 3476
rect 538416 480 538444 3470
rect 542004 480 542032 16546
rect 545500 480 545528 16546
rect 534878 354 534990 480
rect 534460 326 534990 354
rect 534878 -960 534990 326
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 548628 354 548656 16546
rect 552676 480 552704 16546
rect 556172 480 556200 541010
rect 565820 539844 565872 539850
rect 565820 539786 565872 539792
rect 563060 494760 563112 494766
rect 563060 494702 563112 494708
rect 558184 492040 558236 492046
rect 558184 491982 558236 491988
rect 558196 3398 558224 491982
rect 558184 3392 558236 3398
rect 558184 3334 558236 3340
rect 559748 3392 559800 3398
rect 559748 3334 559800 3340
rect 559760 480 559788 3334
rect 549046 354 549158 480
rect 548628 326 549158 354
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563072 354 563100 494702
rect 565832 16574 565860 539786
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 582380 487892 582432 487898
rect 582380 487834 582432 487840
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 569960 483676 570012 483682
rect 569960 483618 570012 483624
rect 569972 16574 570000 483618
rect 580172 471980 580224 471986
rect 580172 471922 580224 471928
rect 580184 471481 580212 471922
rect 580170 471472 580226 471481
rect 580170 471407 580226 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 579804 431928 579856 431934
rect 579804 431870 579856 431876
rect 579816 431633 579844 431870
rect 579802 431624 579858 431633
rect 579802 431559 579858 431568
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 578884 220856 578936 220862
rect 578884 220798 578936 220804
rect 565832 16546 566872 16574
rect 569972 16546 570368 16574
rect 566844 480 566872 16546
rect 570340 480 570368 16546
rect 573916 3596 573968 3602
rect 573916 3538 573968 3544
rect 573928 480 573956 3538
rect 578896 3534 578924 220798
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580264 109744 580316 109750
rect 580264 109686 580316 109692
rect 580276 86193 580304 109686
rect 580262 86184 580318 86193
rect 580262 86119 580318 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 20596 580224 20602
rect 580172 20538 580224 20544
rect 580184 19825 580212 20538
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 582392 16574 582420 487834
rect 582392 16546 583432 16574
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 582196 3664 582248 3670
rect 582196 3606 582248 3612
rect 578884 3528 578936 3534
rect 578884 3470 578936 3476
rect 579804 3528 579856 3534
rect 579804 3470 579856 3476
rect 577412 3460 577464 3466
rect 577412 3402 577464 3408
rect 577424 480 577452 3402
rect 579816 480 579844 3470
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3606
rect 583404 480 583432 16546
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3238 671200 3294 671256
rect 3330 658144 3386 658200
rect 3330 566888 3386 566944
rect 2962 553832 3018 553888
rect 3606 659912 3662 659968
rect 3606 514800 3662 514856
rect 3514 462576 3570 462632
rect 47950 663176 48006 663232
rect 3422 449520 3478 449576
rect 46846 662904 46902 662960
rect 46754 662768 46810 662824
rect 49974 661816 50030 661872
rect 47950 427080 48006 427136
rect 48042 421232 48098 421288
rect 48134 415384 48190 415440
rect 3146 410488 3202 410544
rect 48594 660048 48650 660104
rect 48594 620064 48650 620120
rect 48502 612720 48558 612776
rect 49330 661544 49386 661600
rect 49054 661272 49110 661328
rect 48962 661000 49018 661056
rect 48870 631760 48926 631816
rect 48686 579128 48742 579184
rect 48778 555736 48834 555792
rect 48962 596672 49018 596728
rect 49238 660320 49294 660376
rect 49054 590824 49110 590880
rect 48870 549888 48926 549944
rect 49422 649304 49478 649360
rect 49238 584976 49294 585032
rect 49146 567432 49202 567488
rect 49882 659640 49938 659696
rect 50158 661680 50214 661736
rect 50066 661408 50122 661464
rect 49606 655152 49662 655208
rect 49514 643456 49570 643512
rect 49422 561584 49478 561640
rect 49330 544040 49386 544096
rect 49422 532344 49478 532400
rect 48870 497256 48926 497312
rect 48778 468016 48834 468072
rect 48318 444624 48374 444680
rect 48318 438812 48320 438832
rect 48320 438812 48372 438832
rect 48372 438812 48374 438832
rect 48318 438776 48374 438812
rect 48226 409536 48282 409592
rect 3422 397432 3478 397488
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3514 306176 3570 306232
rect 3606 293120 3662 293176
rect 48318 392012 48374 392048
rect 48318 391992 48320 392012
rect 48320 391992 48372 392012
rect 48372 391992 48374 392012
rect 48318 386144 48374 386200
rect 48226 374448 48282 374504
rect 48134 368600 48190 368656
rect 48042 362752 48098 362808
rect 47950 351056 48006 351112
rect 47858 345208 47914 345264
rect 47858 281288 47914 281344
rect 47950 281152 48006 281208
rect 46846 280608 46902 280664
rect 48134 280472 48190 280528
rect 46754 280064 46810 280120
rect 48686 298424 48742 298480
rect 48778 292576 48834 292632
rect 46570 279928 46626 279984
rect 3146 254088 3202 254144
rect 2778 149776 2834 149832
rect 3514 241032 3570 241088
rect 3514 224168 3570 224224
rect 3422 97552 3478 97608
rect 3422 84632 3478 84688
rect 3698 201864 3754 201920
rect 3790 188808 3846 188864
rect 3606 136720 3662 136776
rect 3514 58520 3570 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 24214 8880 24270 8936
rect 42798 226888 42854 226944
rect 50250 659640 50306 659696
rect 49606 573280 49662 573336
rect 50434 659776 50490 659832
rect 50526 637472 50582 637528
rect 49606 503104 49662 503160
rect 49514 491408 49570 491464
rect 48962 473864 49018 473920
rect 49146 432928 49202 432984
rect 49422 397840 49478 397896
rect 49422 380296 49478 380352
rect 49422 327664 49478 327720
rect 49330 321816 49386 321872
rect 49238 315968 49294 316024
rect 49146 304272 49202 304328
rect 49422 281016 49478 281072
rect 48962 224304 49018 224360
rect 49606 485560 49662 485616
rect 49606 484336 49662 484392
rect 49790 456356 49792 456376
rect 49792 456356 49844 456376
rect 49844 456356 49846 456376
rect 49790 456320 49846 456356
rect 50710 625912 50766 625968
rect 51078 538192 51134 538248
rect 50986 526496 51042 526552
rect 50894 520648 50950 520704
rect 50802 462168 50858 462224
rect 50710 456320 50766 456376
rect 50618 450472 50674 450528
rect 51446 660592 51502 660648
rect 51170 514800 51226 514856
rect 51262 508952 51318 509008
rect 51354 450472 51410 450528
rect 71778 663040 71834 663096
rect 51814 607144 51870 607200
rect 254766 658144 254822 658200
rect 254582 652296 254638 652352
rect 254306 646448 254362 646504
rect 254306 640600 254362 640656
rect 254398 617208 254454 617264
rect 254490 611380 254546 611416
rect 254490 611360 254492 611380
rect 254492 611360 254544 611380
rect 254544 611360 254546 611380
rect 254214 605512 254270 605568
rect 254674 634752 254730 634808
rect 254674 628904 254730 628960
rect 254674 623056 254730 623112
rect 254490 593816 254546 593872
rect 254582 587988 254638 588024
rect 254582 587968 254584 587988
rect 254584 587968 254636 587988
rect 254636 587968 254638 587988
rect 253938 582120 253994 582176
rect 254214 576272 254270 576328
rect 253938 570424 253994 570480
rect 254582 564576 254638 564632
rect 254582 558728 254638 558784
rect 254582 552880 254638 552936
rect 254582 547032 254638 547088
rect 254858 599664 254914 599720
rect 254398 541184 254454 541240
rect 254582 535336 254638 535392
rect 254582 529488 254638 529544
rect 254306 523640 254362 523696
rect 254582 517812 254638 517848
rect 254582 517792 254584 517812
rect 254584 517792 254636 517812
rect 254636 517792 254638 517812
rect 254398 511944 254454 512000
rect 254306 506096 254362 506152
rect 254582 500248 254638 500304
rect 254582 494400 254638 494456
rect 254582 488572 254638 488608
rect 254582 488552 254584 488572
rect 254584 488552 254636 488572
rect 254636 488552 254638 488572
rect 254582 482704 254638 482760
rect 254214 476856 254270 476912
rect 254582 471008 254638 471064
rect 254582 465160 254638 465216
rect 254582 459312 254638 459368
rect 254306 453464 254362 453520
rect 254674 447616 254730 447672
rect 254398 441788 254454 441824
rect 254398 441768 254400 441788
rect 254400 441768 254452 441788
rect 254452 441768 254454 441788
rect 254398 435920 254454 435976
rect 254582 430072 254638 430128
rect 254582 424224 254638 424280
rect 254582 418376 254638 418432
rect 254582 412528 254638 412584
rect 254582 406680 254638 406736
rect 51446 403688 51502 403744
rect 254030 400832 254086 400888
rect 254398 383288 254454 383344
rect 254122 377440 254178 377496
rect 253938 359896 253994 359952
rect 51446 356904 51502 356960
rect 254214 354048 254270 354104
rect 254490 348200 254546 348256
rect 254674 394984 254730 395040
rect 254674 389172 254676 389192
rect 254676 389172 254728 389192
rect 254728 389172 254730 389192
rect 254674 389136 254730 389172
rect 254674 371592 254730 371648
rect 254674 365764 254730 365800
rect 254674 365744 254676 365764
rect 254676 365744 254728 365764
rect 254728 365744 254730 365764
rect 254582 342352 254638 342408
rect 51538 339360 51594 339416
rect 51446 281968 51502 282024
rect 254398 336504 254454 336560
rect 51722 333512 51778 333568
rect 51630 310120 51686 310176
rect 51630 281832 51686 281888
rect 51538 280880 51594 280936
rect 52090 286456 52146 286512
rect 51722 280744 51778 280800
rect 59358 279384 59414 279440
rect 54574 278704 54630 278760
rect 55862 223488 55918 223544
rect 57058 217368 57114 217424
rect 57150 209208 57206 209264
rect 57334 205128 57390 205184
rect 57334 201048 57390 201104
rect 57334 196968 57390 197024
rect 57334 192924 57336 192944
rect 57336 192924 57388 192944
rect 57388 192924 57390 192944
rect 57334 192888 57390 192924
rect 57334 188808 57390 188864
rect 56690 184728 56746 184784
rect 56690 180648 56746 180704
rect 57334 176604 57336 176624
rect 57336 176604 57388 176624
rect 57388 176604 57390 176624
rect 57334 176568 57390 176604
rect 57242 172488 57298 172544
rect 57334 168408 57390 168464
rect 55862 164328 55918 164384
rect 57058 160248 57114 160304
rect 57058 156168 57114 156224
rect 57334 152088 57390 152144
rect 57334 148008 57390 148064
rect 57334 143928 57390 143984
rect 57426 139848 57482 139904
rect 57334 135768 57390 135824
rect 57518 123528 57574 123584
rect 57610 107208 57666 107264
rect 57702 103128 57758 103184
rect 57794 86808 57850 86864
rect 58898 127608 58954 127664
rect 58806 119448 58862 119504
rect 58714 111288 58770 111344
rect 59082 90888 59138 90944
rect 58990 82728 59046 82784
rect 57886 78648 57942 78704
rect 59266 99048 59322 99104
rect 59450 115368 59506 115424
rect 59358 70488 59414 70544
rect 59726 225528 59782 225584
rect 59726 94968 59782 95024
rect 59634 74568 59690 74624
rect 59542 66408 59598 66464
rect 59174 62328 59230 62384
rect 53746 4800 53802 4856
rect 222842 215600 222898 215656
rect 60554 213832 60610 213888
rect 222290 212744 222346 212800
rect 223210 209888 223266 209944
rect 222934 207032 222990 207088
rect 222842 204176 222898 204232
rect 223026 201320 223082 201376
rect 222934 198464 222990 198520
rect 223486 195608 223542 195664
rect 223486 192752 223542 192808
rect 223486 189896 223542 189952
rect 223486 187040 223542 187096
rect 222290 184204 222346 184240
rect 222290 184184 222292 184204
rect 222292 184184 222344 184204
rect 222344 184184 222346 184204
rect 223486 181328 223542 181384
rect 222658 178472 222714 178528
rect 222658 175616 222714 175672
rect 222382 172760 222438 172816
rect 222474 169904 222530 169960
rect 222934 167048 222990 167104
rect 223486 164192 223542 164248
rect 223026 161336 223082 161392
rect 222934 158480 222990 158536
rect 223486 155624 223542 155680
rect 222658 152768 222714 152824
rect 222566 147092 222568 147112
rect 222568 147092 222620 147112
rect 222620 147092 222622 147112
rect 222566 147056 222622 147092
rect 223210 149912 223266 149968
rect 223486 144200 223542 144256
rect 223486 141344 223542 141400
rect 222934 138488 222990 138544
rect 222842 135632 222898 135688
rect 222658 132776 222714 132832
rect 223026 129920 223082 129976
rect 222842 127064 222898 127120
rect 222290 124208 222346 124264
rect 223486 121352 223542 121408
rect 223486 118496 223542 118552
rect 223486 115640 223542 115696
rect 222198 112784 222254 112840
rect 223486 109928 223542 109984
rect 222658 107072 222714 107128
rect 222842 104216 222898 104272
rect 223486 101360 223542 101416
rect 223026 98504 223082 98560
rect 223118 95648 223174 95704
rect 223486 92792 223542 92848
rect 223486 89936 223542 89992
rect 223210 87080 223266 87136
rect 223210 84224 223266 84280
rect 223486 81388 223542 81424
rect 223486 81368 223488 81388
rect 223488 81368 223540 81388
rect 223540 81368 223542 81388
rect 222474 78548 222476 78568
rect 222476 78548 222528 78568
rect 222528 78548 222530 78568
rect 222474 78512 222530 78548
rect 222198 75692 222200 75712
rect 222200 75692 222252 75712
rect 222252 75692 222254 75712
rect 222198 75656 222254 75692
rect 254582 331472 254638 331528
rect 254214 330656 254270 330712
rect 254490 324808 254546 324864
rect 254306 318960 254362 319016
rect 254214 307264 254270 307320
rect 254398 289720 254454 289776
rect 254306 283872 254362 283928
rect 254674 313112 254730 313168
rect 254674 301416 254730 301472
rect 254674 295568 254730 295624
rect 222198 72800 222254 72856
rect 223486 69944 223542 70000
rect 223486 67088 223542 67144
rect 257618 227024 257674 227080
rect 222842 64232 222898 64288
rect 165618 61512 165674 61568
rect 126978 61376 127034 61432
rect 92478 24112 92534 24168
rect 71502 7520 71558 7576
rect 67914 6160 67970 6216
rect 129738 55800 129794 55856
rect 136638 59880 136694 59936
rect 147678 57160 147734 57216
rect 144734 5072 144790 5128
rect 162490 3304 162546 3360
rect 186318 39208 186374 39264
rect 183742 3440 183798 3496
rect 254674 4936 254730 4992
rect 272522 542816 272578 542872
rect 278778 629992 278834 630048
rect 278686 610000 278742 610056
rect 279974 660456 280030 660512
rect 300122 700304 300178 700360
rect 310518 661408 310574 661464
rect 310058 642232 310114 642288
rect 307482 640600 307538 640656
rect 304170 640464 304226 640520
rect 308586 639376 308642 639432
rect 285402 639240 285458 639296
rect 288254 639240 288310 639296
rect 289634 639240 289690 639296
rect 290922 639240 290978 639296
rect 292026 639240 292082 639296
rect 293130 639240 293186 639296
rect 298466 639240 298522 639296
rect 303434 600616 303490 600672
rect 301410 600480 301466 600536
rect 280158 559544 280214 559600
rect 281630 573280 281686 573336
rect 282918 563624 282974 563680
rect 287150 580216 287206 580272
rect 292670 587152 292726 587208
rect 289818 555328 289874 555384
rect 299294 598848 299350 598904
rect 300674 600072 300730 600128
rect 299386 589872 299442 589928
rect 300582 580352 300638 580408
rect 300674 578856 300730 578912
rect 300858 582936 300914 582992
rect 298098 551384 298154 551440
rect 297086 543360 297142 543416
rect 297454 543088 297510 543144
rect 283470 542816 283526 542872
rect 297086 542816 297142 542872
rect 296902 542680 296958 542736
rect 287886 539688 287942 539744
rect 289358 539688 289414 539744
rect 290830 539688 290886 539744
rect 283378 539552 283434 539608
rect 286138 539552 286194 539608
rect 287610 539552 287666 539608
rect 288622 539552 288678 539608
rect 290738 539552 290794 539608
rect 291566 539552 291622 539608
rect 300398 543224 300454 543280
rect 301134 542816 301190 542872
rect 304722 600616 304778 600672
rect 306194 600616 306250 600672
rect 304998 543360 305054 543416
rect 305550 542952 305606 543008
rect 307022 597624 307078 597680
rect 311898 561176 311954 561232
rect 309322 556688 309378 556744
rect 306378 543632 306434 543688
rect 307022 543496 307078 543552
rect 312266 543088 312322 543144
rect 308402 542544 308458 542600
rect 309966 542544 310022 542600
rect 311438 542544 311494 542600
rect 308678 542408 308734 542464
rect 309414 542408 309470 542464
rect 311070 542408 311126 542464
rect 293038 539552 293094 539608
rect 294510 539552 294566 539608
rect 295982 539552 296038 539608
rect 317510 543632 317566 543688
rect 320178 537308 320234 537364
rect 320086 510788 320142 510844
rect 282182 281424 282238 281480
rect 282182 280880 282238 280936
rect 287334 280764 287390 280800
rect 287334 280744 287336 280764
rect 287336 280744 287388 280764
rect 287388 280744 287390 280764
rect 296074 331336 296130 331392
rect 295982 180240 296038 180296
rect 295982 160792 296038 160848
rect 296074 148824 296130 148880
rect 295982 142840 296038 142896
rect 297362 329704 297418 329760
rect 297086 320184 297142 320240
rect 296994 303864 297050 303920
rect 296994 301144 297050 301200
rect 296810 208664 296866 208720
rect 296810 205692 296866 205728
rect 296810 205672 296812 205692
rect 296812 205672 296864 205692
rect 296864 205672 296866 205692
rect 296810 186260 296812 186280
rect 296812 186260 296864 186280
rect 296864 186260 296866 186280
rect 296810 186224 296866 186260
rect 296810 169788 296866 169824
rect 296810 169768 296812 169788
rect 296812 169768 296864 169788
rect 296864 169768 296866 169788
rect 296810 151836 296866 151872
rect 296810 151816 296812 151836
rect 296812 151816 296864 151836
rect 296864 151816 296866 151836
rect 296810 132404 296812 132424
rect 296812 132404 296864 132424
rect 296864 132404 296866 132424
rect 296810 132368 296866 132404
rect 296810 129376 296866 129432
rect 296810 114452 296812 114472
rect 296812 114452 296864 114472
rect 296864 114452 296866 114472
rect 296810 114416 296866 114452
rect 296994 102448 297050 102504
rect 297178 318824 297234 318880
rect 297270 306584 297326 306640
rect 297454 328344 297510 328400
rect 297546 326304 297602 326360
rect 297730 324944 297786 325000
rect 297822 323584 297878 323640
rect 297730 317464 297786 317520
rect 297730 316104 297786 316160
rect 297914 314744 297970 314800
rect 297914 312704 297970 312760
rect 298006 311344 298062 311400
rect 297730 296384 297786 296440
rect 298006 305224 298062 305280
rect 298006 302504 298062 302560
rect 297914 299104 297970 299160
rect 297822 295024 297878 295080
rect 298006 291624 298062 291680
rect 297914 290264 297970 290320
rect 298006 288904 298062 288960
rect 298006 287544 298062 287600
rect 297638 284144 297694 284200
rect 297362 109928 297418 109984
rect 297546 216688 297602 216744
rect 297454 103944 297510 104000
rect 297546 99456 297602 99512
rect 297730 192208 297786 192264
rect 297730 189216 297786 189272
rect 297914 285504 297970 285560
rect 297914 217640 297970 217696
rect 297914 216144 297970 216200
rect 297914 214648 297970 214704
rect 297914 213152 297970 213208
rect 297914 211656 297970 211712
rect 297914 210160 297970 210216
rect 297914 207168 297970 207224
rect 297914 204176 297970 204232
rect 297914 202680 297970 202736
rect 297914 201184 297970 201240
rect 297914 199688 297970 199744
rect 297914 198192 297970 198248
rect 297914 196696 297970 196752
rect 297914 195200 297970 195256
rect 297914 193704 297970 193760
rect 297914 190712 297970 190768
rect 297914 187720 297970 187776
rect 297914 184728 297970 184784
rect 297914 183232 297970 183288
rect 297914 181736 297970 181792
rect 297914 178744 297970 178800
rect 297914 177248 297970 177304
rect 297914 175752 297970 175808
rect 297914 174256 297970 174312
rect 297914 172760 297970 172816
rect 297914 171264 297970 171320
rect 297914 168272 297970 168328
rect 297914 166776 297970 166832
rect 297914 165280 297970 165336
rect 297914 163784 297970 163840
rect 297914 162288 297970 162344
rect 297914 159296 297970 159352
rect 297914 157800 297970 157856
rect 297914 156304 297970 156360
rect 297914 154808 297970 154864
rect 297914 153312 297970 153368
rect 297914 150320 297970 150376
rect 297914 147328 297970 147384
rect 297914 145832 297970 145888
rect 297914 144336 297970 144392
rect 297914 141344 297970 141400
rect 297914 139848 297970 139904
rect 297914 138352 297970 138408
rect 297914 136856 297970 136912
rect 297914 135360 297970 135416
rect 297914 133864 297970 133920
rect 297914 130872 297970 130928
rect 297914 127880 297970 127936
rect 297914 126384 297970 126440
rect 297914 124888 297970 124944
rect 297914 123392 297970 123448
rect 297914 121896 297970 121952
rect 297914 120400 297970 120456
rect 297914 118904 297970 118960
rect 297914 117408 297970 117464
rect 297914 115912 297970 115968
rect 297914 112920 297970 112976
rect 297822 96464 297878 96520
rect 297638 94968 297694 95024
rect 297086 91976 297142 92032
rect 298098 282376 298154 282432
rect 298742 308624 298798 308680
rect 298650 281424 298706 281480
rect 298742 97960 298798 98016
rect 298926 111424 298982 111480
rect 299018 108432 299074 108488
rect 299110 106936 299166 106992
rect 299202 105440 299258 105496
rect 299386 311344 299442 311400
rect 299662 322224 299718 322280
rect 299570 297744 299626 297800
rect 299570 282784 299626 282840
rect 305182 331200 305238 331256
rect 316130 331336 316186 331392
rect 319350 508292 319406 508328
rect 319350 508272 319352 508292
rect 319352 508272 319404 508292
rect 319404 508272 319406 508292
rect 319350 506524 319406 506560
rect 319350 506504 319352 506524
rect 319352 506504 319404 506524
rect 319404 506504 319406 506524
rect 320086 506028 320142 506084
rect 320362 509428 320418 509484
rect 320270 508104 320272 508124
rect 320272 508104 320324 508124
rect 320324 508104 320326 508124
rect 320270 508068 320326 508104
rect 320270 507388 320326 507444
rect 320270 505348 320326 505404
rect 320454 505280 320510 505336
rect 322110 534928 322166 534984
rect 321650 532208 321706 532264
rect 322110 528128 322166 528184
rect 322294 525680 322350 525736
rect 322110 524592 322166 524648
rect 322294 524456 322350 524512
rect 322202 522280 322258 522336
rect 322018 520648 322074 520704
rect 322570 536152 322626 536208
rect 322478 535220 322534 535256
rect 322478 535200 322480 535220
rect 322480 535200 322532 535220
rect 322532 535200 322534 535220
rect 322846 533976 322902 534032
rect 322478 533296 322534 533352
rect 322754 532344 322810 532400
rect 322478 531276 322534 531312
rect 322478 531256 322480 531276
rect 322480 531256 322532 531276
rect 322532 531256 322534 531276
rect 322570 530168 322626 530224
rect 322478 529760 322534 529816
rect 322478 528400 322534 528456
rect 322846 528808 322902 528864
rect 322570 527040 322626 527096
rect 322478 526768 322534 526824
rect 322662 523232 322718 523288
rect 322478 523096 322534 523152
rect 322570 522144 322626 522200
rect 322478 520512 322534 520568
rect 322202 519560 322258 519616
rect 321650 519424 321706 519480
rect 322294 517928 322350 517984
rect 321742 517792 321798 517848
rect 322294 515344 322350 515400
rect 322294 513460 322350 513496
rect 322294 513440 322296 513460
rect 322296 513440 322348 513460
rect 322348 513440 322350 513460
rect 321742 512624 321798 512680
rect 322202 512644 322258 512680
rect 322202 512624 322204 512644
rect 322204 512624 322256 512644
rect 322256 512624 322258 512644
rect 321558 511284 321614 511320
rect 321558 511264 321560 511284
rect 321560 511264 321612 511284
rect 321612 511264 321614 511284
rect 321650 509632 321706 509688
rect 321558 504600 321614 504656
rect 322202 512080 322258 512136
rect 321650 349696 321706 349752
rect 322386 506776 322442 506832
rect 322478 504464 322534 504520
rect 322478 503512 322534 503568
rect 322478 502424 322534 502480
rect 322754 517384 322810 517440
rect 322846 516704 322902 516760
rect 322846 515480 322902 515536
rect 322754 514120 322810 514176
rect 324226 518880 324282 518936
rect 322202 335960 322258 336016
rect 329102 547032 329158 547088
rect 331218 516704 331274 516760
rect 331954 641824 332010 641880
rect 337934 530576 337990 530632
rect 345846 541048 345902 541104
rect 348514 497120 348570 497176
rect 350078 496848 350134 496904
rect 348974 331472 349030 331528
rect 350078 327664 350134 327720
rect 350262 329024 350318 329080
rect 349802 315968 349858 316024
rect 299294 100952 299350 101008
rect 298834 93472 298890 93528
rect 298006 90480 298062 90536
rect 297178 85992 297234 86048
rect 296810 84496 296866 84552
rect 297178 77016 297234 77072
rect 296810 72528 296866 72584
rect 297178 68040 297234 68096
rect 349802 312160 349858 312216
rect 349802 290808 349858 290864
rect 349802 286320 349858 286376
rect 350078 310800 350134 310856
rect 350354 303864 350410 303920
rect 341062 147464 341118 147520
rect 340142 145288 340198 145344
rect 340050 129920 340106 129976
rect 299386 88984 299442 89040
rect 298006 87488 298062 87544
rect 297914 83000 297970 83056
rect 297914 81504 297970 81560
rect 298006 80028 298062 80064
rect 298006 80008 298008 80028
rect 298008 80008 298060 80028
rect 298060 80008 298062 80028
rect 297546 78512 297602 78568
rect 298006 75520 298062 75576
rect 298006 74024 298062 74080
rect 297730 71032 297786 71088
rect 298006 69536 298062 69592
rect 297546 66544 297602 66600
rect 297362 65048 297418 65104
rect 297914 63552 297970 63608
rect 298006 62076 298062 62112
rect 298006 62056 298008 62076
rect 298008 62056 298060 62076
rect 298060 62056 298062 62076
rect 297270 3576 297326 3632
rect 300766 3576 300822 3632
rect 317418 60016 317474 60072
rect 340878 140936 340934 140992
rect 340234 138760 340290 138816
rect 340326 119176 340382 119232
rect 340418 110472 340474 110528
rect 340510 75656 340566 75712
rect 340970 121352 341026 121408
rect 343086 143112 343142 143168
rect 342442 136584 342498 136640
rect 342258 134408 342314 134464
rect 341154 132232 341210 132288
rect 341338 114824 341394 114880
rect 341246 112648 341302 112704
rect 341430 103944 341486 104000
rect 341522 101768 341578 101824
rect 341614 99592 341670 99648
rect 341706 97416 341762 97472
rect 342350 117000 342406 117056
rect 342350 108296 342406 108352
rect 342350 106120 342406 106176
rect 342350 93064 342406 93120
rect 342350 79328 342406 79384
rect 342350 79192 342406 79248
rect 342534 127880 342590 127936
rect 342350 62600 342406 62656
rect 342626 125704 342682 125760
rect 342718 123528 342774 123584
rect 342810 90888 342866 90944
rect 342902 88712 342958 88768
rect 342994 69128 343050 69184
rect 342994 66952 343050 67008
rect 342994 64776 343050 64832
rect 343178 86536 343234 86592
rect 329194 3576 329250 3632
rect 353298 530576 353354 530632
rect 353298 529896 353354 529952
rect 353574 529896 353630 529952
rect 351274 497256 351330 497312
rect 350998 324944 351054 325000
rect 350906 314064 350962 314120
rect 350906 291624 350962 291680
rect 350814 280744 350870 280800
rect 351090 317464 351146 317520
rect 351090 307944 351146 308000
rect 351918 326304 351974 326360
rect 351918 321544 351974 321600
rect 352010 318824 352066 318880
rect 351458 305224 351514 305280
rect 351918 301824 351974 301880
rect 351918 300464 351974 300520
rect 351366 299104 351422 299160
rect 351366 291660 351368 291680
rect 351368 291660 351420 291680
rect 351420 291660 351422 291680
rect 351366 291624 351422 291660
rect 351274 288224 351330 288280
rect 352102 297744 352158 297800
rect 352010 294344 352066 294400
rect 352102 285504 352158 285560
rect 352378 323584 352434 323640
rect 352286 296384 352342 296440
rect 352286 292984 352342 293040
rect 352194 282784 352250 282840
rect 352562 306584 352618 306640
rect 352470 284144 352526 284200
rect 352838 309984 352894 310040
rect 355230 497528 355286 497584
rect 358818 661272 358874 661328
rect 401598 661308 401600 661328
rect 401600 661308 401652 661328
rect 401652 661308 401654 661328
rect 401598 661272 401654 661308
rect 356702 503240 356758 503296
rect 356610 499432 356666 499488
rect 357070 550296 357126 550352
rect 357530 548936 357586 548992
rect 357438 547712 357494 547768
rect 357438 546216 357494 546272
rect 357438 544720 357494 544776
rect 357438 539144 357494 539200
rect 357438 536732 357440 536752
rect 357440 536732 357492 536752
rect 357492 536732 357494 536752
rect 357438 536696 357494 536732
rect 357438 535336 357494 535392
rect 357530 535200 357586 535256
rect 357530 533452 357586 533488
rect 357530 533432 357532 533452
rect 357532 533432 357584 533452
rect 357584 533432 357586 533452
rect 357438 532344 357494 532400
rect 357530 531800 357586 531856
rect 357438 529488 357494 529544
rect 357438 527076 357440 527096
rect 357440 527076 357492 527096
rect 357492 527076 357494 527096
rect 357438 527040 357494 527076
rect 357530 526360 357586 526416
rect 357438 523640 357494 523696
rect 357714 543496 357770 543552
rect 357714 539280 357770 539336
rect 357622 521600 357678 521656
rect 357438 519560 357494 519616
rect 357438 518744 357494 518800
rect 357530 517540 357586 517576
rect 357530 517520 357532 517540
rect 357532 517520 357584 517540
rect 357584 517520 357586 517540
rect 357438 517420 357440 517440
rect 357440 517420 357492 517440
rect 357492 517420 357494 517440
rect 357438 517384 357494 517420
rect 357438 514700 357440 514720
rect 357440 514700 357492 514720
rect 357492 514700 357494 514720
rect 357438 514664 357494 514700
rect 357530 513440 357586 513496
rect 357438 512760 357494 512816
rect 357438 511400 357494 511456
rect 357438 510448 357494 510504
rect 357438 508952 357494 509008
rect 357438 507320 357494 507376
rect 357438 506404 357440 506424
rect 357440 506404 357492 506424
rect 357492 506404 357494 506424
rect 357438 506368 357494 506404
rect 357438 504600 357494 504656
rect 357438 501880 357494 501936
rect 357622 505824 357678 505880
rect 357898 544992 357954 545048
rect 358082 543496 358138 543552
rect 357898 536560 357954 536616
rect 357898 534520 357954 534576
rect 358266 538056 358322 538112
rect 358450 542272 358506 542328
rect 358542 540912 358598 540968
rect 358726 548800 358782 548856
rect 358634 537920 358690 537976
rect 358358 533432 358414 533488
rect 358358 528536 358414 528592
rect 358174 528264 358230 528320
rect 357806 524592 357862 524648
rect 357806 523776 357862 523832
rect 358082 519696 358138 519752
rect 358174 515072 358230 515128
rect 357898 511536 357954 511592
rect 357990 508680 358046 508736
rect 358266 503648 358322 503704
rect 358634 532752 358690 532808
rect 358542 522416 358598 522472
rect 358450 507728 358506 507784
rect 358910 543360 358966 543416
rect 358818 510040 358874 510096
rect 359094 522280 359150 522336
rect 359554 524728 359610 524784
rect 359186 520920 359242 520976
rect 359002 513304 359058 513360
rect 359370 497800 359426 497856
rect 360014 599528 360070 599584
rect 360014 552064 360070 552120
rect 368938 642096 368994 642152
rect 361946 639376 362002 639432
rect 362498 639512 362554 639568
rect 362590 639376 362646 639432
rect 364062 639376 364118 639432
rect 369490 641688 369546 641744
rect 378046 641008 378102 641064
rect 378874 640328 378930 640384
rect 382186 641824 382242 641880
rect 379518 640872 379574 640928
rect 398194 642232 398250 642288
rect 397090 641960 397146 642016
rect 398194 641688 398250 641744
rect 399206 641688 399262 641744
rect 380162 639648 380218 639704
rect 368110 639376 368166 639432
rect 369674 639396 369730 639432
rect 382922 639512 382978 639568
rect 369674 639376 369676 639396
rect 369676 639376 369728 639396
rect 369728 639376 369730 639396
rect 380898 639376 380954 639432
rect 391294 639376 391350 639432
rect 361578 593136 361634 593192
rect 362314 593272 362370 593328
rect 361854 551928 361910 551984
rect 364522 581576 364578 581632
rect 367282 568520 367338 568576
rect 368478 551656 368534 551712
rect 370134 564984 370190 565040
rect 370042 563080 370098 563136
rect 369858 554104 369914 554160
rect 371238 555464 371294 555520
rect 376114 597624 376170 597680
rect 376942 565800 376998 565856
rect 376758 552608 376814 552664
rect 378414 571920 378470 571976
rect 379610 577496 379666 577552
rect 378322 562400 378378 562456
rect 378230 558320 378286 558376
rect 383290 598168 383346 598224
rect 382370 563624 382426 563680
rect 386602 581576 386658 581632
rect 389270 579536 389326 579592
rect 388534 569336 388590 569392
rect 388442 564440 388498 564496
rect 391202 595448 391258 595504
rect 392030 563624 392086 563680
rect 394790 575456 394846 575512
rect 397458 581712 397514 581768
rect 397642 550060 397644 550080
rect 397644 550060 397696 550080
rect 397696 550060 397698 550080
rect 397642 550024 397698 550060
rect 359738 500792 359794 500848
rect 399758 536968 399814 537024
rect 399850 536560 399906 536616
rect 399574 536288 399630 536344
rect 399482 507320 399538 507376
rect 399482 501608 399538 501664
rect 360014 499704 360070 499760
rect 360658 499840 360714 499896
rect 360474 497664 360530 497720
rect 362958 499876 362960 499896
rect 362960 499876 363012 499896
rect 363012 499876 363014 499896
rect 362958 499840 363014 499876
rect 362590 497392 362646 497448
rect 365166 499840 365222 499896
rect 365810 499432 365866 499488
rect 368386 499840 368442 499896
rect 367742 499432 367798 499488
rect 370962 499840 371018 499896
rect 371606 499840 371662 499896
rect 369030 498072 369086 498128
rect 369030 497256 369086 497312
rect 374826 499296 374882 499352
rect 376390 499840 376446 499896
rect 376114 498072 376170 498128
rect 377402 499840 377458 499896
rect 376758 499432 376814 499488
rect 380622 499840 380678 499896
rect 381266 499840 381322 499896
rect 382554 499840 382610 499896
rect 382554 497120 382610 497176
rect 385774 499840 385830 499896
rect 385130 499704 385186 499760
rect 386418 498072 386474 498128
rect 387706 499840 387762 499896
rect 387062 497936 387118 497992
rect 390282 499840 390338 499896
rect 385774 497800 385830 497856
rect 385130 497664 385186 497720
rect 391570 497528 391626 497584
rect 392858 499840 392914 499896
rect 395434 499840 395490 499896
rect 400126 541524 400182 541580
rect 399942 533160 399998 533216
rect 400402 526564 400458 526620
rect 400310 517724 400366 517780
rect 401138 551520 401194 551576
rect 400954 539280 401010 539336
rect 401046 538056 401102 538112
rect 400770 532480 400826 532536
rect 400678 526632 400734 526688
rect 401138 522960 401194 523016
rect 400494 514800 400550 514856
rect 400218 511604 400274 511660
rect 398654 497936 398710 497992
rect 401598 535336 401654 535392
rect 401598 533568 401654 533624
rect 401598 530032 401654 530088
rect 401598 528808 401654 528864
rect 401598 528128 401654 528184
rect 401598 526088 401654 526144
rect 401598 525408 401654 525464
rect 401598 524864 401654 524920
rect 401598 524048 401654 524104
rect 401598 521736 401654 521792
rect 401598 520784 401654 520840
rect 401598 519968 401654 520024
rect 401782 543088 401838 543144
rect 401782 541728 401838 541784
rect 401782 530304 401838 530360
rect 401782 528944 401838 529000
rect 401782 528536 401838 528592
rect 401690 517384 401746 517440
rect 401598 516296 401654 516352
rect 401690 515888 401746 515944
rect 401690 513848 401746 513904
rect 401598 506404 401600 506424
rect 401600 506404 401652 506424
rect 401652 506404 401654 506424
rect 401598 506368 401654 506404
rect 401230 505008 401286 505064
rect 401598 503240 401654 503296
rect 401598 500248 401654 500304
rect 402058 544720 402114 544776
rect 402058 540912 402114 540968
rect 402058 528536 402114 528592
rect 401966 521600 402022 521656
rect 401966 513440 402022 513496
rect 401874 508272 401930 508328
rect 401782 504600 401838 504656
rect 402242 558184 402298 558240
rect 402242 547712 402298 547768
rect 402426 547440 402482 547496
rect 402334 540640 402390 540696
rect 402886 546352 402942 546408
rect 402886 546080 402942 546136
rect 402518 534656 402574 534712
rect 402334 514800 402390 514856
rect 402150 510448 402206 510504
rect 402058 508408 402114 508464
rect 402426 512760 402482 512816
rect 402886 510720 402942 510776
rect 402886 509360 402942 509416
rect 405002 559680 405058 559736
rect 444378 44784 444434 44840
rect 477682 636112 477738 636168
rect 478142 617752 478198 617808
rect 477590 534248 477646 534304
rect 477590 532772 477646 532808
rect 477590 532752 477592 532772
rect 477592 532752 477644 532772
rect 477644 532752 477646 532772
rect 477590 531392 477646 531448
rect 477590 528944 477646 529000
rect 477590 527196 477646 527232
rect 477590 527176 477592 527196
rect 477592 527176 477644 527196
rect 477644 527176 477646 527196
rect 477682 526768 477738 526824
rect 477590 525836 477646 525872
rect 477590 525816 477592 525836
rect 477592 525816 477644 525836
rect 477644 525816 477646 525836
rect 478142 524864 478198 524920
rect 477866 520240 477922 520296
rect 477590 519288 477646 519344
rect 477590 517928 477646 517984
rect 477682 517656 477738 517712
rect 477590 517248 477646 517304
rect 477682 515208 477738 515264
rect 477590 514936 477646 514992
rect 477590 513848 477646 513904
rect 477682 512488 477738 512544
rect 477590 511808 477646 511864
rect 477590 509360 477646 509416
rect 477498 506640 477554 506696
rect 477498 502832 477554 502888
rect 477590 501608 477646 501664
rect 477498 501200 477554 501256
rect 477498 500112 477554 500168
rect 477590 498752 477646 498808
rect 478142 512100 478198 512136
rect 478142 512080 478144 512100
rect 478144 512080 478196 512100
rect 478196 512080 478198 512100
rect 478142 510484 478144 510504
rect 478144 510484 478196 510504
rect 478196 510484 478198 510504
rect 478142 510448 478198 510484
rect 478142 508408 478198 508464
rect 478142 503784 478198 503840
rect 478602 536152 478658 536208
rect 478418 535336 478474 535392
rect 479062 537648 479118 537704
rect 478786 534112 478842 534168
rect 478694 530576 478750 530632
rect 478602 528536 478658 528592
rect 478418 523368 478474 523424
rect 478326 506368 478382 506424
rect 478510 520648 478566 520704
rect 478970 523096 479026 523152
rect 478786 521872 478842 521928
rect 479338 536968 479394 537024
rect 479246 507048 479302 507104
rect 479154 504328 479210 504384
rect 502338 660184 502394 660240
rect 507858 660184 507914 660240
rect 490746 543632 490802 543688
rect 498382 541048 498438 541104
rect 508318 543496 508374 543552
rect 506754 539824 506810 539880
rect 486146 539688 486202 539744
rect 495806 539688 495862 539744
rect 502154 539688 502210 539744
rect 505558 539688 505614 539744
rect 513838 541048 513894 541104
rect 517058 539824 517114 539880
rect 516414 539688 516470 539744
rect 519634 539008 519690 539064
rect 519450 531120 519506 531176
rect 484490 496848 484546 496904
rect 485778 281444 485834 281480
rect 485778 281424 485780 281444
rect 485780 281424 485832 281444
rect 485832 281424 485834 281444
rect 496082 499568 496138 499624
rect 494702 496848 494758 496904
rect 496082 496848 496138 496904
rect 495898 3304 495954 3360
rect 502568 499840 502624 499896
rect 502982 3440 503038 3496
rect 510066 3984 510122 4040
rect 513562 3440 513618 3496
rect 519542 530032 519598 530088
rect 519726 528944 519782 529000
rect 520094 518404 520150 518460
rect 519910 505144 519966 505200
rect 519726 500520 519782 500576
rect 520002 503784 520058 503840
rect 520370 526564 520426 526620
rect 520646 527312 520702 527368
rect 520554 520104 520610 520160
rect 520554 517520 520610 517576
rect 520462 515480 520518 515536
rect 520370 508884 520426 508940
rect 520830 612312 520886 612368
rect 520738 508680 520794 508736
rect 520738 505688 520794 505744
rect 521014 528536 521070 528592
rect 520922 515616 520978 515672
rect 521106 520240 521162 520296
rect 521750 630672 521806 630728
rect 521750 535472 521806 535528
rect 521658 510176 521714 510232
rect 521934 641688 521990 641744
rect 521934 612312 521990 612368
rect 521934 524592 521990 524648
rect 521842 512760 521898 512816
rect 521842 500928 521898 500984
rect 522026 517384 522082 517440
rect 522026 513712 522082 513768
rect 522302 536968 522358 537024
rect 522210 536288 522266 536344
rect 522210 534248 522266 534304
rect 522118 500792 522174 500848
rect 522946 532344 523002 532400
rect 522946 525836 523002 525872
rect 522946 525816 522948 525836
rect 522948 525816 523000 525836
rect 523000 525816 523002 525836
rect 522946 523096 523002 523152
rect 522486 521872 522542 521928
rect 522394 502424 522450 502480
rect 522946 520920 523002 520976
rect 522854 513204 522856 513224
rect 522856 513204 522908 513224
rect 522908 513204 522910 513224
rect 522854 513168 522910 513204
rect 522946 511128 523002 511184
rect 522578 510584 522634 510640
rect 522946 506524 523002 506560
rect 522946 506504 522948 506524
rect 522948 506504 523000 506524
rect 523000 506504 523002 506524
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 580262 564304 580318 564360
rect 580262 553968 580318 554024
rect 580170 537784 580226 537840
rect 579802 524456 579858 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 471416 580226 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 579802 431568 579858 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580262 86128 580318 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect 300117 700362 300183 700365
rect 360694 700362 360700 700364
rect 300117 700360 360700 700362
rect 300117 700304 300122 700360
rect 300178 700304 360700 700360
rect 300117 700302 360700 700304
rect 300117 700299 300183 700302
rect 360694 700300 360700 700302
rect 360764 700300 360770 700364
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3233 671258 3299 671261
rect -960 671256 3299 671258
rect -960 671200 3238 671256
rect 3294 671200 3299 671256
rect -960 671198 3299 671200
rect -960 671108 480 671198
rect 3233 671195 3299 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect 47945 663234 48011 663237
rect 283414 663234 283420 663236
rect 47945 663232 283420 663234
rect 47945 663176 47950 663232
rect 48006 663176 283420 663232
rect 47945 663174 283420 663176
rect 47945 663171 48011 663174
rect 283414 663172 283420 663174
rect 283484 663172 283490 663236
rect 71773 663098 71839 663101
rect 405038 663098 405044 663100
rect 71773 663096 405044 663098
rect 71773 663040 71778 663096
rect 71834 663040 405044 663096
rect 71773 663038 405044 663040
rect 71773 663035 71839 663038
rect 405038 663036 405044 663038
rect 405108 663036 405114 663100
rect 46841 662962 46907 662965
rect 286174 662962 286180 662964
rect 46841 662960 286180 662962
rect 46841 662904 46846 662960
rect 46902 662904 286180 662960
rect 46841 662902 286180 662904
rect 46841 662899 46907 662902
rect 286174 662900 286180 662902
rect 286244 662900 286250 662964
rect 46749 662826 46815 662829
rect 317638 662826 317644 662828
rect 46749 662824 317644 662826
rect 46749 662768 46754 662824
rect 46810 662768 317644 662824
rect 46749 662766 317644 662768
rect 46749 662763 46815 662766
rect 317638 662764 317644 662766
rect 317708 662764 317714 662828
rect 51022 662628 51028 662692
rect 51092 662690 51098 662692
rect 401542 662690 401548 662692
rect 51092 662630 401548 662690
rect 51092 662628 51098 662630
rect 401542 662628 401548 662630
rect 401612 662628 401618 662692
rect 51574 662492 51580 662556
rect 51644 662554 51650 662556
rect 403014 662554 403020 662556
rect 51644 662494 403020 662554
rect 51644 662492 51650 662494
rect 403014 662492 403020 662494
rect 403084 662492 403090 662556
rect 49969 661874 50035 661877
rect 282310 661874 282316 661876
rect 49969 661872 282316 661874
rect 49969 661816 49974 661872
rect 50030 661816 282316 661872
rect 49969 661814 282316 661816
rect 49969 661811 50035 661814
rect 282310 661812 282316 661814
rect 282380 661812 282386 661876
rect 50153 661738 50219 661741
rect 295006 661738 295012 661740
rect 50153 661736 295012 661738
rect 50153 661680 50158 661736
rect 50214 661680 295012 661736
rect 50153 661678 295012 661680
rect 50153 661675 50219 661678
rect 295006 661676 295012 661678
rect 295076 661676 295082 661740
rect 49325 661602 49391 661605
rect 295926 661602 295932 661604
rect 49325 661600 295932 661602
rect 49325 661544 49330 661600
rect 49386 661544 295932 661600
rect 49325 661542 295932 661544
rect 49325 661539 49391 661542
rect 295926 661540 295932 661542
rect 295996 661540 296002 661604
rect 50061 661466 50127 661469
rect 297214 661466 297220 661468
rect 50061 661464 297220 661466
rect 50061 661408 50066 661464
rect 50122 661408 297220 661464
rect 50061 661406 297220 661408
rect 50061 661403 50127 661406
rect 297214 661404 297220 661406
rect 297284 661404 297290 661468
rect 310513 661466 310579 661469
rect 311014 661466 311020 661468
rect 310513 661464 311020 661466
rect 310513 661408 310518 661464
rect 310574 661408 311020 661464
rect 310513 661406 311020 661408
rect 310513 661403 310579 661406
rect 311014 661404 311020 661406
rect 311084 661404 311090 661468
rect 49049 661330 49115 661333
rect 308622 661330 308628 661332
rect 49049 661328 308628 661330
rect 49049 661272 49054 661328
rect 49110 661272 308628 661328
rect 49049 661270 308628 661272
rect 49049 661267 49115 661270
rect 308622 661268 308628 661270
rect 308692 661268 308698 661332
rect 358813 661330 358879 661333
rect 359958 661330 359964 661332
rect 358813 661328 359964 661330
rect 358813 661272 358818 661328
rect 358874 661272 359964 661328
rect 358813 661270 359964 661272
rect 358813 661267 358879 661270
rect 359958 661268 359964 661270
rect 360028 661268 360034 661332
rect 401593 661330 401659 661333
rect 401726 661330 401732 661332
rect 401593 661328 401732 661330
rect 401593 661272 401598 661328
rect 401654 661272 401732 661328
rect 401593 661270 401732 661272
rect 401593 661267 401659 661270
rect 401726 661268 401732 661270
rect 401796 661268 401802 661332
rect 48998 661132 49004 661196
rect 49068 661194 49074 661196
rect 309358 661194 309364 661196
rect 49068 661134 309364 661194
rect 49068 661132 49074 661134
rect 309358 661132 309364 661134
rect 309428 661132 309434 661196
rect 48957 661058 49023 661061
rect 309174 661058 309180 661060
rect 48957 661056 309180 661058
rect 48957 661000 48962 661056
rect 49018 661000 309180 661056
rect 48957 660998 309180 661000
rect 48957 660995 49023 660998
rect 309174 660996 309180 660998
rect 309244 660996 309250 661060
rect 51441 660650 51507 660653
rect 279366 660650 279372 660652
rect 51441 660648 279372 660650
rect 51441 660592 51446 660648
rect 51502 660592 279372 660648
rect 51441 660590 279372 660592
rect 51441 660587 51507 660590
rect 279366 660588 279372 660590
rect 279436 660588 279442 660652
rect 49366 660452 49372 660516
rect 49436 660514 49442 660516
rect 279969 660514 280035 660517
rect 49436 660512 280035 660514
rect 49436 660456 279974 660512
rect 280030 660456 280035 660512
rect 49436 660454 280035 660456
rect 49436 660452 49442 660454
rect 279969 660451 280035 660454
rect 49233 660378 49299 660381
rect 308806 660378 308812 660380
rect 49233 660376 308812 660378
rect 49233 660320 49238 660376
rect 49294 660320 308812 660376
rect 49233 660318 308812 660320
rect 49233 660315 49299 660318
rect 308806 660316 308812 660318
rect 308876 660316 308882 660380
rect 49182 660180 49188 660244
rect 49252 660242 49258 660244
rect 310462 660242 310468 660244
rect 49252 660182 310468 660242
rect 49252 660180 49258 660182
rect 310462 660180 310468 660182
rect 310532 660180 310538 660244
rect 502333 660242 502399 660245
rect 502926 660242 502932 660244
rect 502333 660240 502932 660242
rect 502333 660184 502338 660240
rect 502394 660184 502932 660240
rect 502333 660182 502932 660184
rect 502333 660179 502399 660182
rect 502926 660180 502932 660182
rect 502996 660180 503002 660244
rect 507853 660242 507919 660245
rect 508446 660242 508452 660244
rect 507853 660240 508452 660242
rect 507853 660184 507858 660240
rect 507914 660184 508452 660240
rect 507853 660182 508452 660184
rect 507853 660179 507919 660182
rect 508446 660180 508452 660182
rect 508516 660180 508522 660244
rect 48589 660106 48655 660109
rect 311934 660106 311940 660108
rect 48589 660104 311940 660106
rect 48589 660048 48594 660104
rect 48650 660048 311940 660104
rect 48589 660046 311940 660048
rect 48589 660043 48655 660046
rect 311934 660044 311940 660046
rect 312004 660044 312010 660108
rect 3601 659970 3667 659973
rect 489678 659970 489684 659972
rect 3601 659968 489684 659970
rect 3601 659912 3606 659968
rect 3662 659912 489684 659968
rect 3601 659910 489684 659912
rect 3601 659907 3667 659910
rect 489678 659908 489684 659910
rect 489748 659908 489754 659972
rect 49918 659772 49924 659836
rect 49988 659834 49994 659836
rect 50429 659834 50495 659837
rect 49988 659832 50495 659834
rect 49988 659776 50434 659832
rect 50490 659776 50495 659832
rect 49988 659774 50495 659776
rect 49988 659772 49994 659774
rect 50429 659771 50495 659774
rect 49734 659636 49740 659700
rect 49804 659698 49810 659700
rect 49877 659698 49943 659701
rect 49804 659696 49943 659698
rect 49804 659640 49882 659696
rect 49938 659640 49943 659696
rect 49804 659638 49943 659640
rect 49804 659636 49810 659638
rect 49877 659635 49943 659638
rect 50102 659636 50108 659700
rect 50172 659698 50178 659700
rect 50245 659698 50311 659701
rect 50172 659696 50311 659698
rect 50172 659640 50250 659696
rect 50306 659640 50311 659696
rect 50172 659638 50311 659640
rect 50172 659636 50178 659638
rect 50245 659635 50311 659638
rect -960 658202 480 658292
rect 3325 658202 3391 658205
rect 254761 658202 254827 658205
rect -960 658200 3391 658202
rect -960 658144 3330 658200
rect 3386 658144 3391 658200
rect -960 658142 3391 658144
rect 251804 658200 254827 658202
rect 251804 658144 254766 658200
rect 254822 658144 254827 658200
rect 251804 658142 254827 658144
rect -960 658052 480 658142
rect 3325 658139 3391 658142
rect 254761 658139 254827 658142
rect 583520 657236 584960 657476
rect 49601 655210 49667 655213
rect 49601 655208 52164 655210
rect 49601 655152 49606 655208
rect 49662 655152 52164 655208
rect 49601 655150 52164 655152
rect 49601 655147 49667 655150
rect 254577 652354 254643 652357
rect 251804 652352 254643 652354
rect 251804 652296 254582 652352
rect 254638 652296 254643 652352
rect 251804 652294 254643 652296
rect 254577 652291 254643 652294
rect 49417 649362 49483 649365
rect 49417 649360 52164 649362
rect 49417 649304 49422 649360
rect 49478 649304 52164 649360
rect 49417 649302 52164 649304
rect 49417 649299 49483 649302
rect 254301 646506 254367 646509
rect 251804 646504 254367 646506
rect 251804 646448 254306 646504
rect 254362 646448 254367 646504
rect 251804 646446 254367 646448
rect 254301 646443 254367 646446
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 49509 643514 49575 643517
rect 49509 643512 52164 643514
rect 49509 643456 49514 643512
rect 49570 643456 52164 643512
rect 49509 643454 52164 643456
rect 49509 643451 49575 643454
rect 310053 642290 310119 642293
rect 398189 642290 398255 642293
rect 310053 642288 398255 642290
rect 310053 642232 310058 642288
rect 310114 642232 398194 642288
rect 398250 642232 398255 642288
rect 310053 642230 398255 642232
rect 310053 642227 310119 642230
rect 398189 642227 398255 642230
rect 368933 642154 368999 642157
rect 398598 642154 398604 642156
rect 368933 642152 398604 642154
rect 368933 642096 368938 642152
rect 368994 642096 398604 642152
rect 368933 642094 398604 642096
rect 368933 642091 368999 642094
rect 398598 642092 398604 642094
rect 398668 642092 398674 642156
rect 358854 641956 358860 642020
rect 358924 642018 358930 642020
rect 397085 642018 397151 642021
rect 358924 642016 397151 642018
rect 358924 641960 397090 642016
rect 397146 641960 397151 642016
rect 358924 641958 397151 641960
rect 358924 641956 358930 641958
rect 397085 641955 397151 641958
rect 331949 641882 332015 641885
rect 382181 641882 382247 641885
rect 331949 641880 382247 641882
rect 331949 641824 331954 641880
rect 332010 641824 382186 641880
rect 382242 641824 382247 641880
rect 331949 641822 382247 641824
rect 331949 641819 332015 641822
rect 382181 641819 382247 641822
rect 363454 641684 363460 641748
rect 363524 641746 363530 641748
rect 369485 641746 369551 641749
rect 363524 641744 369551 641746
rect 363524 641688 369490 641744
rect 369546 641688 369551 641744
rect 363524 641686 369551 641688
rect 363524 641684 363530 641686
rect 369485 641683 369551 641686
rect 398189 641746 398255 641749
rect 399201 641746 399267 641749
rect 521929 641746 521995 641749
rect 398189 641744 521995 641746
rect 398189 641688 398194 641744
rect 398250 641688 399206 641744
rect 399262 641688 521934 641744
rect 521990 641688 521995 641744
rect 398189 641686 521995 641688
rect 398189 641683 398255 641686
rect 399201 641683 399267 641686
rect 521929 641683 521995 641686
rect 304758 641004 304764 641068
rect 304828 641066 304834 641068
rect 378041 641066 378107 641069
rect 304828 641064 378107 641066
rect 304828 641008 378046 641064
rect 378102 641008 378107 641064
rect 304828 641006 378107 641008
rect 304828 641004 304834 641006
rect 378041 641003 378107 641006
rect 306230 640868 306236 640932
rect 306300 640930 306306 640932
rect 379513 640930 379579 640933
rect 306300 640928 379579 640930
rect 306300 640872 379518 640928
rect 379574 640872 379579 640928
rect 306300 640870 379579 640872
rect 306300 640868 306306 640870
rect 379513 640867 379579 640870
rect 254301 640658 254367 640661
rect 251804 640656 254367 640658
rect 251804 640600 254306 640656
rect 254362 640600 254367 640656
rect 251804 640598 254367 640600
rect 254301 640595 254367 640598
rect 307477 640658 307543 640661
rect 351126 640658 351132 640660
rect 307477 640656 351132 640658
rect 307477 640600 307482 640656
rect 307538 640600 351132 640656
rect 307477 640598 351132 640600
rect 307477 640595 307543 640598
rect 351126 640596 351132 640598
rect 351196 640596 351202 640660
rect 304165 640522 304231 640525
rect 355174 640522 355180 640524
rect 304165 640520 355180 640522
rect 304165 640464 304170 640520
rect 304226 640464 355180 640520
rect 304165 640462 355180 640464
rect 304165 640459 304231 640462
rect 355174 640460 355180 640462
rect 355244 640460 355250 640524
rect 301446 640324 301452 640388
rect 301516 640386 301522 640388
rect 378869 640386 378935 640389
rect 301516 640384 378935 640386
rect 301516 640328 378874 640384
rect 378930 640328 378935 640384
rect 301516 640326 378935 640328
rect 301516 640324 301522 640326
rect 378869 640323 378935 640326
rect 373950 639782 383670 639842
rect 358670 639644 358676 639708
rect 358740 639706 358746 639708
rect 358740 639646 369870 639706
rect 358740 639644 358746 639646
rect 362493 639570 362559 639573
rect 362718 639570 362724 639572
rect 362493 639568 362724 639570
rect 362493 639512 362498 639568
rect 362554 639512 362724 639568
rect 362493 639510 362724 639512
rect 362493 639507 362559 639510
rect 362718 639508 362724 639510
rect 362788 639508 362794 639572
rect 308581 639434 308647 639437
rect 355358 639434 355364 639436
rect 308581 639432 355364 639434
rect 308581 639376 308586 639432
rect 308642 639376 355364 639432
rect 308581 639374 355364 639376
rect 308581 639371 308647 639374
rect 355358 639372 355364 639374
rect 355428 639372 355434 639436
rect 361941 639434 362007 639437
rect 362585 639436 362651 639437
rect 364057 639436 364123 639437
rect 362350 639434 362356 639436
rect 361941 639432 362356 639434
rect 361941 639376 361946 639432
rect 362002 639376 362356 639432
rect 361941 639374 362356 639376
rect 361941 639371 362007 639374
rect 362350 639372 362356 639374
rect 362420 639372 362426 639436
rect 362534 639434 362540 639436
rect 362494 639374 362540 639434
rect 362604 639432 362651 639436
rect 364006 639434 364012 639436
rect 362646 639376 362651 639432
rect 362534 639372 362540 639374
rect 362604 639372 362651 639376
rect 363966 639374 364012 639434
rect 364076 639432 364123 639436
rect 364118 639376 364123 639432
rect 364006 639372 364012 639374
rect 364076 639372 364123 639376
rect 362585 639371 362651 639372
rect 364057 639371 364123 639372
rect 368105 639434 368171 639437
rect 369669 639434 369735 639437
rect 368105 639432 369735 639434
rect 368105 639376 368110 639432
rect 368166 639376 369674 639432
rect 369730 639376 369735 639432
rect 368105 639374 369735 639376
rect 369810 639434 369870 639646
rect 373950 639434 374010 639782
rect 377254 639644 377260 639708
rect 377324 639706 377330 639708
rect 380157 639706 380223 639709
rect 377324 639704 380223 639706
rect 377324 639648 380162 639704
rect 380218 639648 380223 639704
rect 377324 639646 380223 639648
rect 377324 639644 377330 639646
rect 380157 639643 380223 639646
rect 381118 639508 381124 639572
rect 381188 639570 381194 639572
rect 382917 639570 382983 639573
rect 381188 639568 382983 639570
rect 381188 639512 382922 639568
rect 382978 639512 382983 639568
rect 381188 639510 382983 639512
rect 381188 639508 381194 639510
rect 382917 639507 382983 639510
rect 380893 639434 380959 639437
rect 369810 639374 374010 639434
rect 377630 639432 380959 639434
rect 377630 639376 380898 639432
rect 380954 639376 380959 639432
rect 377630 639374 380959 639376
rect 383610 639434 383670 639782
rect 391289 639434 391355 639437
rect 383610 639432 391355 639434
rect 383610 639376 391294 639432
rect 391350 639376 391355 639432
rect 383610 639374 391355 639376
rect 368105 639371 368171 639374
rect 369669 639371 369735 639374
rect 285397 639300 285463 639301
rect 288249 639300 288315 639301
rect 285397 639296 285444 639300
rect 285508 639298 285514 639300
rect 288198 639298 288204 639300
rect 285397 639240 285402 639296
rect 285397 639236 285444 639240
rect 285508 639238 285554 639298
rect 288158 639238 288204 639298
rect 288268 639296 288315 639300
rect 288310 639240 288315 639296
rect 285508 639236 285514 639238
rect 288198 639236 288204 639238
rect 288268 639236 288315 639240
rect 289486 639236 289492 639300
rect 289556 639298 289562 639300
rect 289629 639298 289695 639301
rect 289556 639296 289695 639298
rect 289556 639240 289634 639296
rect 289690 639240 289695 639296
rect 289556 639238 289695 639240
rect 289556 639236 289562 639238
rect 285397 639235 285463 639236
rect 288249 639235 288315 639236
rect 289629 639235 289695 639238
rect 290917 639300 290983 639301
rect 290917 639296 290964 639300
rect 291028 639298 291034 639300
rect 292021 639298 292087 639301
rect 292430 639298 292436 639300
rect 290917 639240 290922 639296
rect 290917 639236 290964 639240
rect 291028 639238 291074 639298
rect 292021 639296 292436 639298
rect 292021 639240 292026 639296
rect 292082 639240 292436 639296
rect 292021 639238 292436 639240
rect 291028 639236 291034 639238
rect 290917 639235 290983 639236
rect 292021 639235 292087 639238
rect 292430 639236 292436 639238
rect 292500 639236 292506 639300
rect 293125 639298 293191 639301
rect 298461 639300 298527 639301
rect 293718 639298 293724 639300
rect 293125 639296 293724 639298
rect 293125 639240 293130 639296
rect 293186 639240 293724 639296
rect 293125 639238 293724 639240
rect 293125 639235 293191 639238
rect 293718 639236 293724 639238
rect 293788 639236 293794 639300
rect 298461 639296 298508 639300
rect 298572 639298 298578 639300
rect 298461 639240 298466 639296
rect 298461 639236 298508 639240
rect 298572 639238 298618 639298
rect 298572 639236 298578 639238
rect 306966 639236 306972 639300
rect 307036 639298 307042 639300
rect 377630 639298 377690 639374
rect 380893 639371 380959 639374
rect 391289 639371 391355 639374
rect 307036 639238 377690 639298
rect 307036 639236 307042 639238
rect 298461 639235 298527 639236
rect 300710 639100 300716 639164
rect 300780 639162 300786 639164
rect 377254 639162 377260 639164
rect 300780 639102 377260 639162
rect 300780 639100 300786 639102
rect 377254 639100 377260 639102
rect 377324 639100 377330 639164
rect 303470 638964 303476 639028
rect 303540 639026 303546 639028
rect 381118 639026 381124 639028
rect 303540 638966 381124 639026
rect 303540 638964 303546 638966
rect 381118 638964 381124 638966
rect 381188 638964 381194 639028
rect 49366 637604 49372 637668
rect 49436 637666 49442 637668
rect 49436 637606 52164 637666
rect 49436 637604 49442 637606
rect 49366 637468 49372 637532
rect 49436 637530 49442 637532
rect 50521 637530 50587 637533
rect 49436 637528 50587 637530
rect 49436 637472 50526 637528
rect 50582 637472 50587 637528
rect 49436 637470 50587 637472
rect 49436 637468 49442 637470
rect 50521 637467 50587 637470
rect 477677 636170 477743 636173
rect 477677 636168 480148 636170
rect 477677 636112 477682 636168
rect 477738 636112 480148 636168
rect 477677 636110 480148 636112
rect 477677 636107 477743 636110
rect 254669 634810 254735 634813
rect 251804 634808 254735 634810
rect 251804 634752 254674 634808
rect 254730 634752 254735 634808
rect 251804 634750 254735 634752
rect 254669 634747 254735 634750
rect -960 631940 480 632180
rect 48865 631818 48931 631821
rect 48865 631816 52164 631818
rect 48865 631760 48870 631816
rect 48926 631760 52164 631816
rect 48865 631758 52164 631760
rect 48865 631755 48931 631758
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 521745 630730 521811 630733
rect 519892 630728 521811 630730
rect 519892 630672 521750 630728
rect 521806 630672 521811 630728
rect 583520 630716 584960 630806
rect 519892 630670 521811 630672
rect 521745 630667 521811 630670
rect 278773 630050 278839 630053
rect 278773 630048 280140 630050
rect 278773 629992 278778 630048
rect 278834 629992 280140 630048
rect 278773 629990 280140 629992
rect 278773 629987 278839 629990
rect 254669 628962 254735 628965
rect 251804 628960 254735 628962
rect 251804 628904 254674 628960
rect 254730 628904 254735 628960
rect 251804 628902 254735 628904
rect 254669 628899 254735 628902
rect 50705 625970 50771 625973
rect 50705 625968 52164 625970
rect 50705 625912 50710 625968
rect 50766 625912 52164 625968
rect 50705 625910 52164 625912
rect 50705 625907 50771 625910
rect 254669 623114 254735 623117
rect 251804 623112 254735 623114
rect 251804 623056 254674 623112
rect 254730 623056 254735 623112
rect 251804 623054 254735 623056
rect 254669 623051 254735 623054
rect 48589 620122 48655 620125
rect 48589 620120 52164 620122
rect 48589 620064 48594 620120
rect 48650 620064 52164 620120
rect 48589 620062 52164 620064
rect 48589 620059 48655 620062
rect -960 619170 480 619260
rect -960 619110 674 619170
rect -960 619034 480 619110
rect 614 619034 674 619110
rect -960 619020 674 619034
rect 246 618974 674 619020
rect 246 618490 306 618974
rect 246 618430 6930 618490
rect 6870 618354 6930 618430
rect 50102 618354 50108 618356
rect 6870 618294 50108 618354
rect 50102 618292 50108 618294
rect 50172 618292 50178 618356
rect 478137 617810 478203 617813
rect 478137 617808 480148 617810
rect 478137 617752 478142 617808
rect 478198 617752 480148 617808
rect 478137 617750 480148 617752
rect 478137 617747 478203 617750
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect 254393 617266 254459 617269
rect 251804 617264 254459 617266
rect 251804 617208 254398 617264
rect 254454 617208 254459 617264
rect 251804 617206 254459 617208
rect 254393 617203 254459 617206
rect 49182 614212 49188 614276
rect 49252 614274 49258 614276
rect 49252 614214 52164 614274
rect 49252 614212 49258 614214
rect 48497 612778 48563 612781
rect 49550 612778 49556 612780
rect 48497 612776 49556 612778
rect 48497 612720 48502 612776
rect 48558 612720 49556 612776
rect 48497 612718 49556 612720
rect 48497 612715 48563 612718
rect 49550 612716 49556 612718
rect 49620 612716 49626 612780
rect 520825 612370 520891 612373
rect 521929 612370 521995 612373
rect 519892 612368 521995 612370
rect 519892 612312 520830 612368
rect 520886 612312 521934 612368
rect 521990 612312 521995 612368
rect 519892 612310 521995 612312
rect 520825 612307 520891 612310
rect 521929 612307 521995 612310
rect 254485 611418 254551 611421
rect 251804 611416 254551 611418
rect 251804 611360 254490 611416
rect 254546 611360 254551 611416
rect 251804 611358 254551 611360
rect 254485 611355 254551 611358
rect 278681 610058 278747 610061
rect 278681 610056 280140 610058
rect 278681 610000 278686 610056
rect 278742 610000 280140 610056
rect 278681 609998 280140 610000
rect 278681 609995 278747 609998
rect 49550 608364 49556 608428
rect 49620 608426 49626 608428
rect 49620 608366 52164 608426
rect 49620 608364 49626 608366
rect 49550 607140 49556 607204
rect 49620 607202 49626 607204
rect 51809 607202 51875 607205
rect 49620 607200 51875 607202
rect 49620 607144 51814 607200
rect 51870 607144 51875 607200
rect 49620 607142 51875 607144
rect 49620 607140 49626 607142
rect 51809 607139 51875 607142
rect -960 606114 480 606204
rect -960 606054 6930 606114
rect -960 605964 480 606054
rect 6870 605978 6930 606054
rect 49918 605978 49924 605980
rect 6870 605918 49924 605978
rect 49918 605916 49924 605918
rect 49988 605916 49994 605980
rect 254209 605570 254275 605573
rect 251804 605568 254275 605570
rect 251804 605512 254214 605568
rect 254270 605512 254275 605568
rect 251804 605510 254275 605512
rect 254209 605507 254275 605510
rect 583520 604060 584960 604300
rect 48998 602516 49004 602580
rect 49068 602578 49074 602580
rect 49068 602518 52164 602578
rect 49068 602516 49074 602518
rect 49182 601020 49188 601084
rect 49252 601082 49258 601084
rect 51574 601082 51580 601084
rect 49252 601022 51580 601082
rect 49252 601020 49258 601022
rect 51574 601020 51580 601022
rect 51644 601020 51650 601084
rect 303429 600676 303495 600677
rect 304717 600676 304783 600677
rect 306189 600676 306255 600677
rect 303429 600674 303476 600676
rect 303384 600672 303476 600674
rect 303384 600616 303434 600672
rect 303384 600614 303476 600616
rect 303429 600612 303476 600614
rect 303540 600612 303546 600676
rect 304717 600674 304764 600676
rect 304672 600672 304764 600674
rect 304672 600616 304722 600672
rect 304672 600614 304764 600616
rect 304717 600612 304764 600614
rect 304828 600612 304834 600676
rect 306189 600674 306236 600676
rect 306144 600672 306236 600674
rect 306144 600616 306194 600672
rect 306144 600614 306236 600616
rect 306189 600612 306236 600614
rect 306300 600612 306306 600676
rect 303429 600611 303495 600612
rect 304717 600611 304783 600612
rect 306189 600611 306255 600612
rect 301405 600538 301471 600541
rect 306966 600538 306972 600540
rect 301405 600536 306972 600538
rect 301405 600480 301410 600536
rect 301466 600480 306972 600536
rect 301405 600478 306972 600480
rect 301405 600475 301471 600478
rect 306966 600476 306972 600478
rect 307036 600476 307042 600540
rect 300669 600132 300735 600133
rect 300669 600128 300716 600132
rect 300780 600130 300786 600132
rect 300669 600072 300674 600128
rect 300669 600068 300716 600072
rect 300780 600070 300826 600130
rect 300780 600068 300786 600070
rect 300669 600067 300735 600068
rect 254853 599722 254919 599725
rect 251804 599720 254919 599722
rect 251804 599664 254858 599720
rect 254914 599664 254919 599720
rect 251804 599662 254919 599664
rect 254853 599659 254919 599662
rect 360009 599586 360075 599589
rect 369894 599586 369900 599588
rect 360009 599584 369900 599586
rect 360009 599528 360014 599584
rect 360070 599528 369900 599584
rect 360009 599526 369900 599528
rect 360009 599523 360075 599526
rect 369894 599524 369900 599526
rect 369964 599524 369970 599588
rect 299289 598906 299355 598909
rect 301446 598906 301452 598908
rect 299289 598904 301452 598906
rect 299289 598848 299294 598904
rect 299350 598848 301452 598904
rect 299289 598846 301452 598848
rect 299289 598843 299355 598846
rect 301446 598844 301452 598846
rect 301516 598844 301522 598908
rect 382222 598164 382228 598228
rect 382292 598226 382298 598228
rect 383285 598226 383351 598229
rect 382292 598224 383351 598226
rect 382292 598168 383290 598224
rect 383346 598168 383351 598224
rect 382292 598166 383351 598168
rect 382292 598164 382298 598166
rect 383285 598163 383351 598166
rect 307017 597684 307083 597685
rect 306966 597620 306972 597684
rect 307036 597682 307083 597684
rect 307036 597680 307128 597682
rect 307078 597624 307128 597680
rect 307036 597622 307128 597624
rect 307036 597620 307083 597622
rect 368974 597620 368980 597684
rect 369044 597682 369050 597684
rect 376109 597682 376175 597685
rect 369044 597680 376175 597682
rect 369044 597624 376114 597680
rect 376170 597624 376175 597680
rect 369044 597622 376175 597624
rect 369044 597620 369050 597622
rect 307017 597619 307083 597620
rect 376109 597619 376175 597622
rect 48957 596730 49023 596733
rect 48957 596728 52164 596730
rect 48957 596672 48962 596728
rect 49018 596672 52164 596728
rect 48957 596670 52164 596672
rect 48957 596667 49023 596670
rect 362350 595444 362356 595508
rect 362420 595506 362426 595508
rect 391197 595506 391263 595509
rect 362420 595504 391263 595506
rect 362420 595448 391202 595504
rect 391258 595448 391263 595504
rect 362420 595446 391263 595448
rect 362420 595444 362426 595446
rect 391197 595443 391263 595446
rect 254485 593874 254551 593877
rect 251804 593872 254551 593874
rect 251804 593816 254490 593872
rect 254546 593816 254551 593872
rect 251804 593814 254551 593816
rect 254485 593811 254551 593814
rect 362309 593330 362375 593333
rect 362902 593330 362908 593332
rect 362309 593328 362908 593330
rect 362309 593272 362314 593328
rect 362370 593272 362908 593328
rect 362309 593270 362908 593272
rect 362309 593267 362375 593270
rect 362902 593268 362908 593270
rect 362972 593268 362978 593332
rect 361573 593194 361639 593197
rect 363454 593194 363460 593196
rect 361573 593192 363460 593194
rect -960 592908 480 593148
rect 361573 593136 361578 593192
rect 361634 593136 363460 593192
rect 361573 593134 363460 593136
rect 361573 593131 361639 593134
rect 363454 593132 363460 593134
rect 363524 593132 363530 593196
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 49049 590882 49115 590885
rect 49049 590880 52164 590882
rect 49049 590824 49054 590880
rect 49110 590824 52164 590880
rect 583520 590868 584960 590958
rect 49049 590822 52164 590824
rect 49049 590819 49115 590822
rect 299381 589930 299447 589933
rect 380934 589930 380940 589932
rect 299381 589928 380940 589930
rect 299381 589872 299386 589928
rect 299442 589872 380940 589928
rect 299381 589870 380940 589872
rect 299381 589867 299447 589870
rect 380934 589868 380940 589870
rect 381004 589868 381010 589932
rect 254577 588026 254643 588029
rect 251804 588024 254643 588026
rect 251804 587968 254582 588024
rect 254638 587968 254643 588024
rect 251804 587966 254643 587968
rect 254577 587963 254643 587966
rect 292665 587210 292731 587213
rect 376150 587210 376156 587212
rect 292665 587208 376156 587210
rect 292665 587152 292670 587208
rect 292726 587152 376156 587208
rect 292665 587150 376156 587152
rect 292665 587147 292731 587150
rect 376150 587148 376156 587150
rect 376220 587148 376226 587212
rect 49233 585034 49299 585037
rect 49233 585032 52164 585034
rect 49233 584976 49238 585032
rect 49294 584976 52164 585032
rect 49233 584974 52164 584976
rect 49233 584971 49299 584974
rect 300853 582994 300919 582997
rect 384062 582994 384068 582996
rect 300853 582992 384068 582994
rect 300853 582936 300858 582992
rect 300914 582936 384068 582992
rect 300853 582934 384068 582936
rect 300853 582931 300919 582934
rect 384062 582932 384068 582934
rect 384132 582932 384138 582996
rect 253933 582178 253999 582181
rect 251804 582176 253999 582178
rect 251804 582120 253938 582176
rect 253994 582120 253999 582176
rect 251804 582118 253999 582120
rect 253933 582115 253999 582118
rect 364006 581708 364012 581772
rect 364076 581770 364082 581772
rect 397453 581770 397519 581773
rect 364076 581768 397519 581770
rect 364076 581712 397458 581768
rect 397514 581712 397519 581768
rect 364076 581710 397519 581712
rect 364076 581708 364082 581710
rect 397453 581707 397519 581710
rect 292430 581572 292436 581636
rect 292500 581634 292506 581636
rect 364517 581634 364583 581637
rect 292500 581632 364583 581634
rect 292500 581576 364522 581632
rect 364578 581576 364583 581632
rect 292500 581574 364583 581576
rect 292500 581572 292506 581574
rect 364517 581571 364583 581574
rect 373206 581572 373212 581636
rect 373276 581634 373282 581636
rect 386597 581634 386663 581637
rect 373276 581632 386663 581634
rect 373276 581576 386602 581632
rect 386658 581576 386663 581632
rect 373276 581574 386663 581576
rect 373276 581572 373282 581574
rect 386597 581571 386663 581574
rect 300577 580410 300643 580413
rect 394734 580410 394740 580412
rect 300577 580408 394740 580410
rect 300577 580352 300582 580408
rect 300638 580352 394740 580408
rect 300577 580350 394740 580352
rect 300577 580347 300643 580350
rect 394734 580348 394740 580350
rect 394804 580348 394810 580412
rect 287145 580274 287211 580277
rect 389582 580274 389588 580276
rect 287145 580272 389588 580274
rect 287145 580216 287150 580272
rect 287206 580216 389588 580272
rect 287145 580214 389588 580216
rect 287145 580211 287211 580214
rect 389582 580212 389588 580214
rect 389652 580212 389658 580276
rect -960 579852 480 580092
rect 385534 579532 385540 579596
rect 385604 579594 385610 579596
rect 389265 579594 389331 579597
rect 385604 579592 389331 579594
rect 385604 579536 389270 579592
rect 389326 579536 389331 579592
rect 385604 579534 389331 579536
rect 385604 579532 385610 579534
rect 389265 579531 389331 579534
rect 48681 579186 48747 579189
rect 48681 579184 52164 579186
rect 48681 579128 48686 579184
rect 48742 579128 52164 579184
rect 48681 579126 52164 579128
rect 48681 579123 48747 579126
rect 300669 578914 300735 578917
rect 376886 578914 376892 578916
rect 300669 578912 376892 578914
rect 300669 578856 300674 578912
rect 300730 578856 376892 578912
rect 300669 578854 376892 578856
rect 300669 578851 300735 578854
rect 376886 578852 376892 578854
rect 376956 578852 376962 578916
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 379605 577554 379671 577557
rect 391974 577554 391980 577556
rect 379605 577552 391980 577554
rect 379605 577496 379610 577552
rect 379666 577496 391980 577552
rect 379605 577494 391980 577496
rect 379605 577491 379671 577494
rect 391974 577492 391980 577494
rect 392044 577492 392050 577556
rect 583520 577540 584960 577630
rect 254209 576330 254275 576333
rect 251804 576328 254275 576330
rect 251804 576272 254214 576328
rect 254270 576272 254275 576328
rect 251804 576270 254275 576272
rect 254209 576267 254275 576270
rect 393998 575452 394004 575516
rect 394068 575514 394074 575516
rect 394785 575514 394851 575517
rect 394068 575512 394851 575514
rect 394068 575456 394790 575512
rect 394846 575456 394851 575512
rect 394068 575454 394851 575456
rect 394068 575452 394074 575454
rect 394785 575451 394851 575454
rect 49601 573338 49667 573341
rect 281625 573338 281691 573341
rect 391054 573338 391060 573340
rect 49601 573336 52164 573338
rect 49601 573280 49606 573336
rect 49662 573280 52164 573336
rect 49601 573278 52164 573280
rect 281625 573336 391060 573338
rect 281625 573280 281630 573336
rect 281686 573280 391060 573336
rect 281625 573278 391060 573280
rect 49601 573275 49667 573278
rect 281625 573275 281691 573278
rect 391054 573276 391060 573278
rect 391124 573276 391130 573340
rect 361614 571916 361620 571980
rect 361684 571978 361690 571980
rect 378409 571978 378475 571981
rect 361684 571976 378475 571978
rect 361684 571920 378414 571976
rect 378470 571920 378475 571976
rect 361684 571918 378475 571920
rect 361684 571916 361690 571918
rect 378409 571915 378475 571918
rect 253933 570482 253999 570485
rect 251804 570480 253999 570482
rect 251804 570424 253938 570480
rect 253994 570424 253999 570480
rect 251804 570422 253999 570424
rect 253933 570419 253999 570422
rect 377254 569332 377260 569396
rect 377324 569394 377330 569396
rect 388529 569394 388595 569397
rect 377324 569392 388595 569394
rect 377324 569336 388534 569392
rect 388590 569336 388595 569392
rect 377324 569334 388595 569336
rect 377324 569332 377330 569334
rect 388529 569331 388595 569334
rect 290958 569196 290964 569260
rect 291028 569258 291034 569260
rect 380566 569258 380572 569260
rect 291028 569198 380572 569258
rect 291028 569196 291034 569198
rect 380566 569196 380572 569198
rect 380636 569196 380642 569260
rect 366214 568516 366220 568580
rect 366284 568578 366290 568580
rect 367277 568578 367343 568581
rect 366284 568576 367343 568578
rect 366284 568520 367282 568576
rect 367338 568520 367343 568576
rect 366284 568518 367343 568520
rect 366284 568516 366290 568518
rect 367277 568515 367343 568518
rect 49141 567490 49207 567493
rect 49141 567488 52164 567490
rect 49141 567432 49146 567488
rect 49202 567432 52164 567488
rect 49141 567430 52164 567432
rect 49141 567427 49207 567430
rect -960 566946 480 567036
rect 3325 566946 3391 566949
rect -960 566944 3391 566946
rect -960 566888 3330 566944
rect 3386 566888 3391 566944
rect -960 566886 3391 566888
rect -960 566796 480 566886
rect 3325 566883 3391 566886
rect 376937 565858 377003 565861
rect 378726 565858 378732 565860
rect 376937 565856 378732 565858
rect 376937 565800 376942 565856
rect 376998 565800 378732 565856
rect 376937 565798 378732 565800
rect 376937 565795 377003 565798
rect 378726 565796 378732 565798
rect 378796 565796 378802 565860
rect 362534 564980 362540 565044
rect 362604 565042 362610 565044
rect 370129 565042 370195 565045
rect 362604 565040 370195 565042
rect 362604 564984 370134 565040
rect 370190 564984 370195 565040
rect 362604 564982 370195 564984
rect 362604 564980 362610 564982
rect 370129 564979 370195 564982
rect 254577 564634 254643 564637
rect 251804 564632 254643 564634
rect 251804 564576 254582 564632
rect 254638 564576 254643 564632
rect 251804 564574 254643 564576
rect 254577 564571 254643 564574
rect 385718 564436 385724 564500
rect 385788 564498 385794 564500
rect 388437 564498 388503 564501
rect 385788 564496 388503 564498
rect 385788 564440 388442 564496
rect 388498 564440 388503 564496
rect 385788 564438 388503 564440
rect 385788 564436 385794 564438
rect 388437 564435 388503 564438
rect 580257 564362 580323 564365
rect 583520 564362 584960 564452
rect 580257 564360 584960 564362
rect 580257 564304 580262 564360
rect 580318 564304 584960 564360
rect 580257 564302 584960 564304
rect 580257 564299 580323 564302
rect 583520 564212 584960 564302
rect 282913 563682 282979 563685
rect 364742 563682 364748 563684
rect 282913 563680 364748 563682
rect 282913 563624 282918 563680
rect 282974 563624 364748 563680
rect 282913 563622 364748 563624
rect 282913 563619 282979 563622
rect 364742 563620 364748 563622
rect 364812 563620 364818 563684
rect 368238 563620 368244 563684
rect 368308 563682 368314 563684
rect 382365 563682 382431 563685
rect 368308 563680 382431 563682
rect 368308 563624 382370 563680
rect 382426 563624 382431 563680
rect 368308 563622 382431 563624
rect 368308 563620 368314 563622
rect 382365 563619 382431 563622
rect 382774 563620 382780 563684
rect 382844 563682 382850 563684
rect 392025 563682 392091 563685
rect 382844 563680 392091 563682
rect 382844 563624 392030 563680
rect 392086 563624 392091 563680
rect 382844 563622 392091 563624
rect 382844 563620 382850 563622
rect 392025 563619 392091 563622
rect 370037 563138 370103 563141
rect 371550 563138 371556 563140
rect 370037 563136 371556 563138
rect 370037 563080 370042 563136
rect 370098 563080 371556 563136
rect 370037 563078 371556 563080
rect 370037 563075 370103 563078
rect 371550 563076 371556 563078
rect 371620 563076 371626 563140
rect 378317 562458 378383 562461
rect 386454 562458 386460 562460
rect 378317 562456 386460 562458
rect 378317 562400 378322 562456
rect 378378 562400 386460 562456
rect 378317 562398 386460 562400
rect 378317 562395 378383 562398
rect 386454 562396 386460 562398
rect 386524 562396 386530 562460
rect 289486 562260 289492 562324
rect 289556 562322 289562 562324
rect 400622 562322 400628 562324
rect 289556 562262 400628 562322
rect 289556 562260 289562 562262
rect 400622 562260 400628 562262
rect 400692 562260 400698 562324
rect 49417 561642 49483 561645
rect 49417 561640 52164 561642
rect 49417 561584 49422 561640
rect 49478 561584 52164 561640
rect 49417 561582 52164 561584
rect 49417 561579 49483 561582
rect 311893 561234 311959 561237
rect 376334 561234 376340 561236
rect 311893 561232 376340 561234
rect 311893 561176 311898 561232
rect 311954 561176 376340 561232
rect 311893 561174 376340 561176
rect 311893 561171 311959 561174
rect 376334 561172 376340 561174
rect 376404 561172 376410 561236
rect 298502 561036 298508 561100
rect 298572 561098 298578 561100
rect 400438 561098 400444 561100
rect 298572 561038 400444 561098
rect 298572 561036 298578 561038
rect 400438 561036 400444 561038
rect 400508 561036 400514 561100
rect 285438 560900 285444 560964
rect 285508 560962 285514 560964
rect 399150 560962 399156 560964
rect 285508 560902 399156 560962
rect 285508 560900 285514 560902
rect 399150 560900 399156 560902
rect 399220 560900 399226 560964
rect 358302 559676 358308 559740
rect 358372 559738 358378 559740
rect 404997 559738 405063 559741
rect 358372 559736 405063 559738
rect 358372 559680 405002 559736
rect 405058 559680 405063 559736
rect 358372 559678 405063 559680
rect 358372 559676 358378 559678
rect 404997 559675 405063 559678
rect 280153 559602 280219 559605
rect 398782 559602 398788 559604
rect 280153 559600 398788 559602
rect 280153 559544 280158 559600
rect 280214 559544 398788 559600
rect 280153 559542 398788 559544
rect 280153 559539 280219 559542
rect 398782 559540 398788 559542
rect 398852 559540 398858 559604
rect 254577 558786 254643 558789
rect 251804 558784 254643 558786
rect 251804 558728 254582 558784
rect 254638 558728 254643 558784
rect 251804 558726 254643 558728
rect 254577 558723 254643 558726
rect 361430 558316 361436 558380
rect 361500 558378 361506 558380
rect 378225 558378 378291 558381
rect 361500 558376 378291 558378
rect 361500 558320 378230 558376
rect 378286 558320 378291 558376
rect 361500 558318 378291 558320
rect 361500 558316 361506 558318
rect 378225 558315 378291 558318
rect 288198 558180 288204 558244
rect 288268 558242 288274 558244
rect 402237 558242 402303 558245
rect 288268 558240 402303 558242
rect 288268 558184 402242 558240
rect 402298 558184 402303 558240
rect 288268 558182 402303 558184
rect 288268 558180 288274 558182
rect 402237 558179 402303 558182
rect 309317 556746 309383 556749
rect 400254 556746 400260 556748
rect 309317 556744 400260 556746
rect 309317 556688 309322 556744
rect 309378 556688 400260 556744
rect 309317 556686 400260 556688
rect 309317 556683 309383 556686
rect 400254 556684 400260 556686
rect 400324 556684 400330 556748
rect 48773 555794 48839 555797
rect 48773 555792 52164 555794
rect 48773 555736 48778 555792
rect 48834 555736 52164 555792
rect 48773 555734 52164 555736
rect 48773 555731 48839 555734
rect 358118 555460 358124 555524
rect 358188 555522 358194 555524
rect 371233 555522 371299 555525
rect 358188 555520 371299 555522
rect 358188 555464 371238 555520
rect 371294 555464 371299 555520
rect 358188 555462 371299 555464
rect 358188 555460 358194 555462
rect 371233 555459 371299 555462
rect 289813 555386 289879 555389
rect 399334 555386 399340 555388
rect 289813 555384 399340 555386
rect 289813 555328 289818 555384
rect 289874 555328 399340 555384
rect 289813 555326 399340 555328
rect 289813 555323 289879 555326
rect 399334 555324 399340 555326
rect 399404 555324 399410 555388
rect 358486 554100 358492 554164
rect 358556 554162 358562 554164
rect 369853 554162 369919 554165
rect 358556 554160 369919 554162
rect 358556 554104 369858 554160
rect 369914 554104 369919 554160
rect 358556 554102 369919 554104
rect 358556 554100 358562 554102
rect 369853 554099 369919 554102
rect -960 553890 480 553980
rect 359038 553964 359044 554028
rect 359108 554026 359114 554028
rect 580257 554026 580323 554029
rect 359108 554024 580323 554026
rect 359108 553968 580262 554024
rect 580318 553968 580323 554024
rect 359108 553966 580323 553968
rect 359108 553964 359114 553966
rect 580257 553963 580323 553966
rect 2957 553890 3023 553893
rect -960 553888 3023 553890
rect -960 553832 2962 553888
rect 3018 553832 3023 553888
rect -960 553830 3023 553832
rect -960 553740 480 553830
rect 2957 553827 3023 553830
rect 254577 552938 254643 552941
rect 251804 552936 254643 552938
rect 251804 552880 254582 552936
rect 254638 552880 254643 552936
rect 251804 552878 254643 552880
rect 254577 552875 254643 552878
rect 359958 552604 359964 552668
rect 360028 552666 360034 552668
rect 376753 552666 376819 552669
rect 360028 552664 376819 552666
rect 360028 552608 376758 552664
rect 376814 552608 376819 552664
rect 360028 552606 376819 552608
rect 360028 552604 360034 552606
rect 376753 552603 376819 552606
rect 360009 552122 360075 552125
rect 403566 552122 403572 552124
rect 360009 552120 403572 552122
rect 360009 552064 360014 552120
rect 360070 552064 403572 552120
rect 360009 552062 403572 552064
rect 360009 552059 360075 552062
rect 403566 552060 403572 552062
rect 403636 552060 403642 552124
rect 359222 551924 359228 551988
rect 359292 551986 359298 551988
rect 361849 551986 361915 551989
rect 359292 551984 361915 551986
rect 359292 551928 361854 551984
rect 361910 551928 361915 551984
rect 359292 551926 361915 551928
rect 359292 551924 359298 551926
rect 361849 551923 361915 551926
rect 359406 551652 359412 551716
rect 359476 551714 359482 551716
rect 368473 551714 368539 551717
rect 359476 551712 368539 551714
rect 359476 551656 368478 551712
rect 368534 551656 368539 551712
rect 359476 551654 368539 551656
rect 359476 551652 359482 551654
rect 368473 551651 368539 551654
rect 362718 551516 362724 551580
rect 362788 551578 362794 551580
rect 401133 551578 401199 551581
rect 362788 551576 401199 551578
rect 362788 551520 401138 551576
rect 401194 551520 401199 551576
rect 362788 551518 401199 551520
rect 362788 551516 362794 551518
rect 401133 551515 401199 551518
rect 298093 551442 298159 551445
rect 400806 551442 400812 551444
rect 298093 551440 400812 551442
rect 298093 551384 298098 551440
rect 298154 551384 400812 551440
rect 298093 551382 400812 551384
rect 298093 551379 298159 551382
rect 400806 551380 400812 551382
rect 400876 551380 400882 551444
rect 293718 551244 293724 551308
rect 293788 551306 293794 551308
rect 398966 551306 398972 551308
rect 293788 551246 398972 551306
rect 293788 551244 293794 551246
rect 398966 551244 398972 551246
rect 399036 551244 399042 551308
rect 583520 551020 584960 551260
rect 357065 550354 357131 550357
rect 357065 550352 360210 550354
rect 357065 550296 357070 550352
rect 357126 550296 360210 550352
rect 357065 550294 360210 550296
rect 357065 550291 357131 550294
rect 48865 549946 48931 549949
rect 48865 549944 52164 549946
rect 48865 549888 48870 549944
rect 48926 549888 52164 549944
rect 48865 549886 52164 549888
rect 48865 549883 48931 549886
rect 360150 549712 360210 550294
rect 397637 550082 397703 550085
rect 401910 550082 401916 550084
rect 397637 550080 401916 550082
rect 397637 550024 397642 550080
rect 397698 550024 401916 550080
rect 397637 550022 401916 550024
rect 397637 550019 397703 550022
rect 401910 550020 401916 550022
rect 401980 550020 401986 550084
rect 401726 549266 401732 549268
rect 399894 549206 401732 549266
rect 399894 549032 399954 549206
rect 401726 549204 401732 549206
rect 401796 549204 401802 549268
rect 357525 548994 357591 548997
rect 360150 548994 360210 549032
rect 357525 548992 360210 548994
rect 357525 548936 357530 548992
rect 357586 548936 360210 548992
rect 357525 548934 360210 548936
rect 357525 548931 357591 548934
rect 358721 548858 358787 548861
rect 358721 548856 360210 548858
rect 358721 548800 358726 548856
rect 358782 548800 360210 548856
rect 358721 548798 360210 548800
rect 358721 548795 358787 548798
rect 360150 548352 360210 548798
rect 357433 547770 357499 547773
rect 402237 547770 402303 547773
rect 357433 547768 360210 547770
rect 357433 547712 357438 547768
rect 357494 547712 360210 547768
rect 357433 547710 360210 547712
rect 357433 547707 357499 547710
rect 360150 547672 360210 547710
rect 399894 547768 402303 547770
rect 399894 547712 402242 547768
rect 402298 547712 402303 547768
rect 399894 547710 402303 547712
rect 399894 547672 399954 547710
rect 402237 547707 402303 547710
rect 402421 547498 402487 547501
rect 399894 547496 402487 547498
rect 399894 547440 402426 547496
rect 402482 547440 402487 547496
rect 399894 547438 402487 547440
rect 358118 547362 358124 547364
rect 354630 547302 358124 547362
rect 254577 547090 254643 547093
rect 251804 547088 254643 547090
rect 251804 547032 254582 547088
rect 254638 547032 254643 547088
rect 251804 547030 254643 547032
rect 254577 547027 254643 547030
rect 329097 547090 329163 547093
rect 354630 547090 354690 547302
rect 358118 547300 358124 547302
rect 358188 547362 358194 547364
rect 358188 547302 360210 547362
rect 358188 547300 358194 547302
rect 329097 547088 354690 547090
rect 329097 547032 329102 547088
rect 329158 547032 354690 547088
rect 329097 547030 354690 547032
rect 329097 547027 329163 547030
rect 360150 546992 360210 547302
rect 399894 546992 399954 547438
rect 402421 547435 402487 547438
rect 402881 546410 402947 546413
rect 399894 546408 402947 546410
rect 399894 546352 402886 546408
rect 402942 546352 402947 546408
rect 399894 546350 402947 546352
rect 399894 546312 399954 546350
rect 402881 546347 402947 546350
rect 357433 546274 357499 546277
rect 357433 546272 360210 546274
rect 357433 546216 357438 546272
rect 357494 546216 360210 546272
rect 357433 546214 360210 546216
rect 357433 546211 357499 546214
rect 360150 545632 360210 546214
rect 402881 546138 402947 546141
rect 399894 546136 402947 546138
rect 399894 546080 402886 546136
rect 402942 546080 402947 546136
rect 399894 546078 402947 546080
rect 399894 545632 399954 546078
rect 402881 546075 402947 546078
rect 357893 545050 357959 545053
rect 357893 545048 360210 545050
rect 357893 544992 357898 545048
rect 357954 544992 360210 545048
rect 357893 544990 360210 544992
rect 357893 544987 357959 544990
rect 360150 544952 360210 544990
rect 357433 544778 357499 544781
rect 402053 544778 402119 544781
rect 357433 544776 360210 544778
rect 357433 544720 357438 544776
rect 357494 544720 360210 544776
rect 357433 544718 360210 544720
rect 357433 544715 357499 544718
rect 360150 544272 360210 544718
rect 399894 544776 402119 544778
rect 399894 544720 402058 544776
rect 402114 544720 402119 544776
rect 399894 544718 402119 544720
rect 399894 544272 399954 544718
rect 402053 544715 402119 544718
rect 49325 544098 49391 544101
rect 49325 544096 52164 544098
rect 49325 544040 49330 544096
rect 49386 544040 52164 544096
rect 49325 544038 52164 544040
rect 49325 544035 49391 544038
rect 295926 543628 295932 543692
rect 295996 543690 296002 543692
rect 306373 543690 306439 543693
rect 295996 543688 306439 543690
rect 295996 543632 306378 543688
rect 306434 543632 306439 543688
rect 295996 543630 306439 543632
rect 295996 543628 296002 543630
rect 306373 543627 306439 543630
rect 317505 543690 317571 543693
rect 317638 543690 317644 543692
rect 317505 543688 317644 543690
rect 317505 543632 317510 543688
rect 317566 543632 317644 543688
rect 317505 543630 317644 543632
rect 317505 543627 317571 543630
rect 317638 543628 317644 543630
rect 317708 543628 317714 543692
rect 401910 543690 401916 543692
rect 399894 543630 401916 543690
rect 399894 543592 399954 543630
rect 401910 543628 401916 543630
rect 401980 543628 401986 543692
rect 489862 543628 489868 543692
rect 489932 543690 489938 543692
rect 490741 543690 490807 543693
rect 489932 543688 490807 543690
rect 489932 543632 490746 543688
rect 490802 543632 490807 543688
rect 489932 543630 490807 543632
rect 489932 543628 489938 543630
rect 490741 543627 490807 543630
rect 295006 543492 295012 543556
rect 295076 543554 295082 543556
rect 307017 543554 307083 543557
rect 295076 543552 307083 543554
rect 295076 543496 307022 543552
rect 307078 543496 307083 543552
rect 295076 543494 307083 543496
rect 295076 543492 295082 543494
rect 307017 543491 307083 543494
rect 357709 543554 357775 543557
rect 358077 543554 358143 543557
rect 360150 543554 360210 543592
rect 357709 543552 360210 543554
rect 357709 543496 357714 543552
rect 357770 543496 358082 543552
rect 358138 543496 360210 543552
rect 357709 543494 360210 543496
rect 508313 543554 508379 543557
rect 508446 543554 508452 543556
rect 508313 543552 508452 543554
rect 508313 543496 508318 543552
rect 508374 543496 508452 543552
rect 508313 543494 508452 543496
rect 357709 543491 357775 543494
rect 358077 543491 358143 543494
rect 508313 543491 508379 543494
rect 508446 543492 508452 543494
rect 508516 543492 508522 543556
rect 286174 543356 286180 543420
rect 286244 543418 286250 543420
rect 297081 543418 297147 543421
rect 286244 543416 297147 543418
rect 286244 543360 297086 543416
rect 297142 543360 297147 543416
rect 286244 543358 297147 543360
rect 286244 543356 286250 543358
rect 297081 543355 297147 543358
rect 297214 543356 297220 543420
rect 297284 543418 297290 543420
rect 304993 543418 305059 543421
rect 297284 543416 305059 543418
rect 297284 543360 304998 543416
rect 305054 543360 305059 543416
rect 297284 543358 305059 543360
rect 297284 543356 297290 543358
rect 304993 543355 305059 543358
rect 358905 543418 358971 543421
rect 358905 543416 360210 543418
rect 358905 543360 358910 543416
rect 358966 543360 360210 543416
rect 358905 543358 360210 543360
rect 358905 543355 358971 543358
rect 283414 543220 283420 543284
rect 283484 543282 283490 543284
rect 300393 543282 300459 543285
rect 283484 543280 300459 543282
rect 283484 543224 300398 543280
rect 300454 543224 300459 543280
rect 283484 543222 300459 543224
rect 283484 543220 283490 543222
rect 300393 543219 300459 543222
rect 279366 543084 279372 543148
rect 279436 543146 279442 543148
rect 297449 543146 297515 543149
rect 279436 543144 297515 543146
rect 279436 543088 297454 543144
rect 297510 543088 297515 543144
rect 279436 543086 297515 543088
rect 279436 543084 279442 543086
rect 297449 543083 297515 543086
rect 311934 543084 311940 543148
rect 312004 543146 312010 543148
rect 312261 543146 312327 543149
rect 312004 543144 312327 543146
rect 312004 543088 312266 543144
rect 312322 543088 312327 543144
rect 312004 543086 312327 543088
rect 312004 543084 312010 543086
rect 312261 543083 312327 543086
rect 282310 542948 282316 543012
rect 282380 543010 282386 543012
rect 305545 543010 305611 543013
rect 282380 543008 305611 543010
rect 282380 542952 305550 543008
rect 305606 542952 305611 543008
rect 282380 542950 305611 542952
rect 282380 542948 282386 542950
rect 305545 542947 305611 542950
rect 360150 542912 360210 543358
rect 401777 543146 401843 543149
rect 399894 543144 401843 543146
rect 399894 543088 401782 543144
rect 401838 543088 401843 543144
rect 399894 543086 401843 543088
rect 399894 542912 399954 543086
rect 401777 543083 401843 543086
rect 272517 542874 272583 542877
rect 283465 542874 283531 542877
rect 272517 542872 283531 542874
rect 272517 542816 272522 542872
rect 272578 542816 283470 542872
rect 283526 542816 283531 542872
rect 272517 542814 283531 542816
rect 272517 542811 272583 542814
rect 283465 542811 283531 542814
rect 297081 542874 297147 542877
rect 301129 542874 301195 542877
rect 297081 542872 301195 542874
rect 297081 542816 297086 542872
rect 297142 542816 301134 542872
rect 301190 542816 301195 542872
rect 297081 542814 301195 542816
rect 297081 542811 297147 542814
rect 301129 542811 301195 542814
rect 282126 542676 282132 542740
rect 282196 542738 282202 542740
rect 296897 542738 296963 542741
rect 282196 542736 296963 542738
rect 282196 542680 296902 542736
rect 296958 542680 296963 542736
rect 282196 542678 296963 542680
rect 282196 542676 282202 542678
rect 296897 542675 296963 542678
rect 308397 542602 308463 542605
rect 308806 542602 308812 542604
rect 308397 542600 308812 542602
rect 308397 542544 308402 542600
rect 308458 542544 308812 542600
rect 308397 542542 308812 542544
rect 308397 542539 308463 542542
rect 308806 542540 308812 542542
rect 308876 542540 308882 542604
rect 309358 542540 309364 542604
rect 309428 542602 309434 542604
rect 309961 542602 310027 542605
rect 309428 542600 310027 542602
rect 309428 542544 309966 542600
rect 310022 542544 310027 542600
rect 309428 542542 310027 542544
rect 309428 542540 309434 542542
rect 309961 542539 310027 542542
rect 310462 542540 310468 542604
rect 310532 542602 310538 542604
rect 311433 542602 311499 542605
rect 310532 542600 311499 542602
rect 310532 542544 311438 542600
rect 311494 542544 311499 542600
rect 310532 542542 311499 542544
rect 310532 542540 310538 542542
rect 311433 542539 311499 542542
rect 308673 542468 308739 542469
rect 308622 542404 308628 542468
rect 308692 542466 308739 542468
rect 308692 542464 308784 542466
rect 308734 542408 308784 542464
rect 308692 542406 308784 542408
rect 308692 542404 308739 542406
rect 309174 542404 309180 542468
rect 309244 542466 309250 542468
rect 309409 542466 309475 542469
rect 311065 542468 311131 542469
rect 309244 542464 309475 542466
rect 309244 542408 309414 542464
rect 309470 542408 309475 542464
rect 309244 542406 309475 542408
rect 309244 542404 309250 542406
rect 308673 542403 308739 542404
rect 309409 542403 309475 542406
rect 311014 542404 311020 542468
rect 311084 542466 311131 542468
rect 311084 542464 311176 542466
rect 311126 542408 311176 542464
rect 311084 542406 311176 542408
rect 311084 542404 311131 542406
rect 311065 542403 311131 542404
rect 358445 542330 358511 542333
rect 358445 542328 360210 542330
rect 358445 542272 358450 542328
rect 358506 542272 360210 542328
rect 358445 542270 360210 542272
rect 358445 542267 358511 542270
rect 360150 542232 360210 542270
rect 359406 541996 359412 542060
rect 359476 542058 359482 542060
rect 359476 541998 360210 542058
rect 359476 541996 359482 541998
rect 254393 541242 254459 541245
rect 251804 541240 254459 541242
rect 251804 541184 254398 541240
rect 254454 541184 254459 541240
rect 251804 541182 254459 541184
rect 254393 541179 254459 541182
rect 345841 541106 345907 541109
rect 360150 541106 360210 541998
rect 399894 541786 399954 542232
rect 401777 541786 401843 541789
rect 399894 541784 401843 541786
rect 399894 541728 401782 541784
rect 401838 541728 401843 541784
rect 399894 541726 401843 541728
rect 401777 541723 401843 541726
rect 400121 541582 400187 541585
rect 399924 541580 400187 541582
rect 399924 541524 400126 541580
rect 400182 541524 400187 541580
rect 399924 541522 400187 541524
rect 400121 541519 400187 541522
rect 345841 541104 360210 541106
rect 345841 541048 345846 541104
rect 345902 541048 360210 541104
rect 345841 541046 360210 541048
rect 345841 541043 345907 541046
rect 495934 541044 495940 541108
rect 496004 541106 496010 541108
rect 498377 541106 498443 541109
rect 496004 541104 498443 541106
rect 496004 541048 498382 541104
rect 498438 541048 498443 541104
rect 496004 541046 498443 541048
rect 496004 541044 496010 541046
rect 498377 541043 498443 541046
rect 511206 541044 511212 541108
rect 511276 541106 511282 541108
rect 513833 541106 513899 541109
rect 511276 541104 513899 541106
rect 511276 541048 513838 541104
rect 513894 541048 513899 541104
rect 511276 541046 513899 541048
rect 511276 541044 511282 541046
rect 513833 541043 513899 541046
rect 358537 540970 358603 540973
rect 402053 540970 402119 540973
rect 358537 540968 360210 540970
rect -960 540684 480 540924
rect 358537 540912 358542 540968
rect 358598 540912 360210 540968
rect 358537 540910 360210 540912
rect 358537 540907 358603 540910
rect 360150 540872 360210 540910
rect 399894 540968 402119 540970
rect 399894 540912 402058 540968
rect 402114 540912 402119 540968
rect 399894 540910 402119 540912
rect 399894 540872 399954 540910
rect 402053 540907 402119 540910
rect 358302 540636 358308 540700
rect 358372 540698 358378 540700
rect 402329 540698 402395 540701
rect 358372 540638 360210 540698
rect 358372 540636 358378 540638
rect 360150 540192 360210 540638
rect 399894 540696 402395 540698
rect 399894 540640 402334 540696
rect 402390 540640 402395 540696
rect 399894 540638 402395 540640
rect 399894 540192 399954 540638
rect 402329 540635 402395 540638
rect 485630 539820 485636 539884
rect 485700 539882 485706 539884
rect 506749 539882 506815 539885
rect 485700 539880 506815 539882
rect 485700 539824 506754 539880
rect 506810 539824 506815 539880
rect 485700 539822 506815 539824
rect 485700 539820 485706 539822
rect 506749 539819 506815 539822
rect 512494 539820 512500 539884
rect 512564 539882 512570 539884
rect 517053 539882 517119 539885
rect 512564 539880 517119 539882
rect 512564 539824 517058 539880
rect 517114 539824 517119 539880
rect 512564 539822 517119 539824
rect 512564 539820 512570 539822
rect 517053 539819 517119 539822
rect 287278 539684 287284 539748
rect 287348 539746 287354 539748
rect 287881 539746 287947 539749
rect 287348 539744 287947 539746
rect 287348 539688 287886 539744
rect 287942 539688 287947 539744
rect 287348 539686 287947 539688
rect 287348 539684 287354 539686
rect 287881 539683 287947 539686
rect 288566 539684 288572 539748
rect 288636 539746 288642 539748
rect 289353 539746 289419 539749
rect 288636 539744 289419 539746
rect 288636 539688 289358 539744
rect 289414 539688 289419 539744
rect 288636 539686 289419 539688
rect 288636 539684 288642 539686
rect 289353 539683 289419 539686
rect 290590 539684 290596 539748
rect 290660 539746 290666 539748
rect 290825 539746 290891 539749
rect 290660 539744 290891 539746
rect 290660 539688 290830 539744
rect 290886 539688 290891 539744
rect 290660 539686 290891 539688
rect 290660 539684 290666 539686
rect 290825 539683 290891 539686
rect 486141 539746 486207 539749
rect 486366 539746 486372 539748
rect 486141 539744 486372 539746
rect 486141 539688 486146 539744
rect 486202 539688 486372 539744
rect 486141 539686 486372 539688
rect 486141 539683 486207 539686
rect 486366 539684 486372 539686
rect 486436 539684 486442 539748
rect 494646 539684 494652 539748
rect 494716 539746 494722 539748
rect 495801 539746 495867 539749
rect 494716 539744 495867 539746
rect 494716 539688 495806 539744
rect 495862 539688 495867 539744
rect 494716 539686 495867 539688
rect 494716 539684 494722 539686
rect 495801 539683 495867 539686
rect 502149 539748 502215 539749
rect 505553 539748 505619 539749
rect 516409 539748 516475 539749
rect 502149 539744 502196 539748
rect 502260 539746 502266 539748
rect 505502 539746 505508 539748
rect 502149 539688 502154 539744
rect 502149 539684 502196 539688
rect 502260 539686 502306 539746
rect 505462 539686 505508 539746
rect 505572 539744 505619 539748
rect 516358 539746 516364 539748
rect 505614 539688 505619 539744
rect 502260 539684 502266 539686
rect 505502 539684 505508 539686
rect 505572 539684 505619 539688
rect 516318 539686 516364 539746
rect 516428 539744 516475 539748
rect 516470 539688 516475 539744
rect 516358 539684 516364 539686
rect 516428 539684 516475 539688
rect 502149 539683 502215 539684
rect 505553 539683 505619 539684
rect 516409 539683 516475 539684
rect 283373 539610 283439 539613
rect 284886 539610 284892 539612
rect 283373 539608 284892 539610
rect 283373 539552 283378 539608
rect 283434 539552 284892 539608
rect 283373 539550 284892 539552
rect 283373 539547 283439 539550
rect 284886 539548 284892 539550
rect 284956 539548 284962 539612
rect 285990 539548 285996 539612
rect 286060 539610 286066 539612
rect 286133 539610 286199 539613
rect 286060 539608 286199 539610
rect 286060 539552 286138 539608
rect 286194 539552 286199 539608
rect 286060 539550 286199 539552
rect 286060 539548 286066 539550
rect 286133 539547 286199 539550
rect 287605 539612 287671 539613
rect 287605 539608 287652 539612
rect 287716 539610 287722 539612
rect 287605 539552 287610 539608
rect 287605 539548 287652 539552
rect 287716 539550 287762 539610
rect 287716 539548 287722 539550
rect 288382 539548 288388 539612
rect 288452 539610 288458 539612
rect 288617 539610 288683 539613
rect 288452 539608 288683 539610
rect 288452 539552 288622 539608
rect 288678 539552 288683 539608
rect 288452 539550 288683 539552
rect 288452 539548 288458 539550
rect 287605 539547 287671 539548
rect 288617 539547 288683 539550
rect 290733 539612 290799 539613
rect 290733 539608 290780 539612
rect 290844 539610 290850 539612
rect 290733 539552 290738 539608
rect 290733 539548 290780 539552
rect 290844 539550 290890 539610
rect 290844 539548 290850 539550
rect 291142 539548 291148 539612
rect 291212 539610 291218 539612
rect 291561 539610 291627 539613
rect 291212 539608 291627 539610
rect 291212 539552 291566 539608
rect 291622 539552 291627 539608
rect 291212 539550 291627 539552
rect 291212 539548 291218 539550
rect 290733 539547 290799 539548
rect 291561 539547 291627 539550
rect 292614 539548 292620 539612
rect 292684 539610 292690 539612
rect 293033 539610 293099 539613
rect 292684 539608 293099 539610
rect 292684 539552 293038 539608
rect 293094 539552 293099 539608
rect 292684 539550 293099 539552
rect 292684 539548 292690 539550
rect 293033 539547 293099 539550
rect 293902 539548 293908 539612
rect 293972 539610 293978 539612
rect 294505 539610 294571 539613
rect 293972 539608 294571 539610
rect 293972 539552 294510 539608
rect 294566 539552 294571 539608
rect 293972 539550 294571 539552
rect 293972 539548 293978 539550
rect 294505 539547 294571 539550
rect 295374 539548 295380 539612
rect 295444 539610 295450 539612
rect 295977 539610 296043 539613
rect 401542 539610 401548 539612
rect 295444 539608 296043 539610
rect 295444 539552 295982 539608
rect 296038 539552 296043 539608
rect 295444 539550 296043 539552
rect 295444 539548 295450 539550
rect 295977 539547 296043 539550
rect 399894 539550 401548 539610
rect 399894 539512 399954 539550
rect 401542 539548 401548 539550
rect 401612 539548 401618 539612
rect 357709 539338 357775 539341
rect 360150 539338 360210 539512
rect 400949 539338 401015 539341
rect 357709 539336 360210 539338
rect 357709 539280 357714 539336
rect 357770 539280 360210 539336
rect 357709 539278 360210 539280
rect 399894 539336 401015 539338
rect 399894 539280 400954 539336
rect 401010 539280 401015 539336
rect 399894 539278 401015 539280
rect 357709 539275 357775 539278
rect 357433 539202 357499 539205
rect 357433 539200 360210 539202
rect 357433 539144 357438 539200
rect 357494 539144 360210 539200
rect 357433 539142 360210 539144
rect 357433 539139 357499 539142
rect 360150 538832 360210 539142
rect 399894 538832 399954 539278
rect 400949 539275 401015 539278
rect 480118 538386 480178 539512
rect 519678 539069 519738 539512
rect 519629 539064 519738 539069
rect 519629 539008 519634 539064
rect 519690 539008 519738 539064
rect 519629 539006 519738 539008
rect 519629 539003 519695 539006
rect 519862 538522 519922 538832
rect 521878 538522 521884 538524
rect 519862 538462 521884 538522
rect 521878 538460 521884 538462
rect 521948 538460 521954 538524
rect 470550 538326 480178 538386
rect 51073 538250 51139 538253
rect 51073 538248 52164 538250
rect 51073 538192 51078 538248
rect 51134 538192 52164 538248
rect 51073 538190 52164 538192
rect 51073 538187 51139 538190
rect 404854 538188 404860 538252
rect 404924 538250 404930 538252
rect 470550 538250 470610 538326
rect 404924 538190 470610 538250
rect 404924 538188 404930 538190
rect 358261 538114 358327 538117
rect 360150 538114 360210 538152
rect 358261 538112 360210 538114
rect 358261 538056 358266 538112
rect 358322 538056 360210 538112
rect 358261 538054 360210 538056
rect 399894 538114 399954 538152
rect 401041 538114 401107 538117
rect 399894 538112 401107 538114
rect 399894 538056 401046 538112
rect 401102 538056 401107 538112
rect 399894 538054 401107 538056
rect 358261 538051 358327 538054
rect 401041 538051 401107 538054
rect 358629 537978 358695 537981
rect 358629 537976 360210 537978
rect 358629 537920 358634 537976
rect 358690 537920 360210 537976
rect 358629 537918 360210 537920
rect 358629 537915 358695 537918
rect 360150 537472 360210 537918
rect 400622 537842 400628 537844
rect 399894 537782 400628 537842
rect 399894 537472 399954 537782
rect 400622 537780 400628 537782
rect 400692 537780 400698 537844
rect 479057 537706 479123 537709
rect 480118 537706 480178 538152
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 479057 537704 480178 537706
rect 479057 537648 479062 537704
rect 479118 537648 480178 537704
rect 583520 537692 584960 537782
rect 479057 537646 480178 537648
rect 479057 537643 479123 537646
rect 320173 537366 320239 537369
rect 319884 537364 320239 537366
rect 319884 537308 320178 537364
rect 320234 537308 320239 537364
rect 319884 537306 320239 537308
rect 320173 537303 320239 537306
rect 399753 537026 399819 537029
rect 399710 537024 399819 537026
rect 399710 536968 399758 537024
rect 399814 536968 399819 537024
rect 399710 536963 399819 536968
rect 479333 537026 479399 537029
rect 480118 537026 480178 537472
rect 479333 537024 480178 537026
rect 479333 536968 479338 537024
rect 479394 536968 480178 537024
rect 479333 536966 480178 536968
rect 519862 537026 519922 537472
rect 522297 537026 522363 537029
rect 519862 537024 522363 537026
rect 519862 536968 522302 537024
rect 522358 536968 522363 537024
rect 519862 536966 522363 536968
rect 479333 536963 479399 536966
rect 522297 536963 522363 536966
rect 399710 536822 399770 536963
rect 399556 536792 399770 536822
rect 357433 536754 357499 536757
rect 360150 536754 360210 536792
rect 357433 536752 360210 536754
rect 357433 536696 357438 536752
rect 357494 536696 360210 536752
rect 357433 536694 360210 536696
rect 399526 536762 399740 536792
rect 357433 536691 357499 536694
rect 319854 536210 319914 536656
rect 357893 536618 357959 536621
rect 357893 536616 360210 536618
rect 357893 536560 357898 536616
rect 357954 536560 360210 536616
rect 357893 536558 360210 536560
rect 357893 536555 357959 536558
rect 322565 536210 322631 536213
rect 319854 536208 322631 536210
rect 319854 536152 322570 536208
rect 322626 536152 322631 536208
rect 319854 536150 322631 536152
rect 322565 536147 322631 536150
rect 360150 536112 360210 536558
rect 399526 536349 399586 536762
rect 399845 536618 399911 536621
rect 399845 536616 399954 536618
rect 399845 536560 399850 536616
rect 399906 536560 399954 536616
rect 399845 536555 399954 536560
rect 399526 536344 399635 536349
rect 399526 536288 399574 536344
rect 399630 536288 399635 536344
rect 399526 536286 399635 536288
rect 399569 536283 399635 536286
rect 399894 536112 399954 536555
rect 478597 536210 478663 536213
rect 480118 536210 480178 536792
rect 519862 536346 519922 536792
rect 522205 536346 522271 536349
rect 519862 536344 522271 536346
rect 519862 536288 522210 536344
rect 522266 536288 522271 536344
rect 519862 536286 522271 536288
rect 522205 536283 522271 536286
rect 478597 536208 480178 536210
rect 478597 536152 478602 536208
rect 478658 536152 480178 536208
rect 478597 536150 480178 536152
rect 478597 536147 478663 536150
rect 519862 535530 519922 536112
rect 521745 535530 521811 535533
rect 519862 535528 521811 535530
rect 519862 535472 521750 535528
rect 521806 535472 521811 535528
rect 519862 535470 521811 535472
rect 521745 535467 521811 535470
rect 254577 535394 254643 535397
rect 251804 535392 254643 535394
rect 251804 535336 254582 535392
rect 254638 535336 254643 535392
rect 251804 535334 254643 535336
rect 254577 535331 254643 535334
rect 357433 535394 357499 535397
rect 360150 535394 360210 535432
rect 357433 535392 360210 535394
rect 357433 535336 357438 535392
rect 357494 535336 360210 535392
rect 357433 535334 360210 535336
rect 399894 535394 399954 535432
rect 401593 535394 401659 535397
rect 399894 535392 401659 535394
rect 399894 535336 401598 535392
rect 401654 535336 401659 535392
rect 399894 535334 401659 535336
rect 357433 535331 357499 535334
rect 401593 535331 401659 535334
rect 478413 535394 478479 535397
rect 480118 535394 480178 535432
rect 478413 535392 480178 535394
rect 478413 535336 478418 535392
rect 478474 535336 480178 535392
rect 478413 535334 480178 535336
rect 478413 535331 478479 535334
rect 319854 535258 319914 535296
rect 322473 535258 322539 535261
rect 319854 535256 322539 535258
rect 319854 535200 322478 535256
rect 322534 535200 322539 535256
rect 319854 535198 322539 535200
rect 322473 535195 322539 535198
rect 357525 535258 357591 535261
rect 357525 535256 360210 535258
rect 357525 535200 357530 535256
rect 357586 535200 360210 535256
rect 357525 535198 360210 535200
rect 357525 535195 357591 535198
rect 322105 534986 322171 534989
rect 319854 534984 322171 534986
rect 319854 534928 322110 534984
rect 322166 534928 322171 534984
rect 319854 534926 322171 534928
rect 319854 534616 319914 534926
rect 322105 534923 322171 534926
rect 360150 534752 360210 535198
rect 402513 534714 402579 534717
rect 399894 534712 402579 534714
rect 399894 534656 402518 534712
rect 402574 534656 402579 534712
rect 399894 534654 402579 534656
rect 357893 534578 357959 534581
rect 357893 534576 360210 534578
rect 357893 534520 357898 534576
rect 357954 534520 360210 534576
rect 357893 534518 360210 534520
rect 357893 534515 357959 534518
rect 360150 534072 360210 534518
rect 399894 534072 399954 534654
rect 402513 534651 402579 534654
rect 477585 534306 477651 534309
rect 480118 534306 480178 534752
rect 477585 534304 480178 534306
rect 477585 534248 477590 534304
rect 477646 534248 480178 534304
rect 477585 534246 480178 534248
rect 519862 534306 519922 534752
rect 522205 534306 522271 534309
rect 519862 534304 522271 534306
rect 519862 534248 522210 534304
rect 522266 534248 522271 534304
rect 519862 534246 522271 534248
rect 477585 534243 477651 534246
rect 522205 534243 522271 534246
rect 478781 534170 478847 534173
rect 478781 534168 480178 534170
rect 478781 534112 478786 534168
rect 478842 534112 480178 534168
rect 478781 534110 480178 534112
rect 478781 534107 478847 534110
rect 480118 534072 480178 534110
rect 322841 534034 322907 534037
rect 319854 534032 322907 534034
rect 319854 533976 322846 534032
rect 322902 533976 322907 534032
rect 319854 533974 322907 533976
rect 319854 533936 319914 533974
rect 322841 533971 322907 533974
rect 519310 533900 519370 534072
rect 519302 533836 519308 533900
rect 519372 533836 519378 533900
rect 401593 533626 401659 533629
rect 399894 533624 401659 533626
rect 399894 533568 401598 533624
rect 401654 533568 401659 533624
rect 399894 533566 401659 533568
rect 357525 533490 357591 533493
rect 358353 533490 358419 533493
rect 357525 533488 360210 533490
rect 357525 533432 357530 533488
rect 357586 533432 358358 533488
rect 358414 533432 360210 533488
rect 357525 533430 360210 533432
rect 357525 533427 357591 533430
rect 358353 533427 358419 533430
rect 360150 533392 360210 533430
rect 399894 533392 399954 533566
rect 401593 533563 401659 533566
rect 322473 533354 322539 533357
rect 319854 533352 322539 533354
rect 319854 533296 322478 533352
rect 322534 533296 322539 533352
rect 319854 533294 322539 533296
rect 319854 533256 319914 533294
rect 322473 533291 322539 533294
rect 399937 533218 400003 533221
rect 399894 533216 400003 533218
rect 399894 533160 399942 533216
rect 399998 533160 400003 533216
rect 399894 533155 400003 533160
rect 358629 532810 358695 532813
rect 358629 532808 360210 532810
rect 358629 532752 358634 532808
rect 358690 532752 360210 532808
rect 358629 532750 360210 532752
rect 358629 532747 358695 532750
rect 360150 532712 360210 532750
rect 399894 532712 399954 533155
rect 477585 532810 477651 532813
rect 519862 532810 519922 533392
rect 522062 532810 522068 532812
rect 477585 532808 480178 532810
rect 477585 532752 477590 532808
rect 477646 532752 480178 532808
rect 477585 532750 480178 532752
rect 519862 532750 522068 532810
rect 477585 532747 477651 532750
rect 480118 532712 480178 532750
rect 522062 532748 522068 532750
rect 522132 532748 522138 532812
rect 49182 532340 49188 532404
rect 49252 532402 49258 532404
rect 49417 532402 49483 532405
rect 319854 532402 319914 532576
rect 400765 532538 400831 532541
rect 399894 532536 400831 532538
rect 399894 532480 400770 532536
rect 400826 532480 400831 532536
rect 399894 532478 400831 532480
rect 322749 532402 322815 532405
rect 49252 532400 52164 532402
rect 49252 532344 49422 532400
rect 49478 532344 52164 532400
rect 49252 532342 52164 532344
rect 319854 532400 322815 532402
rect 319854 532344 322754 532400
rect 322810 532344 322815 532400
rect 319854 532342 322815 532344
rect 49252 532340 49258 532342
rect 49417 532339 49483 532342
rect 322749 532339 322815 532342
rect 357433 532402 357499 532405
rect 357433 532400 360210 532402
rect 357433 532344 357438 532400
rect 357494 532344 360210 532400
rect 357433 532342 360210 532344
rect 357433 532339 357499 532342
rect 321645 532266 321711 532269
rect 319854 532264 321711 532266
rect 319854 532208 321650 532264
rect 321706 532208 321711 532264
rect 319854 532206 321711 532208
rect 319854 531896 319914 532206
rect 321645 532203 321711 532206
rect 360150 532032 360210 532342
rect 399894 532032 399954 532478
rect 400765 532475 400831 532478
rect 522941 532402 523007 532405
rect 519862 532400 523007 532402
rect 519862 532344 522946 532400
rect 523002 532344 523007 532400
rect 519862 532342 523007 532344
rect 519862 532032 519922 532342
rect 522941 532339 523007 532342
rect 357525 531858 357591 531861
rect 400806 531858 400812 531860
rect 357525 531856 360210 531858
rect 357525 531800 357530 531856
rect 357586 531800 360210 531856
rect 357525 531798 360210 531800
rect 357525 531795 357591 531798
rect 360150 531352 360210 531798
rect 399894 531798 400812 531858
rect 399894 531352 399954 531798
rect 400806 531796 400812 531798
rect 400876 531796 400882 531860
rect 405038 531524 405044 531588
rect 405108 531586 405114 531588
rect 480118 531586 480178 532032
rect 405108 531526 480178 531586
rect 405108 531524 405114 531526
rect 477585 531450 477651 531453
rect 477585 531448 480178 531450
rect 477585 531392 477590 531448
rect 477646 531392 480178 531448
rect 477585 531390 480178 531392
rect 477585 531387 477651 531390
rect 480118 531352 480178 531390
rect 322473 531314 322539 531317
rect 319854 531312 322539 531314
rect 319854 531256 322478 531312
rect 322534 531256 322539 531312
rect 319854 531254 322539 531256
rect 319854 531216 319914 531254
rect 322473 531251 322539 531254
rect 519494 531181 519554 531352
rect 519445 531176 519554 531181
rect 519445 531120 519450 531176
rect 519506 531120 519554 531176
rect 519445 531118 519554 531120
rect 519445 531115 519511 531118
rect 337929 530634 337995 530637
rect 353293 530634 353359 530637
rect 337929 530632 353359 530634
rect 337929 530576 337934 530632
rect 337990 530576 353298 530632
rect 353354 530576 353359 530632
rect 337929 530574 353359 530576
rect 337929 530571 337995 530574
rect 353293 530571 353359 530574
rect 359222 530572 359228 530636
rect 359292 530634 359298 530636
rect 359292 530574 360210 530634
rect 359292 530572 359298 530574
rect 319854 530226 319914 530536
rect 322565 530226 322631 530229
rect 319854 530224 322631 530226
rect 319854 530168 322570 530224
rect 322626 530168 322631 530224
rect 319854 530166 322631 530168
rect 322565 530163 322631 530166
rect 353293 529954 353359 529957
rect 353569 529954 353635 529957
rect 360150 529954 360210 530574
rect 399894 530362 399954 530672
rect 478689 530634 478755 530637
rect 478689 530632 480178 530634
rect 478689 530576 478694 530632
rect 478750 530576 480178 530632
rect 478689 530574 480178 530576
rect 478689 530571 478755 530574
rect 401777 530362 401843 530365
rect 399894 530360 401843 530362
rect 399894 530304 401782 530360
rect 401838 530304 401843 530360
rect 399894 530302 401843 530304
rect 401777 530299 401843 530302
rect 401593 530090 401659 530093
rect 399894 530088 401659 530090
rect 399894 530032 401598 530088
rect 401654 530032 401659 530088
rect 399894 530030 401659 530032
rect 399894 529992 399954 530030
rect 401593 530027 401659 530030
rect 480118 529992 480178 530574
rect 519494 530093 519554 530672
rect 519494 530088 519603 530093
rect 519494 530032 519542 530088
rect 519598 530032 519603 530088
rect 519494 530030 519603 530032
rect 519537 530027 519603 530030
rect 353293 529952 360210 529954
rect 353293 529896 353298 529952
rect 353354 529896 353574 529952
rect 353630 529896 360210 529952
rect 353293 529894 360210 529896
rect 353293 529891 353359 529894
rect 353569 529891 353635 529894
rect 319854 529818 319914 529856
rect 322473 529818 322539 529821
rect 319854 529816 322539 529818
rect 319854 529760 322478 529816
rect 322534 529760 322539 529816
rect 319854 529758 322539 529760
rect 322473 529755 322539 529758
rect 254577 529546 254643 529549
rect 251804 529544 254643 529546
rect 251804 529488 254582 529544
rect 254638 529488 254643 529544
rect 251804 529486 254643 529488
rect 254577 529483 254643 529486
rect 357433 529546 357499 529549
rect 357433 529544 360210 529546
rect 357433 529488 357438 529544
rect 357494 529488 360210 529544
rect 357433 529486 360210 529488
rect 357433 529483 357499 529486
rect 360150 529312 360210 529486
rect 319854 528866 319914 529176
rect 399894 529002 399954 529312
rect 401777 529002 401843 529005
rect 399894 529000 401843 529002
rect 399894 528944 401782 529000
rect 401838 528944 401843 529000
rect 399894 528942 401843 528944
rect 401777 528939 401843 528942
rect 477585 529002 477651 529005
rect 480118 529002 480178 529312
rect 477585 529000 480178 529002
rect 477585 528944 477590 529000
rect 477646 528944 480178 529000
rect 477585 528942 480178 528944
rect 519678 529005 519738 529312
rect 519678 529000 519787 529005
rect 519678 528944 519726 529000
rect 519782 528944 519787 529000
rect 519678 528942 519787 528944
rect 477585 528939 477651 528942
rect 519721 528939 519787 528942
rect 322841 528866 322907 528869
rect 401593 528866 401659 528869
rect 319854 528864 322907 528866
rect 319854 528808 322846 528864
rect 322902 528808 322907 528864
rect 319854 528806 322907 528808
rect 322841 528803 322907 528806
rect 399894 528864 401659 528866
rect 399894 528808 401598 528864
rect 401654 528808 401659 528864
rect 399894 528806 401659 528808
rect 399894 528632 399954 528806
rect 401593 528803 401659 528806
rect 358353 528594 358419 528597
rect 360150 528594 360210 528632
rect 358353 528592 360210 528594
rect 358353 528536 358358 528592
rect 358414 528536 360210 528592
rect 358353 528534 360210 528536
rect 401777 528594 401843 528597
rect 402053 528594 402119 528597
rect 401777 528592 402119 528594
rect 401777 528536 401782 528592
rect 401838 528536 402058 528592
rect 402114 528536 402119 528592
rect 401777 528534 402119 528536
rect 358353 528531 358419 528534
rect 401777 528531 401843 528534
rect 402053 528531 402119 528534
rect 478597 528594 478663 528597
rect 480118 528594 480178 528632
rect 478597 528592 480178 528594
rect 478597 528536 478602 528592
rect 478658 528536 480178 528592
rect 478597 528534 480178 528536
rect 519862 528594 519922 528632
rect 521009 528594 521075 528597
rect 519862 528592 521075 528594
rect 519862 528536 521014 528592
rect 521070 528536 521075 528592
rect 519862 528534 521075 528536
rect 478597 528531 478663 528534
rect 521009 528531 521075 528534
rect 319854 528458 319914 528496
rect 322473 528458 322539 528461
rect 319854 528456 322539 528458
rect 319854 528400 322478 528456
rect 322534 528400 322539 528456
rect 319854 528398 322539 528400
rect 322473 528395 322539 528398
rect 358169 528322 358235 528325
rect 358169 528320 360210 528322
rect 358169 528264 358174 528320
rect 358230 528264 360210 528320
rect 358169 528262 360210 528264
rect 358169 528259 358235 528262
rect 322105 528186 322171 528189
rect 319854 528184 322171 528186
rect 319854 528128 322110 528184
rect 322166 528128 322171 528184
rect 319854 528126 322171 528128
rect -960 527764 480 528004
rect 319854 527816 319914 528126
rect 322105 528123 322171 528126
rect 360150 527952 360210 528262
rect 401593 528186 401659 528189
rect 399894 528184 401659 528186
rect 399894 528128 401598 528184
rect 401654 528128 401659 528184
rect 399894 528126 401659 528128
rect 399894 527952 399954 528126
rect 401593 528123 401659 528126
rect 358670 527716 358676 527780
rect 358740 527778 358746 527780
rect 358740 527718 360210 527778
rect 358740 527716 358746 527718
rect 360150 527272 360210 527718
rect 399334 527716 399340 527780
rect 399404 527716 399410 527780
rect 399342 527272 399402 527716
rect 519862 527370 519922 527952
rect 520641 527370 520707 527373
rect 519862 527368 520707 527370
rect 519862 527312 520646 527368
rect 520702 527312 520707 527368
rect 519862 527310 520707 527312
rect 520641 527307 520707 527310
rect 477585 527234 477651 527237
rect 480118 527234 480178 527272
rect 477585 527232 480178 527234
rect 477585 527176 477590 527232
rect 477646 527176 480178 527232
rect 477585 527174 480178 527176
rect 477585 527171 477651 527174
rect 319854 527098 319914 527136
rect 322565 527098 322631 527101
rect 319854 527096 322631 527098
rect 319854 527040 322570 527096
rect 322626 527040 322631 527096
rect 319854 527038 322631 527040
rect 322565 527035 322631 527038
rect 357433 527098 357499 527101
rect 357433 527096 360210 527098
rect 357433 527040 357438 527096
rect 357494 527040 360210 527096
rect 357433 527038 360210 527040
rect 357433 527035 357499 527038
rect 322473 526826 322539 526829
rect 319854 526824 322539 526826
rect 319854 526768 322478 526824
rect 322534 526768 322539 526824
rect 319854 526766 322539 526768
rect 50981 526554 51047 526557
rect 50981 526552 52164 526554
rect 50981 526496 50986 526552
rect 51042 526496 52164 526552
rect 50981 526494 52164 526496
rect 50981 526491 51047 526494
rect 319854 526456 319914 526766
rect 322473 526763 322539 526766
rect 360150 526592 360210 527038
rect 477677 526826 477743 526829
rect 477677 526824 480178 526826
rect 477677 526768 477682 526824
rect 477738 526768 480178 526824
rect 477677 526766 480178 526768
rect 477677 526763 477743 526766
rect 400673 526690 400739 526693
rect 400446 526688 400739 526690
rect 400446 526632 400678 526688
rect 400734 526632 400739 526688
rect 400446 526630 400739 526632
rect 400446 526625 400506 526630
rect 400673 526627 400739 526630
rect 400397 526622 400506 526625
rect 399924 526620 400506 526622
rect 399924 526564 400402 526620
rect 400458 526564 400506 526620
rect 480118 526592 480178 526766
rect 520365 526622 520431 526625
rect 519892 526620 520431 526622
rect 399924 526562 400506 526564
rect 519892 526564 520370 526620
rect 520426 526564 520431 526620
rect 519892 526562 520431 526564
rect 400397 526559 400463 526562
rect 520365 526559 520431 526562
rect 357525 526418 357591 526421
rect 357525 526416 360210 526418
rect 357525 526360 357530 526416
rect 357586 526360 360210 526416
rect 357525 526358 360210 526360
rect 357525 526355 357591 526358
rect 360150 525912 360210 526358
rect 401593 526146 401659 526149
rect 399894 526144 401659 526146
rect 399894 526088 401598 526144
rect 401654 526088 401659 526144
rect 399894 526086 401659 526088
rect 399894 525912 399954 526086
rect 401593 526083 401659 526086
rect 477585 525874 477651 525877
rect 480118 525874 480178 525912
rect 477585 525872 480178 525874
rect 477585 525816 477590 525872
rect 477646 525816 480178 525872
rect 477585 525814 480178 525816
rect 519862 525874 519922 525912
rect 522941 525874 523007 525877
rect 519862 525872 523007 525874
rect 519862 525816 522946 525872
rect 523002 525816 523007 525872
rect 519862 525814 523007 525816
rect 477585 525811 477651 525814
rect 522941 525811 523007 525814
rect 319854 525738 319914 525776
rect 322289 525738 322355 525741
rect 319854 525736 322355 525738
rect 319854 525680 322294 525736
rect 322350 525680 322355 525736
rect 319854 525678 322355 525680
rect 322289 525675 322355 525678
rect 401593 525466 401659 525469
rect 399894 525464 401659 525466
rect 399894 525408 401598 525464
rect 401654 525408 401659 525464
rect 399894 525406 401659 525408
rect 399894 525232 399954 525406
rect 401593 525403 401659 525406
rect 319854 524650 319914 525096
rect 359549 524786 359615 524789
rect 360150 524786 360210 525232
rect 401593 524922 401659 524925
rect 359549 524784 360210 524786
rect 359549 524728 359554 524784
rect 359610 524728 360210 524784
rect 359549 524726 360210 524728
rect 399894 524920 401659 524922
rect 399894 524864 401598 524920
rect 401654 524864 401659 524920
rect 399894 524862 401659 524864
rect 359549 524723 359615 524726
rect 322105 524650 322171 524653
rect 319854 524648 322171 524650
rect 319854 524592 322110 524648
rect 322166 524592 322171 524648
rect 319854 524590 322171 524592
rect 322105 524587 322171 524590
rect 357801 524650 357867 524653
rect 357801 524648 360210 524650
rect 357801 524592 357806 524648
rect 357862 524592 360210 524648
rect 357801 524590 360210 524592
rect 357801 524587 357867 524590
rect 360150 524552 360210 524590
rect 399894 524552 399954 524862
rect 401593 524859 401659 524862
rect 478137 524922 478203 524925
rect 480118 524922 480178 525232
rect 478137 524920 480178 524922
rect 478137 524864 478142 524920
rect 478198 524864 480178 524920
rect 478137 524862 480178 524864
rect 478137 524859 478203 524862
rect 519862 524650 519922 525232
rect 521929 524650 521995 524653
rect 519862 524648 521995 524650
rect 519862 524592 521934 524648
rect 521990 524592 521995 524648
rect 519862 524590 521995 524592
rect 521929 524587 521995 524590
rect 322289 524514 322355 524517
rect 319854 524512 322355 524514
rect 319854 524456 322294 524512
rect 322350 524456 322355 524512
rect 319854 524454 322355 524456
rect 319854 524416 319914 524454
rect 322289 524451 322355 524454
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect 401593 524106 401659 524109
rect 399894 524104 401659 524106
rect 399894 524048 401598 524104
rect 401654 524048 401659 524104
rect 399894 524046 401659 524048
rect 399894 523872 399954 524046
rect 401593 524043 401659 524046
rect 357801 523834 357867 523837
rect 360150 523834 360210 523872
rect 357801 523832 360210 523834
rect 357801 523776 357806 523832
rect 357862 523776 360210 523832
rect 357801 523774 360210 523776
rect 357801 523771 357867 523774
rect 254301 523698 254367 523701
rect 251804 523696 254367 523698
rect 251804 523640 254306 523696
rect 254362 523640 254367 523696
rect 251804 523638 254367 523640
rect 254301 523635 254367 523638
rect 319854 523290 319914 523736
rect 357433 523698 357499 523701
rect 357433 523696 360210 523698
rect 357433 523640 357438 523696
rect 357494 523640 360210 523696
rect 357433 523638 360210 523640
rect 357433 523635 357499 523638
rect 322657 523290 322723 523293
rect 319854 523288 322723 523290
rect 319854 523232 322662 523288
rect 322718 523232 322723 523288
rect 319854 523230 322723 523232
rect 322657 523227 322723 523230
rect 360150 523192 360210 523638
rect 478413 523426 478479 523429
rect 480118 523426 480178 523872
rect 519310 523428 519370 523872
rect 478413 523424 480178 523426
rect 478413 523368 478418 523424
rect 478474 523368 480178 523424
rect 478413 523366 480178 523368
rect 478413 523363 478479 523366
rect 519302 523364 519308 523428
rect 519372 523364 519378 523428
rect 400438 523222 400444 523224
rect 399924 523162 400444 523222
rect 400438 523160 400444 523162
rect 400508 523160 400514 523224
rect 322473 523154 322539 523157
rect 319854 523152 322539 523154
rect 319854 523096 322478 523152
rect 322534 523096 322539 523152
rect 319854 523094 322539 523096
rect 319854 523056 319914 523094
rect 322473 523091 322539 523094
rect 478965 523154 479031 523157
rect 480118 523154 480178 523192
rect 478965 523152 480178 523154
rect 478965 523096 478970 523152
rect 479026 523096 480178 523152
rect 478965 523094 480178 523096
rect 519862 523154 519922 523192
rect 522941 523154 523007 523157
rect 519862 523152 523007 523154
rect 519862 523096 522946 523152
rect 523002 523096 523007 523152
rect 519862 523094 523007 523096
rect 478965 523091 479031 523094
rect 522941 523091 523007 523094
rect 401133 523018 401199 523021
rect 399894 523016 401199 523018
rect 399894 522960 401138 523016
rect 401194 522960 401199 523016
rect 399894 522958 401199 522960
rect 399894 522512 399954 522958
rect 401133 522955 401199 522958
rect 358537 522474 358603 522477
rect 360150 522474 360210 522512
rect 358537 522472 360210 522474
rect 358537 522416 358542 522472
rect 358598 522416 360210 522472
rect 358537 522414 360210 522416
rect 358537 522411 358603 522414
rect 319854 522338 319914 522376
rect 322197 522338 322263 522341
rect 319854 522336 322263 522338
rect 319854 522280 322202 522336
rect 322258 522280 322263 522336
rect 319854 522278 322263 522280
rect 322197 522275 322263 522278
rect 359089 522338 359155 522341
rect 359089 522336 360210 522338
rect 359089 522280 359094 522336
rect 359150 522280 360210 522336
rect 359089 522278 360210 522280
rect 359089 522275 359155 522278
rect 322565 522202 322631 522205
rect 319854 522200 322631 522202
rect 319854 522144 322570 522200
rect 322626 522144 322631 522200
rect 319854 522142 322631 522144
rect 319854 521696 319914 522142
rect 322565 522139 322631 522142
rect 360150 521832 360210 522278
rect 478781 521930 478847 521933
rect 480118 521930 480178 522512
rect 478781 521928 480178 521930
rect 478781 521872 478786 521928
rect 478842 521872 480178 521928
rect 478781 521870 480178 521872
rect 519862 521930 519922 522512
rect 522481 521930 522547 521933
rect 519862 521928 522547 521930
rect 519862 521872 522486 521928
rect 522542 521872 522547 521928
rect 519862 521870 522547 521872
rect 478781 521867 478847 521870
rect 522481 521867 522547 521870
rect 399894 521794 399954 521832
rect 401593 521794 401659 521797
rect 399894 521792 401659 521794
rect 399894 521736 401598 521792
rect 401654 521736 401659 521792
rect 399894 521734 401659 521736
rect 401593 521731 401659 521734
rect 357617 521658 357683 521661
rect 401961 521658 402027 521661
rect 357617 521656 360210 521658
rect 357617 521600 357622 521656
rect 357678 521600 360210 521656
rect 357617 521598 360210 521600
rect 357617 521595 357683 521598
rect 360150 521152 360210 521598
rect 399894 521656 402027 521658
rect 399894 521600 401966 521656
rect 402022 521600 402027 521656
rect 399894 521598 402027 521600
rect 399894 521152 399954 521598
rect 401961 521595 402027 521598
rect 50889 520706 50955 520709
rect 319854 520706 319914 521016
rect 359181 520978 359247 520981
rect 359181 520976 360210 520978
rect 359181 520920 359186 520976
rect 359242 520920 360210 520976
rect 359181 520918 360210 520920
rect 359181 520915 359247 520918
rect 322013 520706 322079 520709
rect 50889 520704 52164 520706
rect 50889 520648 50894 520704
rect 50950 520648 52164 520704
rect 50889 520646 52164 520648
rect 319854 520704 322079 520706
rect 319854 520648 322018 520704
rect 322074 520648 322079 520704
rect 319854 520646 322079 520648
rect 50889 520643 50955 520646
rect 322013 520643 322079 520646
rect 322473 520570 322539 520573
rect 319854 520568 322539 520570
rect 319854 520512 322478 520568
rect 322534 520512 322539 520568
rect 319854 520510 322539 520512
rect 319854 520336 319914 520510
rect 322473 520507 322539 520510
rect 360150 520472 360210 520918
rect 401593 520842 401659 520845
rect 399894 520840 401659 520842
rect 399894 520784 401598 520840
rect 401654 520784 401659 520840
rect 399894 520782 401659 520784
rect 399894 520472 399954 520782
rect 401593 520779 401659 520782
rect 478505 520706 478571 520709
rect 480118 520706 480178 521152
rect 519862 520978 519922 521152
rect 522941 520978 523007 520981
rect 519862 520976 523007 520978
rect 519862 520920 522946 520976
rect 523002 520920 523007 520976
rect 519862 520918 523007 520920
rect 522941 520915 523007 520918
rect 478505 520704 480178 520706
rect 478505 520648 478510 520704
rect 478566 520648 480178 520704
rect 478505 520646 480178 520648
rect 478505 520643 478571 520646
rect 477861 520298 477927 520301
rect 480118 520298 480178 520472
rect 477861 520296 480178 520298
rect 477861 520240 477866 520296
rect 477922 520240 480178 520296
rect 477861 520238 480178 520240
rect 519862 520298 519922 520472
rect 521101 520298 521167 520301
rect 519862 520296 521167 520298
rect 519862 520240 521106 520296
rect 521162 520240 521167 520296
rect 519862 520238 521167 520240
rect 477861 520235 477927 520238
rect 521101 520235 521167 520238
rect 520549 520162 520615 520165
rect 519862 520160 520615 520162
rect 519862 520104 520554 520160
rect 520610 520104 520615 520160
rect 519862 520102 520615 520104
rect 401593 520026 401659 520029
rect 399894 520024 401659 520026
rect 399894 519968 401598 520024
rect 401654 519968 401659 520024
rect 399894 519966 401659 519968
rect 399894 519792 399954 519966
rect 401593 519963 401659 519966
rect 519862 519792 519922 520102
rect 520549 520099 520615 520102
rect 358077 519754 358143 519757
rect 360150 519754 360210 519792
rect 358077 519752 360210 519754
rect 358077 519696 358082 519752
rect 358138 519696 360210 519752
rect 358077 519694 360210 519696
rect 358077 519691 358143 519694
rect 319854 519618 319914 519656
rect 322197 519618 322263 519621
rect 319854 519616 322263 519618
rect 319854 519560 322202 519616
rect 322258 519560 322263 519616
rect 319854 519558 322263 519560
rect 322197 519555 322263 519558
rect 357433 519618 357499 519621
rect 357433 519616 360210 519618
rect 357433 519560 357438 519616
rect 357494 519560 360210 519616
rect 357433 519558 360210 519560
rect 357433 519555 357499 519558
rect 321645 519482 321711 519485
rect 319854 519480 321711 519482
rect 319854 519424 321650 519480
rect 321706 519424 321711 519480
rect 319854 519422 321711 519424
rect 319854 518976 319914 519422
rect 321645 519419 321711 519422
rect 360150 519112 360210 519558
rect 477585 519346 477651 519349
rect 480118 519346 480178 519792
rect 477585 519344 480178 519346
rect 477585 519288 477590 519344
rect 477646 519288 480178 519344
rect 477585 519286 480178 519288
rect 477585 519283 477651 519286
rect 324221 518938 324287 518941
rect 349102 518938 349108 518940
rect 324221 518936 349108 518938
rect 324221 518880 324226 518936
rect 324282 518880 349108 518936
rect 324221 518878 349108 518880
rect 324221 518875 324287 518878
rect 349102 518876 349108 518878
rect 349172 518876 349178 518940
rect 357433 518802 357499 518805
rect 357433 518800 360210 518802
rect 357433 518744 357438 518800
rect 357494 518744 360210 518800
rect 357433 518742 360210 518744
rect 357433 518739 357499 518742
rect 360150 518432 360210 518742
rect 399334 518604 399340 518668
rect 399404 518604 399410 518668
rect 399342 518432 399402 518604
rect 520089 518462 520155 518465
rect 519892 518460 520155 518462
rect 319854 517986 319914 518296
rect 322289 517986 322355 517989
rect 319854 517984 322355 517986
rect 319854 517928 322294 517984
rect 322350 517928 322355 517984
rect 319854 517926 322355 517928
rect 322289 517923 322355 517926
rect 477585 517986 477651 517989
rect 480118 517986 480178 518432
rect 519892 518404 520094 518460
rect 520150 518404 520155 518460
rect 519892 518402 520155 518404
rect 520089 518399 520155 518402
rect 477585 517984 480178 517986
rect 477585 517928 477590 517984
rect 477646 517928 480178 517984
rect 477585 517926 480178 517928
rect 477585 517923 477651 517926
rect 254577 517850 254643 517853
rect 321737 517850 321803 517853
rect 251804 517848 254643 517850
rect 251804 517792 254582 517848
rect 254638 517792 254643 517848
rect 251804 517790 254643 517792
rect 254577 517787 254643 517790
rect 319854 517848 321803 517850
rect 319854 517792 321742 517848
rect 321798 517792 321803 517848
rect 319854 517790 321803 517792
rect 319854 517616 319914 517790
rect 321737 517787 321803 517790
rect 400305 517782 400371 517785
rect 399924 517780 400371 517782
rect 357525 517578 357591 517581
rect 360150 517578 360210 517752
rect 399924 517724 400310 517780
rect 400366 517724 400371 517780
rect 399924 517722 400371 517724
rect 400305 517719 400371 517722
rect 477677 517714 477743 517717
rect 480118 517714 480178 517752
rect 477677 517712 480178 517714
rect 477677 517656 477682 517712
rect 477738 517656 480178 517712
rect 477677 517654 480178 517656
rect 477677 517651 477743 517654
rect 357525 517576 360210 517578
rect 357525 517520 357530 517576
rect 357586 517520 360210 517576
rect 357525 517518 360210 517520
rect 519862 517578 519922 517752
rect 520549 517578 520615 517581
rect 519862 517576 520615 517578
rect 519862 517520 520554 517576
rect 520610 517520 520615 517576
rect 519862 517518 520615 517520
rect 357525 517515 357591 517518
rect 520549 517515 520615 517518
rect 322749 517442 322815 517445
rect 319854 517440 322815 517442
rect 319854 517384 322754 517440
rect 322810 517384 322815 517440
rect 319854 517382 322815 517384
rect 319854 516936 319914 517382
rect 322749 517379 322815 517382
rect 357433 517442 357499 517445
rect 401685 517442 401751 517445
rect 522021 517442 522087 517445
rect 357433 517440 360210 517442
rect 357433 517384 357438 517440
rect 357494 517384 360210 517440
rect 357433 517382 360210 517384
rect 357433 517379 357499 517382
rect 360150 517072 360210 517382
rect 399894 517440 401751 517442
rect 399894 517384 401690 517440
rect 401746 517384 401751 517440
rect 399894 517382 401751 517384
rect 399894 517072 399954 517382
rect 401685 517379 401751 517382
rect 519862 517440 522087 517442
rect 519862 517384 522026 517440
rect 522082 517384 522087 517440
rect 519862 517382 522087 517384
rect 477585 517306 477651 517309
rect 477585 517304 480178 517306
rect 477585 517248 477590 517304
rect 477646 517248 480178 517304
rect 477585 517246 480178 517248
rect 477585 517243 477651 517246
rect 480118 517072 480178 517246
rect 519862 517072 519922 517382
rect 522021 517379 522087 517382
rect 358486 516898 358492 516900
rect 354630 516838 358492 516898
rect 322841 516762 322907 516765
rect 319854 516760 322907 516762
rect 319854 516704 322846 516760
rect 322902 516704 322907 516760
rect 319854 516702 322907 516704
rect 319854 516256 319914 516702
rect 322841 516699 322907 516702
rect 331213 516762 331279 516765
rect 354630 516762 354690 516838
rect 358486 516836 358492 516838
rect 358556 516898 358562 516900
rect 358556 516838 360210 516898
rect 358556 516836 358562 516838
rect 331213 516760 354690 516762
rect 331213 516704 331218 516760
rect 331274 516704 354690 516760
rect 331213 516702 354690 516704
rect 331213 516699 331279 516702
rect 360150 516392 360210 516838
rect 399894 516354 399954 516392
rect 401593 516354 401659 516357
rect 399894 516352 401659 516354
rect 399894 516296 401598 516352
rect 401654 516296 401659 516352
rect 399894 516294 401659 516296
rect 401593 516291 401659 516294
rect 401685 515946 401751 515949
rect 399894 515944 401751 515946
rect 399894 515888 401690 515944
rect 401746 515888 401751 515944
rect 399894 515886 401751 515888
rect 399894 515712 399954 515886
rect 401685 515883 401751 515886
rect 319854 515538 319914 515576
rect 322841 515538 322907 515541
rect 319854 515536 322907 515538
rect 319854 515480 322846 515536
rect 322902 515480 322907 515536
rect 319854 515478 322907 515480
rect 322841 515475 322907 515478
rect 322289 515402 322355 515405
rect 319854 515400 322355 515402
rect 319854 515344 322294 515400
rect 322350 515344 322355 515400
rect 319854 515342 322355 515344
rect -960 514858 480 514948
rect 319854 514896 319914 515342
rect 322289 515339 322355 515342
rect 358169 515130 358235 515133
rect 360150 515130 360210 515712
rect 477677 515266 477743 515269
rect 480118 515266 480178 515712
rect 519862 515674 519922 515712
rect 520917 515674 520983 515677
rect 519862 515672 520983 515674
rect 519862 515616 520922 515672
rect 520978 515616 520983 515672
rect 519862 515614 520983 515616
rect 520917 515611 520983 515614
rect 520457 515538 520523 515541
rect 477677 515264 480178 515266
rect 477677 515208 477682 515264
rect 477738 515208 480178 515264
rect 477677 515206 480178 515208
rect 519862 515536 520523 515538
rect 519862 515480 520462 515536
rect 520518 515480 520523 515536
rect 519862 515478 520523 515480
rect 477677 515203 477743 515206
rect 358169 515128 360210 515130
rect 358169 515072 358174 515128
rect 358230 515072 360210 515128
rect 358169 515070 360210 515072
rect 358169 515067 358235 515070
rect 519862 515032 519922 515478
rect 520457 515475 520523 515478
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 51165 514858 51231 514861
rect 399894 514858 399954 515032
rect 477585 514994 477651 514997
rect 480118 514994 480178 515032
rect 477585 514992 480178 514994
rect 477585 514936 477590 514992
rect 477646 514936 480178 514992
rect 477585 514934 480178 514936
rect 477585 514931 477651 514934
rect 400489 514858 400555 514861
rect 402329 514858 402395 514861
rect 51165 514856 52164 514858
rect 51165 514800 51170 514856
rect 51226 514800 52164 514856
rect 51165 514798 52164 514800
rect 399894 514856 402395 514858
rect 399894 514800 400494 514856
rect 400550 514800 402334 514856
rect 402390 514800 402395 514856
rect 399894 514798 402395 514800
rect 51165 514795 51231 514798
rect 400489 514795 400555 514798
rect 402329 514795 402395 514798
rect 357433 514722 357499 514725
rect 357433 514720 360210 514722
rect 357433 514664 357438 514720
rect 357494 514664 360210 514720
rect 357433 514662 360210 514664
rect 357433 514659 357499 514662
rect 360150 514352 360210 514662
rect 319854 514178 319914 514216
rect 322749 514178 322815 514181
rect 319854 514176 322815 514178
rect 319854 514120 322754 514176
rect 322810 514120 322815 514176
rect 319854 514118 322815 514120
rect 322749 514115 322815 514118
rect 399894 513906 399954 514352
rect 401685 513906 401751 513909
rect 399894 513904 401751 513906
rect 399894 513848 401690 513904
rect 401746 513848 401751 513904
rect 399894 513846 401751 513848
rect 401685 513843 401751 513846
rect 477585 513906 477651 513909
rect 480118 513906 480178 514352
rect 477585 513904 480178 513906
rect 477585 513848 477590 513904
rect 477646 513848 480178 513904
rect 477585 513846 480178 513848
rect 477585 513843 477651 513846
rect 519862 513770 519922 514352
rect 522021 513770 522087 513773
rect 519862 513768 522087 513770
rect 519862 513712 522026 513768
rect 522082 513712 522087 513768
rect 519862 513710 522087 513712
rect 522021 513707 522087 513710
rect 319854 513498 319914 513536
rect 322289 513498 322355 513501
rect 319854 513496 322355 513498
rect 319854 513440 322294 513496
rect 322350 513440 322355 513496
rect 319854 513438 322355 513440
rect 322289 513435 322355 513438
rect 357525 513498 357591 513501
rect 360150 513498 360210 513672
rect 357525 513496 360210 513498
rect 357525 513440 357530 513496
rect 357586 513440 360210 513496
rect 357525 513438 360210 513440
rect 399894 513498 399954 513672
rect 401961 513498 402027 513501
rect 399894 513496 402027 513498
rect 399894 513440 401966 513496
rect 402022 513440 402027 513496
rect 399894 513438 402027 513440
rect 357525 513435 357591 513438
rect 401961 513435 402027 513438
rect 358997 513362 359063 513365
rect 403014 513362 403020 513364
rect 358997 513360 360210 513362
rect 358997 513304 359002 513360
rect 359058 513304 360210 513360
rect 358997 513302 360210 513304
rect 358997 513299 359063 513302
rect 360150 512992 360210 513302
rect 399894 513302 403020 513362
rect 399894 512992 399954 513302
rect 403014 513300 403020 513302
rect 403084 513300 403090 513364
rect 522849 513226 522915 513229
rect 519862 513224 522915 513226
rect 519862 513168 522854 513224
rect 522910 513168 522915 513224
rect 519862 513166 522915 513168
rect 519862 512992 519922 513166
rect 522849 513163 522915 513166
rect 319854 512682 319914 512856
rect 357433 512818 357499 512821
rect 402421 512818 402487 512821
rect 357433 512816 360210 512818
rect 357433 512760 357438 512816
rect 357494 512760 360210 512816
rect 357433 512758 360210 512760
rect 357433 512755 357499 512758
rect 321737 512682 321803 512685
rect 322197 512682 322263 512685
rect 319854 512680 322263 512682
rect 319854 512624 321742 512680
rect 321798 512624 322202 512680
rect 322258 512624 322263 512680
rect 319854 512622 322263 512624
rect 321737 512619 321803 512622
rect 322197 512619 322263 512622
rect 360150 512312 360210 512758
rect 399894 512816 402487 512818
rect 399894 512760 402426 512816
rect 402482 512760 402487 512816
rect 399894 512758 402487 512760
rect 399894 512312 399954 512758
rect 402421 512755 402487 512758
rect 477677 512546 477743 512549
rect 480118 512546 480178 512992
rect 521837 512818 521903 512821
rect 477677 512544 480178 512546
rect 477677 512488 477682 512544
rect 477738 512488 480178 512544
rect 477677 512486 480178 512488
rect 519862 512816 521903 512818
rect 519862 512760 521842 512816
rect 521898 512760 521903 512816
rect 519862 512758 521903 512760
rect 477677 512483 477743 512486
rect 519862 512312 519922 512758
rect 521837 512755 521903 512758
rect 319854 512138 319914 512176
rect 322197 512138 322263 512141
rect 319854 512136 322263 512138
rect 319854 512080 322202 512136
rect 322258 512080 322263 512136
rect 319854 512078 322263 512080
rect 322197 512075 322263 512078
rect 478137 512138 478203 512141
rect 480118 512138 480178 512312
rect 478137 512136 480178 512138
rect 478137 512080 478142 512136
rect 478198 512080 480178 512136
rect 478137 512078 480178 512080
rect 478137 512075 478203 512078
rect 254393 512002 254459 512005
rect 251804 512000 254459 512002
rect 251804 511944 254398 512000
rect 254454 511944 254459 512000
rect 251804 511942 254459 511944
rect 254393 511939 254459 511942
rect 477585 511866 477651 511869
rect 477585 511864 480178 511866
rect 477585 511808 477590 511864
rect 477646 511808 480178 511864
rect 477585 511806 480178 511808
rect 477585 511803 477651 511806
rect 400213 511662 400279 511665
rect 399924 511660 400279 511662
rect 357893 511594 357959 511597
rect 360150 511594 360210 511632
rect 399924 511604 400218 511660
rect 400274 511604 400279 511660
rect 480118 511632 480178 511806
rect 399924 511602 400279 511604
rect 400213 511599 400279 511602
rect 357893 511592 360210 511594
rect 357893 511536 357898 511592
rect 357954 511536 360210 511592
rect 357893 511534 360210 511536
rect 357893 511531 357959 511534
rect 319854 511322 319914 511496
rect 357433 511458 357499 511461
rect 357433 511456 360210 511458
rect 357433 511400 357438 511456
rect 357494 511400 360210 511456
rect 357433 511398 360210 511400
rect 357433 511395 357499 511398
rect 321553 511322 321619 511325
rect 319854 511320 321619 511322
rect 319854 511264 321558 511320
rect 321614 511264 321619 511320
rect 319854 511262 321619 511264
rect 321553 511259 321619 511262
rect 360150 510952 360210 511398
rect 519862 511186 519922 511632
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 522941 511186 523007 511189
rect 519862 511184 523007 511186
rect 519862 511128 522946 511184
rect 523002 511128 523007 511184
rect 583520 511172 584960 511262
rect 519862 511126 523007 511128
rect 522941 511123 523007 511126
rect 320081 510846 320147 510849
rect 319884 510844 320147 510846
rect 319884 510788 320086 510844
rect 320142 510788 320147 510844
rect 319884 510786 320147 510788
rect 320081 510783 320147 510786
rect 399894 510778 399954 510952
rect 402881 510778 402947 510781
rect 399894 510776 402947 510778
rect 399894 510720 402886 510776
rect 402942 510720 402947 510776
rect 399894 510718 402947 510720
rect 402881 510715 402947 510718
rect 519862 510642 519922 510952
rect 522573 510642 522639 510645
rect 519862 510640 522639 510642
rect 519862 510584 522578 510640
rect 522634 510584 522639 510640
rect 519862 510582 522639 510584
rect 522573 510579 522639 510582
rect 357433 510506 357499 510509
rect 402145 510506 402211 510509
rect 357433 510504 360210 510506
rect 357433 510448 357438 510504
rect 357494 510448 360210 510504
rect 357433 510446 360210 510448
rect 357433 510443 357499 510446
rect 360150 510272 360210 510446
rect 399894 510504 402211 510506
rect 399894 510448 402150 510504
rect 402206 510448 402211 510504
rect 399894 510446 402211 510448
rect 399894 510272 399954 510446
rect 402145 510443 402211 510446
rect 478137 510506 478203 510509
rect 478137 510504 480178 510506
rect 478137 510448 478142 510504
rect 478198 510448 480178 510504
rect 478137 510446 480178 510448
rect 478137 510443 478203 510446
rect 480118 510272 480178 510446
rect 521653 510234 521719 510237
rect 519862 510232 521719 510234
rect 519862 510176 521658 510232
rect 521714 510176 521719 510232
rect 519862 510174 521719 510176
rect 319854 509690 319914 510136
rect 358813 510098 358879 510101
rect 358813 510096 360210 510098
rect 358813 510040 358818 510096
rect 358874 510040 360210 510096
rect 358813 510038 360210 510040
rect 358813 510035 358879 510038
rect 321645 509690 321711 509693
rect 319854 509688 321711 509690
rect 319854 509632 321650 509688
rect 321706 509632 321711 509688
rect 319854 509630 321711 509632
rect 321645 509627 321711 509630
rect 360150 509592 360210 510038
rect 519862 509592 519922 510174
rect 521653 510171 521719 510174
rect 320357 509486 320423 509489
rect 319884 509484 320423 509486
rect 319884 509428 320362 509484
rect 320418 509428 320423 509484
rect 319884 509426 320423 509428
rect 320357 509423 320423 509426
rect 399894 509418 399954 509592
rect 402881 509418 402947 509421
rect 399894 509416 402947 509418
rect 399894 509360 402886 509416
rect 402942 509360 402947 509416
rect 399894 509358 402947 509360
rect 402881 509355 402947 509358
rect 477585 509418 477651 509421
rect 480118 509418 480178 509592
rect 477585 509416 480178 509418
rect 477585 509360 477590 509416
rect 477646 509360 480178 509416
rect 477585 509358 480178 509360
rect 477585 509355 477651 509358
rect 51257 509010 51323 509013
rect 357433 509010 357499 509013
rect 51257 509008 52164 509010
rect 51257 508952 51262 509008
rect 51318 508952 52164 509008
rect 51257 508950 52164 508952
rect 357433 509008 360210 509010
rect 357433 508952 357438 509008
rect 357494 508952 360210 509008
rect 357433 508950 360210 508952
rect 51257 508947 51323 508950
rect 357433 508947 357499 508950
rect 360150 508912 360210 508950
rect 520365 508942 520431 508945
rect 519892 508940 520431 508942
rect 319302 508333 319362 508776
rect 357985 508738 358051 508741
rect 357985 508736 360210 508738
rect 357985 508680 357990 508736
rect 358046 508680 360210 508736
rect 357985 508678 360210 508680
rect 357985 508675 358051 508678
rect 319302 508328 319411 508333
rect 319302 508272 319350 508328
rect 319406 508272 319411 508328
rect 319302 508270 319411 508272
rect 319345 508267 319411 508270
rect 360150 508232 360210 508678
rect 399894 508466 399954 508912
rect 402053 508466 402119 508469
rect 399894 508464 402119 508466
rect 399894 508408 402058 508464
rect 402114 508408 402119 508464
rect 399894 508406 402119 508408
rect 402053 508403 402119 508406
rect 478137 508466 478203 508469
rect 480118 508466 480178 508912
rect 519892 508884 520370 508940
rect 520426 508884 520431 508940
rect 519892 508882 520431 508884
rect 520365 508879 520431 508882
rect 520733 508738 520799 508741
rect 478137 508464 480178 508466
rect 478137 508408 478142 508464
rect 478198 508408 480178 508464
rect 478137 508406 480178 508408
rect 519862 508736 520799 508738
rect 519862 508680 520738 508736
rect 520794 508680 520799 508736
rect 519862 508678 520799 508680
rect 478137 508403 478203 508406
rect 401869 508330 401935 508333
rect 399894 508328 401935 508330
rect 399894 508272 401874 508328
rect 401930 508272 401935 508328
rect 399894 508270 401935 508272
rect 399894 508232 399954 508270
rect 401869 508267 401935 508270
rect 519862 508232 519922 508678
rect 520733 508675 520799 508678
rect 320265 508126 320331 508129
rect 319884 508124 320331 508126
rect 319884 508068 320270 508124
rect 320326 508068 320331 508124
rect 319884 508066 320331 508068
rect 320265 508063 320331 508066
rect 358445 507786 358511 507789
rect 358445 507784 360210 507786
rect 358445 507728 358450 507784
rect 358506 507728 360210 507784
rect 358445 507726 360210 507728
rect 358445 507723 358511 507726
rect 360150 507552 360210 507726
rect 399334 507724 399340 507788
rect 399404 507724 399410 507788
rect 399342 507552 399402 507724
rect 320265 507446 320331 507449
rect 319884 507444 320331 507446
rect 319884 507388 320270 507444
rect 320326 507388 320331 507444
rect 319884 507386 320331 507388
rect 320265 507383 320331 507386
rect 357433 507378 357499 507381
rect 399477 507378 399543 507381
rect 357433 507376 360210 507378
rect 357433 507320 357438 507376
rect 357494 507320 360210 507376
rect 357433 507318 360210 507320
rect 357433 507315 357499 507318
rect 360150 506872 360210 507318
rect 399477 507376 399586 507378
rect 399477 507320 399482 507376
rect 399538 507320 399586 507376
rect 399477 507315 399586 507320
rect 399526 506872 399586 507315
rect 479241 507106 479307 507109
rect 480118 507106 480178 507552
rect 479241 507104 480178 507106
rect 479241 507048 479246 507104
rect 479302 507048 480178 507104
rect 479241 507046 480178 507048
rect 479241 507043 479307 507046
rect 322381 506834 322447 506837
rect 319302 506832 322447 506834
rect 319302 506776 322386 506832
rect 322442 506776 322447 506832
rect 319302 506774 322447 506776
rect 319302 506565 319362 506774
rect 322381 506771 322447 506774
rect 477493 506698 477559 506701
rect 480118 506698 480178 506872
rect 477493 506696 480178 506698
rect 477493 506640 477498 506696
rect 477554 506640 480178 506696
rect 477493 506638 480178 506640
rect 477493 506635 477559 506638
rect 319302 506560 319411 506565
rect 319302 506504 319350 506560
rect 319406 506504 319411 506560
rect 319302 506502 319411 506504
rect 519862 506562 519922 506872
rect 522941 506562 523007 506565
rect 519862 506560 523007 506562
rect 519862 506504 522946 506560
rect 523002 506504 523007 506560
rect 519862 506502 523007 506504
rect 319345 506499 319411 506502
rect 522941 506499 523007 506502
rect 357433 506426 357499 506429
rect 401593 506426 401659 506429
rect 357433 506424 360210 506426
rect 357433 506368 357438 506424
rect 357494 506368 360210 506424
rect 357433 506366 360210 506368
rect 357433 506363 357499 506366
rect 360150 506192 360210 506366
rect 399894 506424 401659 506426
rect 399894 506368 401598 506424
rect 401654 506368 401659 506424
rect 399894 506366 401659 506368
rect 399894 506192 399954 506366
rect 401593 506363 401659 506366
rect 478321 506426 478387 506429
rect 478321 506424 480178 506426
rect 478321 506368 478326 506424
rect 478382 506368 480178 506424
rect 478321 506366 480178 506368
rect 478321 506363 478387 506366
rect 480118 506192 480178 506366
rect 254301 506154 254367 506157
rect 251804 506152 254367 506154
rect 251804 506096 254306 506152
rect 254362 506096 254367 506152
rect 251804 506094 254367 506096
rect 254301 506091 254367 506094
rect 320081 506086 320147 506089
rect 319884 506084 320147 506086
rect 319884 506028 320086 506084
rect 320142 506028 320147 506084
rect 319884 506026 320147 506028
rect 320081 506023 320147 506026
rect 399518 505956 399524 506020
rect 399588 505956 399594 506020
rect 357617 505882 357683 505885
rect 357617 505880 360210 505882
rect 357617 505824 357622 505880
rect 357678 505824 360210 505880
rect 357617 505822 360210 505824
rect 357617 505819 357683 505822
rect 360150 505512 360210 505822
rect 399526 505512 399586 505956
rect 519862 505746 519922 506192
rect 520733 505746 520799 505749
rect 519862 505744 520799 505746
rect 519862 505688 520738 505744
rect 520794 505688 520799 505744
rect 519862 505686 520799 505688
rect 520733 505683 520799 505686
rect 320265 505406 320331 505409
rect 319884 505404 320466 505406
rect 319884 505348 320270 505404
rect 320326 505348 320466 505404
rect 319884 505346 320466 505348
rect 320265 505343 320331 505346
rect 320406 505341 320466 505346
rect 320406 505336 320515 505341
rect 320406 505280 320454 505336
rect 320510 505280 320515 505336
rect 320406 505278 320515 505280
rect 320449 505275 320515 505278
rect 519862 505205 519922 505512
rect 519862 505200 519971 505205
rect 519862 505144 519910 505200
rect 519966 505144 519971 505200
rect 519862 505142 519971 505144
rect 519905 505139 519971 505142
rect 359038 505004 359044 505068
rect 359108 505066 359114 505068
rect 401225 505066 401291 505069
rect 359108 505006 360210 505066
rect 359108 505004 359114 505006
rect 360150 504832 360210 505006
rect 399894 505064 401291 505066
rect 399894 505008 401230 505064
rect 401286 505008 401291 505064
rect 399894 505006 401291 505008
rect 399894 504832 399954 505006
rect 401225 505003 401291 505006
rect 319854 504658 319914 504696
rect 321553 504658 321619 504661
rect 319854 504656 321619 504658
rect 319854 504600 321558 504656
rect 321614 504600 321619 504656
rect 319854 504598 321619 504600
rect 321553 504595 321619 504598
rect 357433 504658 357499 504661
rect 401777 504658 401843 504661
rect 357433 504656 360210 504658
rect 357433 504600 357438 504656
rect 357494 504600 360210 504656
rect 357433 504598 360210 504600
rect 357433 504595 357499 504598
rect 322473 504522 322539 504525
rect 319854 504520 322539 504522
rect 319854 504464 322478 504520
rect 322534 504464 322539 504520
rect 319854 504462 322539 504464
rect 319854 504016 319914 504462
rect 322473 504459 322539 504462
rect 360150 504152 360210 504598
rect 399894 504656 401843 504658
rect 399894 504600 401782 504656
rect 401838 504600 401843 504656
rect 399894 504598 401843 504600
rect 399894 504152 399954 504598
rect 401777 504595 401843 504598
rect 479149 504386 479215 504389
rect 480118 504386 480178 504832
rect 479149 504384 480178 504386
rect 479149 504328 479154 504384
rect 479210 504328 480178 504384
rect 479149 504326 480178 504328
rect 479149 504323 479215 504326
rect 478137 503842 478203 503845
rect 480118 503842 480178 504152
rect 478137 503840 480178 503842
rect 478137 503784 478142 503840
rect 478198 503784 480178 503840
rect 478137 503782 480178 503784
rect 519862 503842 519922 504152
rect 519997 503842 520063 503845
rect 519862 503840 520063 503842
rect 519862 503784 520002 503840
rect 520058 503784 520063 503840
rect 519862 503782 520063 503784
rect 478137 503779 478203 503782
rect 519997 503779 520063 503782
rect 358261 503706 358327 503709
rect 358261 503704 360210 503706
rect 358261 503648 358266 503704
rect 358322 503648 360210 503704
rect 358261 503646 360210 503648
rect 358261 503643 358327 503646
rect 322473 503570 322539 503573
rect 319854 503568 322539 503570
rect 319854 503512 322478 503568
rect 322534 503512 322539 503568
rect 319854 503510 322539 503512
rect 319854 503336 319914 503510
rect 322473 503507 322539 503510
rect 360150 503472 360210 503646
rect 356697 503298 356763 503301
rect 401593 503298 401659 503301
rect 356697 503296 360210 503298
rect 356697 503240 356702 503296
rect 356758 503240 360210 503296
rect 356697 503238 360210 503240
rect 356697 503235 356763 503238
rect 49601 503164 49667 503165
rect 49550 503162 49556 503164
rect 49474 503102 49556 503162
rect 49620 503162 49667 503164
rect 49620 503160 52164 503162
rect 49662 503104 52164 503160
rect 49550 503100 49556 503102
rect 49620 503102 52164 503104
rect 49620 503100 49667 503102
rect 49601 503099 49667 503100
rect 360150 502792 360210 503238
rect 399894 503296 401659 503298
rect 399894 503240 401598 503296
rect 401654 503240 401659 503296
rect 399894 503238 401659 503240
rect 399894 502792 399954 503238
rect 401593 503235 401659 503238
rect 477493 502890 477559 502893
rect 480118 502890 480178 503472
rect 519862 503026 519922 503472
rect 521694 503026 521700 503028
rect 519862 502966 521700 503026
rect 521694 502964 521700 502966
rect 521764 502964 521770 503028
rect 477493 502888 480178 502890
rect 477493 502832 477498 502888
rect 477554 502832 480178 502888
rect 477493 502830 480178 502832
rect 477493 502827 477559 502830
rect 319854 502482 319914 502656
rect 322473 502482 322539 502485
rect 319854 502480 322539 502482
rect 319854 502424 322478 502480
rect 322534 502424 322539 502480
rect 319854 502422 322539 502424
rect 519862 502482 519922 502792
rect 522389 502482 522455 502485
rect 519862 502480 522455 502482
rect 519862 502424 522394 502480
rect 522450 502424 522455 502480
rect 519862 502422 522455 502424
rect 322473 502419 322539 502422
rect 522389 502419 522455 502422
rect 358854 502284 358860 502348
rect 358924 502346 358930 502348
rect 358924 502286 360210 502346
rect 358924 502284 358930 502286
rect 360150 502112 360210 502286
rect 357433 501938 357499 501941
rect 357433 501936 360210 501938
rect -960 501802 480 501892
rect 357433 501880 357438 501936
rect 357494 501880 360210 501936
rect 357433 501878 360210 501880
rect 357433 501875 357499 501878
rect -960 501742 674 501802
rect -960 501666 480 501742
rect 614 501666 674 501742
rect -960 501652 674 501666
rect 246 501606 674 501652
rect 246 501122 306 501606
rect 360150 501432 360210 501878
rect 399526 501669 399586 502112
rect 399477 501664 399586 501669
rect 399477 501608 399482 501664
rect 399538 501608 399586 501664
rect 399477 501606 399586 501608
rect 477585 501666 477651 501669
rect 480118 501666 480178 502112
rect 477585 501664 480178 501666
rect 477585 501608 477590 501664
rect 477646 501608 480178 501664
rect 477585 501606 480178 501608
rect 399477 501603 399543 501606
rect 477585 501603 477651 501606
rect 400254 501462 400260 501464
rect 399924 501402 400260 501462
rect 400254 501400 400260 501402
rect 400324 501400 400330 501464
rect 477493 501258 477559 501261
rect 480118 501258 480178 501432
rect 477493 501256 480178 501258
rect 477493 501200 477498 501256
rect 477554 501200 480178 501256
rect 477493 501198 480178 501200
rect 477493 501195 477559 501198
rect 246 501062 6930 501122
rect 6870 500986 6930 501062
rect 49734 500986 49740 500988
rect 6870 500926 49740 500986
rect 49734 500924 49740 500926
rect 49804 500924 49810 500988
rect 519862 500986 519922 501432
rect 521837 500986 521903 500989
rect 519862 500984 521903 500986
rect 519862 500928 521842 500984
rect 521898 500928 521903 500984
rect 519862 500926 521903 500928
rect 521837 500923 521903 500926
rect 359733 500850 359799 500853
rect 522113 500850 522179 500853
rect 359733 500848 360210 500850
rect 359733 500792 359738 500848
rect 359794 500792 360210 500848
rect 359733 500790 360210 500792
rect 359733 500787 359799 500790
rect 360150 500752 360210 500790
rect 519862 500848 522179 500850
rect 519862 500792 522118 500848
rect 522174 500792 522179 500848
rect 519862 500790 522179 500792
rect 519862 500752 519922 500790
rect 522113 500787 522179 500790
rect 254577 500306 254643 500309
rect 251804 500304 254643 500306
rect 251804 500248 254582 500304
rect 254638 500248 254643 500304
rect 251804 500246 254643 500248
rect 399894 500306 399954 500752
rect 401593 500306 401659 500309
rect 399894 500304 401659 500306
rect 399894 500248 401598 500304
rect 401654 500248 401659 500304
rect 399894 500246 401659 500248
rect 254577 500243 254643 500246
rect 401593 500243 401659 500246
rect 477493 500170 477559 500173
rect 480118 500170 480178 500752
rect 519721 500578 519787 500581
rect 477493 500168 480178 500170
rect 477493 500112 477498 500168
rect 477554 500112 480178 500168
rect 477493 500110 480178 500112
rect 519678 500576 519787 500578
rect 519678 500520 519726 500576
rect 519782 500520 519787 500576
rect 519678 500515 519787 500520
rect 477493 500107 477559 500110
rect 519678 500072 519738 500515
rect 360653 499898 360719 499901
rect 362953 499900 363019 499901
rect 361430 499898 361436 499900
rect 360653 499896 361436 499898
rect 360653 499840 360658 499896
rect 360714 499840 361436 499896
rect 360653 499838 361436 499840
rect 360653 499835 360719 499838
rect 361430 499836 361436 499838
rect 361500 499836 361506 499900
rect 362902 499898 362908 499900
rect 362862 499838 362908 499898
rect 362972 499896 363019 499900
rect 363014 499840 363019 499896
rect 362902 499836 362908 499838
rect 362972 499836 363019 499840
rect 364742 499836 364748 499900
rect 364812 499898 364818 499900
rect 365161 499898 365227 499901
rect 364812 499896 365227 499898
rect 364812 499840 365166 499896
rect 365222 499840 365227 499896
rect 364812 499838 365227 499840
rect 364812 499836 364818 499838
rect 362953 499835 363019 499836
rect 365161 499835 365227 499838
rect 368238 499836 368244 499900
rect 368308 499898 368314 499900
rect 368381 499898 368447 499901
rect 368308 499896 368447 499898
rect 368308 499840 368386 499896
rect 368442 499840 368447 499896
rect 368308 499838 368447 499840
rect 368308 499836 368314 499838
rect 368381 499835 368447 499838
rect 369894 499836 369900 499900
rect 369964 499898 369970 499900
rect 370957 499898 371023 499901
rect 371601 499900 371667 499901
rect 369964 499896 371023 499898
rect 369964 499840 370962 499896
rect 371018 499840 371023 499896
rect 369964 499838 371023 499840
rect 369964 499836 369970 499838
rect 370957 499835 371023 499838
rect 371550 499836 371556 499900
rect 371620 499898 371667 499900
rect 371620 499896 371712 499898
rect 371662 499840 371712 499896
rect 371620 499838 371712 499840
rect 371620 499836 371667 499838
rect 376150 499836 376156 499900
rect 376220 499898 376226 499900
rect 376385 499898 376451 499901
rect 376220 499896 376451 499898
rect 376220 499840 376390 499896
rect 376446 499840 376451 499896
rect 376220 499838 376451 499840
rect 376220 499836 376226 499838
rect 371601 499835 371667 499836
rect 376385 499835 376451 499838
rect 376886 499836 376892 499900
rect 376956 499898 376962 499900
rect 377397 499898 377463 499901
rect 380617 499900 380683 499901
rect 376956 499896 377463 499898
rect 376956 499840 377402 499896
rect 377458 499840 377463 499896
rect 376956 499838 377463 499840
rect 376956 499836 376962 499838
rect 377397 499835 377463 499838
rect 380566 499836 380572 499900
rect 380636 499898 380683 499900
rect 380636 499896 380728 499898
rect 380678 499840 380728 499896
rect 380636 499838 380728 499840
rect 380636 499836 380683 499838
rect 380934 499836 380940 499900
rect 381004 499898 381010 499900
rect 381261 499898 381327 499901
rect 381004 499896 381327 499898
rect 381004 499840 381266 499896
rect 381322 499840 381327 499896
rect 381004 499838 381327 499840
rect 381004 499836 381010 499838
rect 380617 499835 380683 499836
rect 381261 499835 381327 499838
rect 382549 499898 382615 499901
rect 382774 499898 382780 499900
rect 382549 499896 382780 499898
rect 382549 499840 382554 499896
rect 382610 499840 382780 499896
rect 382549 499838 382780 499840
rect 382549 499835 382615 499838
rect 382774 499836 382780 499838
rect 382844 499836 382850 499900
rect 385534 499836 385540 499900
rect 385604 499898 385610 499900
rect 385769 499898 385835 499901
rect 385604 499896 385835 499898
rect 385604 499840 385774 499896
rect 385830 499840 385835 499896
rect 385604 499838 385835 499840
rect 385604 499836 385610 499838
rect 385769 499835 385835 499838
rect 386454 499836 386460 499900
rect 386524 499898 386530 499900
rect 387701 499898 387767 499901
rect 386524 499896 387767 499898
rect 386524 499840 387706 499896
rect 387762 499840 387767 499896
rect 386524 499838 387767 499840
rect 386524 499836 386530 499838
rect 387701 499835 387767 499838
rect 389582 499836 389588 499900
rect 389652 499898 389658 499900
rect 390277 499898 390343 499901
rect 389652 499896 390343 499898
rect 389652 499840 390282 499896
rect 390338 499840 390343 499896
rect 389652 499838 390343 499840
rect 389652 499836 389658 499838
rect 390277 499835 390343 499838
rect 391974 499836 391980 499900
rect 392044 499898 392050 499900
rect 392853 499898 392919 499901
rect 392044 499896 392919 499898
rect 392044 499840 392858 499896
rect 392914 499840 392919 499896
rect 392044 499838 392919 499840
rect 392044 499836 392050 499838
rect 392853 499835 392919 499838
rect 394734 499836 394740 499900
rect 394804 499898 394810 499900
rect 395429 499898 395495 499901
rect 394804 499896 395495 499898
rect 394804 499840 395434 499896
rect 395490 499840 395495 499896
rect 394804 499838 395495 499840
rect 394804 499836 394810 499838
rect 395429 499835 395495 499838
rect 398598 499836 398604 499900
rect 398668 499898 398674 499900
rect 399342 499898 399402 500072
rect 398668 499838 399402 499898
rect 502563 499898 502629 499901
rect 502926 499898 502932 499900
rect 502563 499896 502932 499898
rect 502563 499840 502568 499896
rect 502624 499840 502932 499896
rect 502563 499838 502932 499840
rect 398668 499836 398674 499838
rect 502563 499835 502629 499838
rect 502926 499836 502932 499838
rect 502996 499836 503002 499900
rect 360009 499762 360075 499765
rect 361614 499762 361620 499764
rect 360009 499760 361620 499762
rect 360009 499704 360014 499760
rect 360070 499704 361620 499760
rect 360009 499702 361620 499704
rect 360009 499699 360075 499702
rect 361614 499700 361620 499702
rect 361684 499700 361690 499764
rect 385125 499762 385191 499765
rect 385718 499762 385724 499764
rect 385125 499760 385724 499762
rect 385125 499704 385130 499760
rect 385186 499704 385724 499760
rect 385125 499702 385724 499704
rect 385125 499699 385191 499702
rect 385718 499700 385724 499702
rect 385788 499700 385794 499764
rect 495934 499564 495940 499628
rect 496004 499626 496010 499628
rect 496077 499626 496143 499629
rect 496004 499624 496143 499626
rect 496004 499568 496082 499624
rect 496138 499568 496143 499624
rect 496004 499566 496143 499568
rect 496004 499564 496010 499566
rect 496077 499563 496143 499566
rect 356605 499490 356671 499493
rect 365805 499490 365871 499493
rect 366214 499490 366220 499492
rect 356605 499488 366220 499490
rect 356605 499432 356610 499488
rect 356666 499432 365810 499488
rect 365866 499432 366220 499488
rect 356605 499430 366220 499432
rect 356605 499427 356671 499430
rect 365805 499427 365871 499430
rect 366214 499428 366220 499430
rect 366284 499428 366290 499492
rect 367737 499490 367803 499493
rect 368974 499490 368980 499492
rect 367737 499488 368980 499490
rect 367737 499432 367742 499488
rect 367798 499432 368980 499488
rect 367737 499430 368980 499432
rect 367737 499427 367803 499430
rect 368974 499428 368980 499430
rect 369044 499428 369050 499492
rect 376334 499428 376340 499492
rect 376404 499490 376410 499492
rect 376753 499490 376819 499493
rect 376404 499488 376819 499490
rect 376404 499432 376758 499488
rect 376814 499432 376819 499488
rect 376404 499430 376819 499432
rect 376404 499428 376410 499430
rect 376753 499427 376819 499430
rect 360694 499292 360700 499356
rect 360764 499354 360770 499356
rect 374821 499354 374887 499357
rect 360764 499352 374887 499354
rect 360764 499296 374826 499352
rect 374882 499296 374887 499352
rect 360764 499294 374887 499296
rect 360764 499292 360770 499294
rect 374821 499291 374887 499294
rect 298318 498748 298324 498812
rect 298388 498810 298394 498812
rect 477585 498810 477651 498813
rect 298388 498808 477651 498810
rect 298388 498752 477590 498808
rect 477646 498752 477651 498808
rect 298388 498750 477651 498752
rect 298388 498748 298394 498750
rect 477585 498747 477651 498750
rect 369025 498130 369091 498133
rect 373206 498130 373212 498132
rect 369025 498128 373212 498130
rect 369025 498072 369030 498128
rect 369086 498072 373212 498128
rect 369025 498070 373212 498072
rect 369025 498067 369091 498070
rect 373206 498068 373212 498070
rect 373276 498068 373282 498132
rect 376109 498130 376175 498133
rect 377254 498130 377260 498132
rect 376109 498128 377260 498130
rect 376109 498072 376114 498128
rect 376170 498072 377260 498128
rect 376109 498070 377260 498072
rect 376109 498067 376175 498070
rect 377254 498068 377260 498070
rect 377324 498068 377330 498132
rect 384062 498068 384068 498132
rect 384132 498130 384138 498132
rect 386413 498130 386479 498133
rect 384132 498128 386479 498130
rect 384132 498072 386418 498128
rect 386474 498072 386479 498128
rect 384132 498070 386479 498072
rect 384132 498068 384138 498070
rect 386413 498067 386479 498070
rect 378726 497932 378732 497996
rect 378796 497994 378802 497996
rect 387057 497994 387123 497997
rect 378796 497992 387123 497994
rect 378796 497936 387062 497992
rect 387118 497936 387123 497992
rect 378796 497934 387123 497936
rect 378796 497932 378802 497934
rect 387057 497931 387123 497934
rect 391054 497932 391060 497996
rect 391124 497994 391130 497996
rect 398649 497994 398715 497997
rect 391124 497992 398715 497994
rect 391124 497936 398654 497992
rect 398710 497936 398715 497992
rect 391124 497934 398715 497936
rect 391124 497932 391130 497934
rect 398649 497931 398715 497934
rect 359365 497858 359431 497861
rect 385769 497858 385835 497861
rect 359365 497856 385835 497858
rect 359365 497800 359370 497856
rect 359426 497800 385774 497856
rect 385830 497800 385835 497856
rect 583520 497844 584960 498084
rect 359365 497798 385835 497800
rect 359365 497795 359431 497798
rect 385769 497795 385835 497798
rect 360469 497722 360535 497725
rect 385125 497722 385191 497725
rect 360469 497720 385191 497722
rect 360469 497664 360474 497720
rect 360530 497664 385130 497720
rect 385186 497664 385191 497720
rect 360469 497662 385191 497664
rect 360469 497659 360535 497662
rect 385125 497659 385191 497662
rect 355225 497586 355291 497589
rect 391565 497586 391631 497589
rect 393998 497586 394004 497588
rect 355225 497584 394004 497586
rect 355225 497528 355230 497584
rect 355286 497528 391570 497584
rect 391626 497528 394004 497584
rect 355225 497526 394004 497528
rect 355225 497523 355291 497526
rect 391565 497523 391631 497526
rect 393998 497524 394004 497526
rect 394068 497524 394074 497588
rect 362585 497450 362651 497453
rect 382222 497450 382228 497452
rect 362585 497448 382228 497450
rect 362585 497392 362590 497448
rect 362646 497392 382228 497448
rect 362585 497390 382228 497392
rect 362585 497387 362651 497390
rect 382222 497388 382228 497390
rect 382292 497388 382298 497452
rect 48865 497314 48931 497317
rect 351269 497314 351335 497317
rect 369025 497314 369091 497317
rect 48865 497312 52164 497314
rect 48865 497256 48870 497312
rect 48926 497256 52164 497312
rect 48865 497254 52164 497256
rect 351269 497312 369091 497314
rect 351269 497256 351274 497312
rect 351330 497256 369030 497312
rect 369086 497256 369091 497312
rect 351269 497254 369091 497256
rect 48865 497251 48931 497254
rect 351269 497251 351335 497254
rect 369025 497251 369091 497254
rect 348509 497178 348575 497181
rect 382549 497178 382615 497181
rect 348509 497176 382615 497178
rect 348509 497120 348514 497176
rect 348570 497120 382554 497176
rect 382610 497120 382615 497176
rect 348509 497118 382615 497120
rect 348509 497115 348575 497118
rect 382549 497115 382615 497118
rect 349286 496844 349292 496908
rect 349356 496906 349362 496908
rect 350073 496906 350139 496909
rect 349356 496904 350139 496906
rect 349356 496848 350078 496904
rect 350134 496848 350139 496904
rect 349356 496846 350139 496848
rect 349356 496844 349362 496846
rect 350073 496843 350139 496846
rect 484342 496844 484348 496908
rect 484412 496906 484418 496908
rect 484485 496906 484551 496909
rect 485630 496906 485636 496908
rect 484412 496904 485636 496906
rect 484412 496848 484490 496904
rect 484546 496848 485636 496904
rect 484412 496846 485636 496848
rect 484412 496844 484418 496846
rect 484485 496843 484551 496846
rect 485630 496844 485636 496846
rect 485700 496844 485706 496908
rect 494697 496906 494763 496909
rect 496077 496906 496143 496909
rect 494697 496904 496143 496906
rect 494697 496848 494702 496904
rect 494758 496848 496082 496904
rect 496138 496848 496143 496904
rect 494697 496846 496143 496848
rect 494697 496843 494763 496846
rect 496077 496843 496143 496846
rect 254577 494458 254643 494461
rect 251804 494456 254643 494458
rect 251804 494400 254582 494456
rect 254638 494400 254643 494456
rect 251804 494398 254643 494400
rect 254577 494395 254643 494398
rect 49509 491466 49575 491469
rect 49509 491464 52164 491466
rect 49509 491408 49514 491464
rect 49570 491408 52164 491464
rect 49509 491406 52164 491408
rect 49509 491403 49575 491406
rect -960 488596 480 488836
rect 254577 488610 254643 488613
rect 251804 488608 254643 488610
rect 251804 488552 254582 488608
rect 254638 488552 254643 488608
rect 251804 488550 254643 488552
rect 254577 488547 254643 488550
rect 49601 485618 49667 485621
rect 51022 485618 51028 485620
rect 49601 485616 51028 485618
rect 49601 485560 49606 485616
rect 49662 485560 51028 485616
rect 49601 485558 51028 485560
rect 49601 485555 49667 485558
rect 51022 485556 51028 485558
rect 51092 485618 51098 485620
rect 51092 485558 52164 485618
rect 51092 485556 51098 485558
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 49601 484396 49667 484397
rect 49550 484332 49556 484396
rect 49620 484394 49667 484396
rect 49620 484392 49712 484394
rect 49662 484336 49712 484392
rect 49620 484334 49712 484336
rect 49620 484332 49667 484334
rect 49601 484331 49667 484332
rect 254577 482762 254643 482765
rect 251804 482760 254643 482762
rect 251804 482704 254582 482760
rect 254638 482704 254643 482760
rect 251804 482702 254643 482704
rect 254577 482699 254643 482702
rect 49366 479708 49372 479772
rect 49436 479770 49442 479772
rect 49436 479710 52164 479770
rect 49436 479708 49442 479710
rect 254209 476914 254275 476917
rect 251804 476912 254275 476914
rect 251804 476856 254214 476912
rect 254270 476856 254275 476912
rect 251804 476854 254275 476856
rect 254209 476851 254275 476854
rect -960 475540 480 475780
rect 48957 473922 49023 473925
rect 48957 473920 52164 473922
rect 48957 473864 48962 473920
rect 49018 473864 52164 473920
rect 48957 473862 52164 473864
rect 48957 473859 49023 473862
rect 580165 471474 580231 471477
rect 583520 471474 584960 471564
rect 580165 471472 584960 471474
rect 580165 471416 580170 471472
rect 580226 471416 584960 471472
rect 580165 471414 584960 471416
rect 580165 471411 580231 471414
rect 583520 471324 584960 471414
rect 254577 471066 254643 471069
rect 251804 471064 254643 471066
rect 251804 471008 254582 471064
rect 254638 471008 254643 471064
rect 251804 471006 254643 471008
rect 254577 471003 254643 471006
rect 48773 468074 48839 468077
rect 48773 468072 52164 468074
rect 48773 468016 48778 468072
rect 48834 468016 52164 468072
rect 48773 468014 52164 468016
rect 48773 468011 48839 468014
rect 254577 465218 254643 465221
rect 251804 465216 254643 465218
rect 251804 465160 254582 465216
rect 254638 465160 254643 465216
rect 251804 465158 254643 465160
rect 254577 465155 254643 465158
rect -960 462634 480 462724
rect 3509 462634 3575 462637
rect -960 462632 3575 462634
rect -960 462576 3514 462632
rect 3570 462576 3575 462632
rect -960 462574 3575 462576
rect -960 462484 480 462574
rect 3509 462571 3575 462574
rect 50797 462226 50863 462229
rect 50797 462224 52164 462226
rect 50797 462168 50802 462224
rect 50858 462168 52164 462224
rect 50797 462166 52164 462168
rect 50797 462163 50863 462166
rect 254577 459370 254643 459373
rect 251804 459368 254643 459370
rect 251804 459312 254582 459368
rect 254638 459312 254643 459368
rect 251804 459310 254643 459312
rect 254577 459307 254643 459310
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 49785 456378 49851 456381
rect 50705 456378 50771 456381
rect 49785 456376 52164 456378
rect 49785 456320 49790 456376
rect 49846 456320 50710 456376
rect 50766 456320 52164 456376
rect 49785 456318 52164 456320
rect 49785 456315 49851 456318
rect 50705 456315 50771 456318
rect 254301 453522 254367 453525
rect 251804 453520 254367 453522
rect 251804 453464 254306 453520
rect 254362 453464 254367 453520
rect 251804 453462 254367 453464
rect 254301 453459 254367 453462
rect 50613 450530 50679 450533
rect 51349 450530 51415 450533
rect 50613 450528 52164 450530
rect 50613 450472 50618 450528
rect 50674 450472 51354 450528
rect 51410 450472 52164 450528
rect 50613 450470 52164 450472
rect 50613 450467 50679 450470
rect 51349 450467 51415 450470
rect -960 449578 480 449668
rect 3417 449578 3483 449581
rect -960 449576 3483 449578
rect -960 449520 3422 449576
rect 3478 449520 3483 449576
rect -960 449518 3483 449520
rect -960 449428 480 449518
rect 3417 449515 3483 449518
rect 254669 447674 254735 447677
rect 251804 447672 254735 447674
rect 251804 447616 254674 447672
rect 254730 447616 254735 447672
rect 251804 447614 254735 447616
rect 254669 447611 254735 447614
rect 48313 444682 48379 444685
rect 48313 444680 52164 444682
rect 48313 444624 48318 444680
rect 48374 444624 52164 444680
rect 583520 444668 584960 444908
rect 48313 444622 52164 444624
rect 48313 444619 48379 444622
rect 254393 441826 254459 441829
rect 251804 441824 254459 441826
rect 251804 441768 254398 441824
rect 254454 441768 254459 441824
rect 251804 441766 254459 441768
rect 254393 441763 254459 441766
rect 48313 438834 48379 438837
rect 48313 438832 52164 438834
rect 48313 438776 48318 438832
rect 48374 438776 52164 438832
rect 48313 438774 52164 438776
rect 48313 438771 48379 438774
rect -960 436508 480 436748
rect 254393 435978 254459 435981
rect 251804 435976 254459 435978
rect 251804 435920 254398 435976
rect 254454 435920 254459 435976
rect 251804 435918 254459 435920
rect 254393 435915 254459 435918
rect 49141 432986 49207 432989
rect 49141 432984 52164 432986
rect 49141 432928 49146 432984
rect 49202 432928 52164 432984
rect 49141 432926 52164 432928
rect 49141 432923 49207 432926
rect 579797 431626 579863 431629
rect 583520 431626 584960 431716
rect 579797 431624 584960 431626
rect 579797 431568 579802 431624
rect 579858 431568 584960 431624
rect 579797 431566 584960 431568
rect 579797 431563 579863 431566
rect 583520 431476 584960 431566
rect 254577 430130 254643 430133
rect 251804 430128 254643 430130
rect 251804 430072 254582 430128
rect 254638 430072 254643 430128
rect 251804 430070 254643 430072
rect 254577 430067 254643 430070
rect 47945 427138 48011 427141
rect 47945 427136 52164 427138
rect 47945 427080 47950 427136
rect 48006 427080 52164 427136
rect 47945 427078 52164 427080
rect 47945 427075 48011 427078
rect 254577 424282 254643 424285
rect 251804 424280 254643 424282
rect 251804 424224 254582 424280
rect 254638 424224 254643 424280
rect 251804 424222 254643 424224
rect 254577 424219 254643 424222
rect -960 423452 480 423692
rect 48037 421290 48103 421293
rect 48037 421288 52164 421290
rect 48037 421232 48042 421288
rect 48098 421232 52164 421288
rect 48037 421230 52164 421232
rect 48037 421227 48103 421230
rect 254577 418434 254643 418437
rect 251804 418432 254643 418434
rect 251804 418376 254582 418432
rect 254638 418376 254643 418432
rect 251804 418374 254643 418376
rect 254577 418371 254643 418374
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 48129 415442 48195 415445
rect 48129 415440 52164 415442
rect 48129 415384 48134 415440
rect 48190 415384 52164 415440
rect 48129 415382 52164 415384
rect 48129 415379 48195 415382
rect 254577 412586 254643 412589
rect 251804 412584 254643 412586
rect 251804 412528 254582 412584
rect 254638 412528 254643 412584
rect 251804 412526 254643 412528
rect 254577 412523 254643 412526
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 48221 409594 48287 409597
rect 48221 409592 52164 409594
rect 48221 409536 48226 409592
rect 48282 409536 52164 409592
rect 48221 409534 52164 409536
rect 48221 409531 48287 409534
rect 254577 406738 254643 406741
rect 251804 406736 254643 406738
rect 251804 406680 254582 406736
rect 254638 406680 254643 406736
rect 251804 406678 254643 406680
rect 254577 406675 254643 406678
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 51441 403746 51507 403749
rect 51441 403744 52164 403746
rect 51441 403688 51446 403744
rect 51502 403688 52164 403744
rect 51441 403686 52164 403688
rect 51441 403683 51507 403686
rect 254025 400890 254091 400893
rect 251804 400888 254091 400890
rect 251804 400832 254030 400888
rect 254086 400832 254091 400888
rect 251804 400830 254091 400832
rect 254025 400827 254091 400830
rect 49417 397898 49483 397901
rect 49417 397896 52164 397898
rect 49417 397840 49422 397896
rect 49478 397840 52164 397896
rect 49417 397838 52164 397840
rect 49417 397835 49483 397838
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 254669 395042 254735 395045
rect 251804 395040 254735 395042
rect 251804 394984 254674 395040
rect 254730 394984 254735 395040
rect 251804 394982 254735 394984
rect 254669 394979 254735 394982
rect 48313 392050 48379 392053
rect 48313 392048 52164 392050
rect 48313 391992 48318 392048
rect 48374 391992 52164 392048
rect 48313 391990 52164 391992
rect 48313 391987 48379 391990
rect 583520 391628 584960 391868
rect 254669 389194 254735 389197
rect 251804 389192 254735 389194
rect 251804 389136 254674 389192
rect 254730 389136 254735 389192
rect 251804 389134 254735 389136
rect 254669 389131 254735 389134
rect 48313 386202 48379 386205
rect 48313 386200 52164 386202
rect 48313 386144 48318 386200
rect 48374 386144 52164 386200
rect 48313 386142 52164 386144
rect 48313 386139 48379 386142
rect -960 384284 480 384524
rect 254393 383346 254459 383349
rect 251804 383344 254459 383346
rect 251804 383288 254398 383344
rect 254454 383288 254459 383344
rect 251804 383286 254459 383288
rect 254393 383283 254459 383286
rect 49417 380354 49483 380357
rect 49417 380352 52164 380354
rect 49417 380296 49422 380352
rect 49478 380296 52164 380352
rect 49417 380294 52164 380296
rect 49417 380291 49483 380294
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 254117 377498 254183 377501
rect 251804 377496 254183 377498
rect 251804 377440 254122 377496
rect 254178 377440 254183 377496
rect 251804 377438 254183 377440
rect 254117 377435 254183 377438
rect 48221 374506 48287 374509
rect 48221 374504 52164 374506
rect 48221 374448 48226 374504
rect 48282 374448 52164 374504
rect 48221 374446 52164 374448
rect 48221 374443 48287 374446
rect 254669 371650 254735 371653
rect 251804 371648 254735 371650
rect 251804 371592 254674 371648
rect 254730 371592 254735 371648
rect 251804 371590 254735 371592
rect 254669 371587 254735 371590
rect -960 371228 480 371468
rect 48129 368658 48195 368661
rect 48129 368656 52164 368658
rect 48129 368600 48134 368656
rect 48190 368600 52164 368656
rect 48129 368598 52164 368600
rect 48129 368595 48195 368598
rect 254669 365802 254735 365805
rect 251804 365800 254735 365802
rect 251804 365744 254674 365800
rect 254730 365744 254735 365800
rect 251804 365742 254735 365744
rect 254669 365739 254735 365742
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 48037 362810 48103 362813
rect 48037 362808 52164 362810
rect 48037 362752 48042 362808
rect 48098 362752 52164 362808
rect 48037 362750 52164 362752
rect 48037 362747 48103 362750
rect 253933 359954 253999 359957
rect 251804 359952 253999 359954
rect 251804 359896 253938 359952
rect 253994 359896 253999 359952
rect 251804 359894 253999 359896
rect 253933 359891 253999 359894
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 51441 356962 51507 356965
rect 51441 356960 52164 356962
rect 51441 356904 51446 356960
rect 51502 356904 52164 356960
rect 51441 356902 52164 356904
rect 51441 356899 51507 356902
rect 254209 354106 254275 354109
rect 251804 354104 254275 354106
rect 251804 354048 254214 354104
rect 254270 354048 254275 354104
rect 251804 354046 254275 354048
rect 254209 354043 254275 354046
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 47945 351114 48011 351117
rect 47945 351112 52164 351114
rect 47945 351056 47950 351112
rect 48006 351056 52164 351112
rect 47945 351054 52164 351056
rect 47945 351051 48011 351054
rect 298502 349692 298508 349756
rect 298572 349754 298578 349756
rect 321645 349754 321711 349757
rect 298572 349752 321711 349754
rect 298572 349696 321650 349752
rect 321706 349696 321711 349752
rect 298572 349694 321711 349696
rect 298572 349692 298578 349694
rect 321645 349691 321711 349694
rect 254485 348258 254551 348261
rect 251804 348256 254551 348258
rect 251804 348200 254490 348256
rect 254546 348200 254551 348256
rect 251804 348198 254551 348200
rect 254485 348195 254551 348198
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 47853 345266 47919 345269
rect 47853 345264 52164 345266
rect 47853 345208 47858 345264
rect 47914 345208 52164 345264
rect 47853 345206 52164 345208
rect 47853 345203 47919 345206
rect 254577 342410 254643 342413
rect 251804 342408 254643 342410
rect 251804 342352 254582 342408
rect 254638 342352 254643 342408
rect 251804 342350 254643 342352
rect 254577 342347 254643 342350
rect 51533 339418 51599 339421
rect 51533 339416 52164 339418
rect 51533 339360 51538 339416
rect 51594 339360 52164 339416
rect 51533 339358 52164 339360
rect 51533 339355 51599 339358
rect 583520 338452 584960 338692
rect 254393 336562 254459 336565
rect 251804 336560 254459 336562
rect 251804 336504 254398 336560
rect 254454 336504 254459 336560
rect 251804 336502 254459 336504
rect 254393 336499 254459 336502
rect 299790 335956 299796 336020
rect 299860 336018 299866 336020
rect 322197 336018 322263 336021
rect 299860 336016 322263 336018
rect 299860 335960 322202 336016
rect 322258 335960 322263 336016
rect 299860 335958 322263 335960
rect 299860 335956 299866 335958
rect 322197 335955 322263 335958
rect 51717 333570 51783 333573
rect 51717 333568 52164 333570
rect 51717 333512 51722 333568
rect 51778 333512 52164 333568
rect 51717 333510 52164 333512
rect 51717 333507 51783 333510
rect -960 332196 480 332436
rect 254577 331530 254643 331533
rect 348969 331530 349035 331533
rect 254577 331528 349035 331530
rect 254577 331472 254582 331528
rect 254638 331472 348974 331528
rect 349030 331472 349035 331528
rect 254577 331470 349035 331472
rect 254577 331467 254643 331470
rect 348969 331467 349035 331470
rect 296069 331394 296135 331397
rect 316125 331394 316191 331397
rect 296069 331392 316191 331394
rect 296069 331336 296074 331392
rect 296130 331336 316130 331392
rect 316186 331336 316191 331392
rect 296069 331334 316191 331336
rect 296069 331331 296135 331334
rect 316125 331331 316191 331334
rect 299606 331196 299612 331260
rect 299676 331258 299682 331260
rect 305177 331258 305243 331261
rect 299676 331256 305243 331258
rect 299676 331200 305182 331256
rect 305238 331200 305243 331256
rect 299676 331198 305243 331200
rect 299676 331196 299682 331198
rect 305177 331195 305243 331198
rect 254209 330714 254275 330717
rect 251804 330712 254275 330714
rect 251804 330656 254214 330712
rect 254270 330656 254275 330712
rect 251804 330654 254275 330656
rect 254209 330651 254275 330654
rect 297357 329762 297423 329765
rect 297357 329760 300196 329762
rect 297357 329704 297362 329760
rect 297418 329704 300196 329760
rect 297357 329702 300196 329704
rect 297357 329699 297423 329702
rect 350257 329082 350323 329085
rect 349876 329080 350323 329082
rect 349876 329024 350262 329080
rect 350318 329024 350323 329080
rect 349876 329022 350323 329024
rect 350257 329019 350323 329022
rect 297449 328402 297515 328405
rect 297449 328400 300196 328402
rect 297449 328344 297454 328400
rect 297510 328344 300196 328400
rect 297449 328342 300196 328344
rect 297449 328339 297515 328342
rect 49417 327722 49483 327725
rect 350073 327722 350139 327725
rect 49417 327720 52164 327722
rect 49417 327664 49422 327720
rect 49478 327664 52164 327720
rect 49417 327662 52164 327664
rect 349876 327720 350139 327722
rect 349876 327664 350078 327720
rect 350134 327664 350139 327720
rect 349876 327662 350139 327664
rect 49417 327659 49483 327662
rect 350073 327659 350139 327662
rect 297541 326362 297607 326365
rect 351913 326362 351979 326365
rect 297541 326360 300196 326362
rect 297541 326304 297546 326360
rect 297602 326304 300196 326360
rect 297541 326302 300196 326304
rect 349876 326360 351979 326362
rect 349876 326304 351918 326360
rect 351974 326304 351979 326360
rect 349876 326302 351979 326304
rect 297541 326299 297607 326302
rect 351913 326299 351979 326302
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 297725 325002 297791 325005
rect 350993 325002 351059 325005
rect 297725 325000 300196 325002
rect 297725 324944 297730 325000
rect 297786 324944 300196 325000
rect 297725 324942 300196 324944
rect 349876 325000 351059 325002
rect 349876 324944 350998 325000
rect 351054 324944 351059 325000
rect 349876 324942 351059 324944
rect 297725 324939 297791 324942
rect 350993 324939 351059 324942
rect 254485 324866 254551 324869
rect 251804 324864 254551 324866
rect 251804 324808 254490 324864
rect 254546 324808 254551 324864
rect 251804 324806 254551 324808
rect 254485 324803 254551 324806
rect 297817 323642 297883 323645
rect 352373 323642 352439 323645
rect 297817 323640 300196 323642
rect 297817 323584 297822 323640
rect 297878 323584 300196 323640
rect 297817 323582 300196 323584
rect 349876 323640 352439 323642
rect 349876 323584 352378 323640
rect 352434 323584 352439 323640
rect 349876 323582 352439 323584
rect 297817 323579 297883 323582
rect 352373 323579 352439 323582
rect 299657 322282 299723 322285
rect 299657 322280 300196 322282
rect 299657 322224 299662 322280
rect 299718 322224 300196 322280
rect 299657 322222 300196 322224
rect 299657 322219 299723 322222
rect 49325 321874 49391 321877
rect 49325 321872 52164 321874
rect 49325 321816 49330 321872
rect 49386 321816 52164 321872
rect 49325 321814 52164 321816
rect 49325 321811 49391 321814
rect 351913 321602 351979 321605
rect 349876 321600 351979 321602
rect 349876 321544 351918 321600
rect 351974 321544 351979 321600
rect 349876 321542 351979 321544
rect 351913 321539 351979 321542
rect 297081 320242 297147 320245
rect 351862 320242 351868 320244
rect 297081 320240 300196 320242
rect 297081 320184 297086 320240
rect 297142 320184 300196 320240
rect 297081 320182 300196 320184
rect 349876 320182 351868 320242
rect 297081 320179 297147 320182
rect 351862 320180 351868 320182
rect 351932 320180 351938 320244
rect -960 319140 480 319380
rect 254301 319018 254367 319021
rect 251804 319016 254367 319018
rect 251804 318960 254306 319016
rect 254362 318960 254367 319016
rect 251804 318958 254367 318960
rect 254301 318955 254367 318958
rect 297173 318882 297239 318885
rect 352005 318882 352071 318885
rect 297173 318880 300196 318882
rect 297173 318824 297178 318880
rect 297234 318824 300196 318880
rect 297173 318822 300196 318824
rect 349876 318880 352071 318882
rect 349876 318824 352010 318880
rect 352066 318824 352071 318880
rect 349876 318822 352071 318824
rect 297173 318819 297239 318822
rect 352005 318819 352071 318822
rect 297725 317522 297791 317525
rect 351085 317522 351151 317525
rect 297725 317520 300196 317522
rect 297725 317464 297730 317520
rect 297786 317464 300196 317520
rect 297725 317462 300196 317464
rect 349876 317520 351151 317522
rect 349876 317464 351090 317520
rect 351146 317464 351151 317520
rect 349876 317462 351151 317464
rect 297725 317459 297791 317462
rect 351085 317459 351151 317462
rect 297725 316162 297791 316165
rect 297725 316160 300196 316162
rect 297725 316104 297730 316160
rect 297786 316104 300196 316160
rect 297725 316102 300196 316104
rect 297725 316099 297791 316102
rect 49233 316026 49299 316029
rect 349797 316026 349863 316029
rect 49233 316024 52164 316026
rect 49233 315968 49238 316024
rect 49294 315968 52164 316024
rect 49233 315966 52164 315968
rect 349797 316024 349906 316026
rect 349797 315968 349802 316024
rect 349858 315968 349906 316024
rect 49233 315963 49299 315966
rect 349797 315963 349906 315968
rect 349846 315452 349906 315963
rect 297909 314802 297975 314805
rect 297909 314800 300196 314802
rect 297909 314744 297914 314800
rect 297970 314744 300196 314800
rect 297909 314742 300196 314744
rect 297909 314739 297975 314742
rect 350901 314122 350967 314125
rect 349876 314120 350967 314122
rect 349876 314064 350906 314120
rect 350962 314064 350967 314120
rect 349876 314062 350967 314064
rect 350901 314059 350967 314062
rect 254669 313170 254735 313173
rect 251804 313168 254735 313170
rect 251804 313112 254674 313168
rect 254730 313112 254735 313168
rect 251804 313110 254735 313112
rect 254669 313107 254735 313110
rect 297909 312762 297975 312765
rect 297909 312760 300196 312762
rect 297909 312704 297914 312760
rect 297970 312704 300196 312760
rect 297909 312702 300196 312704
rect 297909 312699 297975 312702
rect 349846 312221 349906 312732
rect 349797 312216 349906 312221
rect 349797 312160 349802 312216
rect 349858 312160 349906 312216
rect 349797 312158 349906 312160
rect 349797 312155 349863 312158
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 298001 311402 298067 311405
rect 299381 311402 299447 311405
rect 298001 311400 300196 311402
rect 298001 311344 298006 311400
rect 298062 311344 299386 311400
rect 299442 311344 300196 311400
rect 298001 311342 300196 311344
rect 298001 311339 298067 311342
rect 299381 311339 299447 311342
rect 349846 310858 349906 311372
rect 350073 310858 350139 310861
rect 349846 310856 350139 310858
rect 349846 310800 350078 310856
rect 350134 310800 350139 310856
rect 349846 310798 350139 310800
rect 350073 310795 350139 310798
rect 51625 310178 51691 310181
rect 51625 310176 52164 310178
rect 51625 310120 51630 310176
rect 51686 310120 52164 310176
rect 51625 310118 52164 310120
rect 51625 310115 51691 310118
rect 297214 309980 297220 310044
rect 297284 310042 297290 310044
rect 352833 310042 352899 310045
rect 297284 309982 300196 310042
rect 349876 310040 352899 310042
rect 349876 309984 352838 310040
rect 352894 309984 352899 310040
rect 349876 309982 352899 309984
rect 297284 309980 297290 309982
rect 352833 309979 352899 309982
rect 298737 308682 298803 308685
rect 298737 308680 300196 308682
rect 298737 308624 298742 308680
rect 298798 308624 300196 308680
rect 298737 308622 300196 308624
rect 298737 308619 298803 308622
rect 351085 308002 351151 308005
rect 349876 308000 351151 308002
rect 349876 307944 351090 308000
rect 351146 307944 351151 308000
rect 349876 307942 351151 307944
rect 351085 307939 351151 307942
rect 254209 307322 254275 307325
rect 251804 307320 254275 307322
rect 251804 307264 254214 307320
rect 254270 307264 254275 307320
rect 251804 307262 254275 307264
rect 254209 307259 254275 307262
rect 297265 306642 297331 306645
rect 352557 306642 352623 306645
rect 297265 306640 300196 306642
rect 297265 306584 297270 306640
rect 297326 306584 300196 306640
rect 297265 306582 300196 306584
rect 349876 306640 352623 306642
rect 349876 306584 352562 306640
rect 352618 306584 352623 306640
rect 349876 306582 352623 306584
rect 297265 306579 297331 306582
rect 352557 306579 352623 306582
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 298001 305282 298067 305285
rect 351453 305282 351519 305285
rect 298001 305280 300196 305282
rect 298001 305224 298006 305280
rect 298062 305224 300196 305280
rect 298001 305222 300196 305224
rect 349876 305280 351519 305282
rect 349876 305224 351458 305280
rect 351514 305224 351519 305280
rect 349876 305222 351519 305224
rect 298001 305219 298067 305222
rect 351453 305219 351519 305222
rect 49141 304330 49207 304333
rect 49141 304328 52164 304330
rect 49141 304272 49146 304328
rect 49202 304272 52164 304328
rect 49141 304270 52164 304272
rect 49141 304267 49207 304270
rect 296989 303922 297055 303925
rect 350349 303922 350415 303925
rect 296989 303920 300196 303922
rect 296989 303864 296994 303920
rect 297050 303864 300196 303920
rect 296989 303862 300196 303864
rect 349876 303920 350415 303922
rect 349876 303864 350354 303920
rect 350410 303864 350415 303920
rect 349876 303862 350415 303864
rect 296989 303859 297055 303862
rect 350349 303859 350415 303862
rect 298001 302562 298067 302565
rect 298001 302560 300196 302562
rect 298001 302504 298006 302560
rect 298062 302504 300196 302560
rect 298001 302502 300196 302504
rect 298001 302499 298067 302502
rect 351913 301882 351979 301885
rect 349876 301880 351979 301882
rect 349876 301824 351918 301880
rect 351974 301824 351979 301880
rect 349876 301822 351979 301824
rect 351913 301819 351979 301822
rect 254669 301474 254735 301477
rect 251804 301472 254735 301474
rect 251804 301416 254674 301472
rect 254730 301416 254735 301472
rect 251804 301414 254735 301416
rect 254669 301411 254735 301414
rect 296989 301202 297055 301205
rect 296989 301200 300196 301202
rect 296989 301144 296994 301200
rect 297050 301144 300196 301200
rect 296989 301142 300196 301144
rect 296989 301139 297055 301142
rect 351913 300522 351979 300525
rect 349876 300520 351979 300522
rect 349876 300464 351918 300520
rect 351974 300464 351979 300520
rect 349876 300462 351979 300464
rect 351913 300459 351979 300462
rect 297909 299162 297975 299165
rect 351361 299162 351427 299165
rect 297909 299160 300196 299162
rect 297909 299104 297914 299160
rect 297970 299104 300196 299160
rect 297909 299102 300196 299104
rect 349876 299160 351427 299162
rect 349876 299104 351366 299160
rect 351422 299104 351427 299160
rect 349876 299102 351427 299104
rect 297909 299099 297975 299102
rect 351361 299099 351427 299102
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 48681 298482 48747 298485
rect 48681 298480 52164 298482
rect 48681 298424 48686 298480
rect 48742 298424 52164 298480
rect 48681 298422 52164 298424
rect 48681 298419 48747 298422
rect 299565 297802 299631 297805
rect 352097 297802 352163 297805
rect 299565 297800 300196 297802
rect 299565 297744 299570 297800
rect 299626 297744 300196 297800
rect 299565 297742 300196 297744
rect 349876 297800 352163 297802
rect 349876 297744 352102 297800
rect 352158 297744 352163 297800
rect 349876 297742 352163 297744
rect 299565 297739 299631 297742
rect 352097 297739 352163 297742
rect 297725 296442 297791 296445
rect 352281 296442 352347 296445
rect 297725 296440 300196 296442
rect 297725 296384 297730 296440
rect 297786 296384 300196 296440
rect 297725 296382 300196 296384
rect 349876 296440 352347 296442
rect 349876 296384 352286 296440
rect 352342 296384 352347 296440
rect 349876 296382 352347 296384
rect 297725 296379 297791 296382
rect 352281 296379 352347 296382
rect 254669 295626 254735 295629
rect 251804 295624 254735 295626
rect 251804 295568 254674 295624
rect 254730 295568 254735 295624
rect 251804 295566 254735 295568
rect 254669 295563 254735 295566
rect 297817 295082 297883 295085
rect 297817 295080 300196 295082
rect 297817 295024 297822 295080
rect 297878 295024 300196 295080
rect 297817 295022 300196 295024
rect 297817 295019 297883 295022
rect 352005 294402 352071 294405
rect 349876 294400 352071 294402
rect 349876 294344 352010 294400
rect 352066 294344 352071 294400
rect 349876 294342 352071 294344
rect 352005 294339 352071 294342
rect -960 293178 480 293268
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 352281 293042 352347 293045
rect 349876 293040 352347 293042
rect 48773 292634 48839 292637
rect 48773 292632 52164 292634
rect 48773 292576 48778 292632
rect 48834 292576 52164 292632
rect 48773 292574 52164 292576
rect 48773 292571 48839 292574
rect 284886 292572 284892 292636
rect 284956 292634 284962 292636
rect 300166 292634 300226 293012
rect 349876 292984 352286 293040
rect 352342 292984 352347 293040
rect 349876 292982 352347 292984
rect 352281 292979 352347 292982
rect 284956 292574 300226 292634
rect 284956 292572 284962 292574
rect 298001 291682 298067 291685
rect 350901 291682 350967 291685
rect 351361 291682 351427 291685
rect 298001 291680 300196 291682
rect 298001 291624 298006 291680
rect 298062 291624 300196 291680
rect 298001 291622 300196 291624
rect 349876 291680 351427 291682
rect 349876 291624 350906 291680
rect 350962 291624 351366 291680
rect 351422 291624 351427 291680
rect 349876 291622 351427 291624
rect 298001 291619 298067 291622
rect 350901 291619 350967 291622
rect 351361 291619 351427 291622
rect 349797 290866 349863 290869
rect 349797 290864 349906 290866
rect 349797 290808 349802 290864
rect 349858 290808 349906 290864
rect 349797 290803 349906 290808
rect 297909 290322 297975 290325
rect 297909 290320 300196 290322
rect 297909 290264 297914 290320
rect 297970 290264 300196 290320
rect 349846 290292 349906 290803
rect 297909 290262 300196 290264
rect 297909 290259 297975 290262
rect 254393 289778 254459 289781
rect 251804 289776 254459 289778
rect 251804 289720 254398 289776
rect 254454 289720 254459 289776
rect 251804 289718 254459 289720
rect 254393 289715 254459 289718
rect 298001 288962 298067 288965
rect 298001 288960 300196 288962
rect 298001 288904 298006 288960
rect 298062 288904 300196 288960
rect 298001 288902 300196 288904
rect 298001 288899 298067 288902
rect 351269 288282 351335 288285
rect 349876 288280 351335 288282
rect 349876 288224 351274 288280
rect 351330 288224 351335 288280
rect 349876 288222 351335 288224
rect 351269 288219 351335 288222
rect 298001 287602 298067 287605
rect 298001 287600 300196 287602
rect 298001 287544 298006 287600
rect 298062 287544 300196 287600
rect 298001 287542 300196 287544
rect 298001 287539 298067 287542
rect 51950 286726 52164 286786
rect 51950 286514 52010 286726
rect 52085 286514 52151 286517
rect 51950 286512 52151 286514
rect 51950 286456 52090 286512
rect 52146 286456 52151 286512
rect 51950 286454 52151 286456
rect 52085 286451 52151 286454
rect 349846 286381 349906 286892
rect 349797 286376 349906 286381
rect 349797 286320 349802 286376
rect 349858 286320 349906 286376
rect 349797 286318 349906 286320
rect 349797 286315 349863 286318
rect 297909 285562 297975 285565
rect 352097 285562 352163 285565
rect 297909 285560 300196 285562
rect 297909 285504 297914 285560
rect 297970 285504 300196 285560
rect 297909 285502 300196 285504
rect 349876 285560 352163 285562
rect 349876 285504 352102 285560
rect 352158 285504 352163 285560
rect 349876 285502 352163 285504
rect 297909 285499 297975 285502
rect 352097 285499 352163 285502
rect 583520 285276 584960 285516
rect 297633 284202 297699 284205
rect 352465 284202 352531 284205
rect 297633 284200 300196 284202
rect 297633 284144 297638 284200
rect 297694 284144 300196 284200
rect 297633 284142 300196 284144
rect 349876 284200 352531 284202
rect 349876 284144 352470 284200
rect 352526 284144 352531 284200
rect 349876 284142 352531 284144
rect 297633 284139 297699 284142
rect 352465 284139 352531 284142
rect 254301 283930 254367 283933
rect 251804 283928 254367 283930
rect 251804 283872 254306 283928
rect 254362 283872 254367 283928
rect 251804 283870 254367 283872
rect 254301 283867 254367 283870
rect 299565 282842 299631 282845
rect 352189 282842 352255 282845
rect 299565 282840 300196 282842
rect 299565 282784 299570 282840
rect 299626 282784 300196 282840
rect 299565 282782 300196 282784
rect 349876 282840 352255 282842
rect 349876 282784 352194 282840
rect 352250 282784 352255 282840
rect 349876 282782 352255 282784
rect 299565 282779 299631 282782
rect 352189 282779 352255 282782
rect 298093 282434 298159 282437
rect 298318 282434 298324 282436
rect 298093 282432 298324 282434
rect 298093 282376 298098 282432
rect 298154 282376 298324 282432
rect 298093 282374 298324 282376
rect 298093 282371 298159 282374
rect 298318 282372 298324 282374
rect 298388 282372 298394 282436
rect 51441 282026 51507 282029
rect 291142 282026 291148 282028
rect 51441 282024 291148 282026
rect 51441 281968 51446 282024
rect 51502 281968 291148 282024
rect 51441 281966 291148 281968
rect 51441 281963 51507 281966
rect 291142 281964 291148 281966
rect 291212 281964 291218 282028
rect 51625 281890 51691 281893
rect 285990 281890 285996 281892
rect 51625 281888 285996 281890
rect 51625 281832 51630 281888
rect 51686 281832 285996 281888
rect 51625 281830 285996 281832
rect 51625 281827 51691 281830
rect 285990 281828 285996 281830
rect 286060 281828 286066 281892
rect 282177 281482 282243 281485
rect 288566 281482 288572 281484
rect 282177 281480 288572 281482
rect 282177 281424 282182 281480
rect 282238 281424 288572 281480
rect 282177 281422 288572 281424
rect 282177 281419 282243 281422
rect 288566 281420 288572 281422
rect 288636 281420 288642 281484
rect 298645 281482 298711 281485
rect 485773 281482 485839 281485
rect 486366 281482 486372 281484
rect 298645 281480 300196 281482
rect 298645 281424 298650 281480
rect 298706 281424 300196 281480
rect 298645 281422 300196 281424
rect 485773 281480 486372 281482
rect 485773 281424 485778 281480
rect 485834 281424 486372 281480
rect 485773 281422 486372 281424
rect 298645 281419 298711 281422
rect 485773 281419 485839 281422
rect 486366 281420 486372 281422
rect 486436 281420 486442 281484
rect 47853 281346 47919 281349
rect 290774 281346 290780 281348
rect 47853 281344 290780 281346
rect 47853 281288 47858 281344
rect 47914 281288 290780 281344
rect 47853 281286 290780 281288
rect 47853 281283 47919 281286
rect 290774 281284 290780 281286
rect 290844 281284 290850 281348
rect 47945 281210 48011 281213
rect 290590 281210 290596 281212
rect 47945 281208 290596 281210
rect 47945 281152 47950 281208
rect 48006 281152 290596 281208
rect 47945 281150 290596 281152
rect 47945 281147 48011 281150
rect 290590 281148 290596 281150
rect 290660 281148 290666 281212
rect 49417 281074 49483 281077
rect 287278 281074 287284 281076
rect 49417 281072 287284 281074
rect 49417 281016 49422 281072
rect 49478 281016 287284 281072
rect 49417 281014 287284 281016
rect 49417 281011 49483 281014
rect 287278 281012 287284 281014
rect 287348 281012 287354 281076
rect 51533 280938 51599 280941
rect 282177 280938 282243 280941
rect 288382 280938 288388 280940
rect 51533 280936 282243 280938
rect 51533 280880 51538 280936
rect 51594 280880 282182 280936
rect 282238 280880 282243 280936
rect 51533 280878 282243 280880
rect 51533 280875 51599 280878
rect 282177 280875 282243 280878
rect 287010 280878 288388 280938
rect 51717 280802 51783 280805
rect 287010 280802 287070 280878
rect 288382 280876 288388 280878
rect 288452 280876 288458 280940
rect 51717 280800 287070 280802
rect 51717 280744 51722 280800
rect 51778 280744 287070 280800
rect 51717 280742 287070 280744
rect 287329 280802 287395 280805
rect 287646 280802 287652 280804
rect 287329 280800 287652 280802
rect 287329 280744 287334 280800
rect 287390 280744 287652 280800
rect 287329 280742 287652 280744
rect 51717 280739 51783 280742
rect 287329 280739 287395 280742
rect 287646 280740 287652 280742
rect 287716 280740 287722 280804
rect 350809 280802 350875 280805
rect 349876 280800 350875 280802
rect 349876 280744 350814 280800
rect 350870 280744 350875 280800
rect 349876 280742 350875 280744
rect 350809 280739 350875 280742
rect 46841 280666 46907 280669
rect 282126 280666 282132 280668
rect 46841 280664 282132 280666
rect 46841 280608 46846 280664
rect 46902 280608 282132 280664
rect 46841 280606 282132 280608
rect 46841 280603 46907 280606
rect 282126 280604 282132 280606
rect 282196 280604 282202 280668
rect 48129 280530 48195 280533
rect 292614 280530 292620 280532
rect 48129 280528 292620 280530
rect 48129 280472 48134 280528
rect 48190 280472 292620 280528
rect 48129 280470 292620 280472
rect 48129 280467 48195 280470
rect 292614 280468 292620 280470
rect 292684 280468 292690 280532
rect -960 279972 480 280212
rect 46749 280122 46815 280125
rect 295374 280122 295380 280124
rect 46749 280120 295380 280122
rect 46749 280064 46754 280120
rect 46810 280064 295380 280120
rect 46749 280062 295380 280064
rect 46749 280059 46815 280062
rect 295374 280060 295380 280062
rect 295444 280060 295450 280124
rect 46565 279986 46631 279989
rect 293902 279986 293908 279988
rect 46565 279984 293908 279986
rect 46565 279928 46570 279984
rect 46626 279928 293908 279984
rect 46565 279926 293908 279928
rect 46565 279923 46631 279926
rect 293902 279924 293908 279926
rect 293972 279924 293978 279988
rect 59353 279442 59419 279445
rect 297214 279442 297220 279444
rect 59353 279440 297220 279442
rect 59353 279384 59358 279440
rect 59414 279384 297220 279440
rect 59353 279382 297220 279384
rect 59353 279379 59419 279382
rect 297214 279380 297220 279382
rect 297284 279380 297290 279444
rect 49366 278700 49372 278764
rect 49436 278762 49442 278764
rect 54569 278762 54635 278765
rect 49436 278760 54635 278762
rect 49436 278704 54574 278760
rect 54630 278704 54635 278760
rect 49436 278702 54635 278704
rect 49436 278700 49442 278702
rect 54569 278699 54635 278702
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267052 480 267292
rect 583520 258906 584960 258996
rect 583342 258846 584960 258906
rect 583342 258770 583402 258846
rect 583520 258770 584960 258846
rect 583342 258756 584960 258770
rect 583342 258710 583586 258756
rect 355358 258028 355364 258092
rect 355428 258028 355434 258092
rect 355366 257954 355426 258028
rect 583526 257954 583586 258710
rect 355366 257894 583586 257954
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 57830 227020 57836 227084
rect 57900 227082 57906 227084
rect 257613 227082 257679 227085
rect 57900 227080 257679 227082
rect 57900 227024 257618 227080
rect 257674 227024 257679 227080
rect 57900 227022 257679 227024
rect 57900 227020 57906 227022
rect 257613 227019 257679 227022
rect 42793 226946 42859 226949
rect 522062 226946 522068 226948
rect 42793 226944 522068 226946
rect 42793 226888 42798 226944
rect 42854 226888 522068 226944
rect 42793 226886 522068 226888
rect 42793 226883 42859 226886
rect 522062 226884 522068 226886
rect 522132 226884 522138 226948
rect 59721 225586 59787 225589
rect 351862 225586 351868 225588
rect 59721 225584 351868 225586
rect 59721 225528 59726 225584
rect 59782 225528 351868 225584
rect 59721 225526 351868 225528
rect 59721 225523 59787 225526
rect 351862 225524 351868 225526
rect 351932 225524 351938 225588
rect 48957 224362 49023 224365
rect 521878 224362 521884 224364
rect 48957 224360 521884 224362
rect 48957 224304 48962 224360
rect 49018 224304 521884 224360
rect 48957 224302 521884 224304
rect 48957 224299 49023 224302
rect 521878 224300 521884 224302
rect 521948 224300 521954 224364
rect 3509 224226 3575 224229
rect 519118 224226 519124 224228
rect 3509 224224 519124 224226
rect 3509 224168 3514 224224
rect 3570 224168 519124 224224
rect 3509 224166 519124 224168
rect 3509 224163 3575 224166
rect 519118 224164 519124 224166
rect 519188 224164 519194 224228
rect 49550 223484 49556 223548
rect 49620 223546 49626 223548
rect 55857 223546 55923 223549
rect 49620 223544 55923 223546
rect 49620 223488 55862 223544
rect 55918 223488 55923 223544
rect 49620 223486 55923 223488
rect 49620 223484 49626 223486
rect 55857 223483 55923 223486
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 351126 218044 351132 218108
rect 351196 218106 351202 218108
rect 583526 218106 583586 218862
rect 351196 218046 583586 218106
rect 351196 218044 351202 218046
rect 297909 217698 297975 217701
rect 297909 217696 300196 217698
rect 297909 217640 297914 217696
rect 297970 217640 300196 217696
rect 297909 217638 300196 217640
rect 297909 217635 297975 217638
rect 57053 217426 57119 217429
rect 57053 217424 60076 217426
rect 57053 217368 57058 217424
rect 57114 217368 60076 217424
rect 57053 217366 60076 217368
rect 57053 217363 57119 217366
rect 297541 216746 297607 216749
rect 299606 216746 299612 216748
rect 297541 216744 299612 216746
rect 297541 216688 297546 216744
rect 297602 216688 299612 216744
rect 297541 216686 299612 216688
rect 297541 216683 297607 216686
rect 299606 216684 299612 216686
rect 299676 216684 299682 216748
rect 297909 216202 297975 216205
rect 297909 216200 300196 216202
rect 297909 216144 297914 216200
rect 297970 216144 300196 216200
rect 297909 216142 300196 216144
rect 297909 216139 297975 216142
rect 222837 215658 222903 215661
rect 219788 215656 222903 215658
rect 219788 215600 222842 215656
rect 222898 215600 222903 215656
rect 219788 215598 222903 215600
rect 222837 215595 222903 215598
rect -960 214828 480 215068
rect 297909 214706 297975 214709
rect 297909 214704 300196 214706
rect 297909 214648 297914 214704
rect 297970 214648 300196 214704
rect 297909 214646 300196 214648
rect 297909 214643 297975 214646
rect 60549 213890 60615 213893
rect 60549 213888 60658 213890
rect 60549 213832 60554 213888
rect 60610 213832 60658 213888
rect 60549 213827 60658 213832
rect 60598 213316 60658 213827
rect 297909 213210 297975 213213
rect 297909 213208 300196 213210
rect 297909 213152 297914 213208
rect 297970 213152 300196 213208
rect 297909 213150 300196 213152
rect 297909 213147 297975 213150
rect 222285 212802 222351 212805
rect 219788 212800 222351 212802
rect 219788 212744 222290 212800
rect 222346 212744 222351 212800
rect 219788 212742 222351 212744
rect 222285 212739 222351 212742
rect 297909 211714 297975 211717
rect 297909 211712 300196 211714
rect 297909 211656 297914 211712
rect 297970 211656 300196 211712
rect 297909 211654 300196 211656
rect 297909 211651 297975 211654
rect 297909 210218 297975 210221
rect 297909 210216 300196 210218
rect 297909 210160 297914 210216
rect 297970 210160 300196 210216
rect 297909 210158 300196 210160
rect 297909 210155 297975 210158
rect 223205 209946 223271 209949
rect 219788 209944 223271 209946
rect 219788 209888 223210 209944
rect 223266 209888 223271 209944
rect 219788 209886 223271 209888
rect 223205 209883 223271 209886
rect 57145 209266 57211 209269
rect 57145 209264 60076 209266
rect 57145 209208 57150 209264
rect 57206 209208 60076 209264
rect 57145 209206 60076 209208
rect 57145 209203 57211 209206
rect 296805 208722 296871 208725
rect 296805 208720 300196 208722
rect 296805 208664 296810 208720
rect 296866 208664 300196 208720
rect 296805 208662 300196 208664
rect 296805 208659 296871 208662
rect 297909 207226 297975 207229
rect 297909 207224 300196 207226
rect 297909 207168 297914 207224
rect 297970 207168 300196 207224
rect 297909 207166 300196 207168
rect 297909 207163 297975 207166
rect 222929 207090 222995 207093
rect 219788 207088 222995 207090
rect 219788 207032 222934 207088
rect 222990 207032 222995 207088
rect 219788 207030 222995 207032
rect 222929 207027 222995 207030
rect 296805 205730 296871 205733
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 296805 205728 300196 205730
rect 296805 205672 296810 205728
rect 296866 205672 300196 205728
rect 296805 205670 300196 205672
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 296805 205667 296871 205670
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 57329 205186 57395 205189
rect 57329 205184 60076 205186
rect 57329 205128 57334 205184
rect 57390 205128 60076 205184
rect 57329 205126 60076 205128
rect 57329 205123 57395 205126
rect 222837 204234 222903 204237
rect 219788 204232 222903 204234
rect 219788 204176 222842 204232
rect 222898 204176 222903 204232
rect 219788 204174 222903 204176
rect 222837 204171 222903 204174
rect 297909 204234 297975 204237
rect 297909 204232 300196 204234
rect 297909 204176 297914 204232
rect 297970 204176 300196 204232
rect 297909 204174 300196 204176
rect 297909 204171 297975 204174
rect 297909 202738 297975 202741
rect 297909 202736 300196 202738
rect 297909 202680 297914 202736
rect 297970 202680 300196 202736
rect 297909 202678 300196 202680
rect 297909 202675 297975 202678
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 223021 201378 223087 201381
rect 219788 201376 223087 201378
rect 219788 201320 223026 201376
rect 223082 201320 223087 201376
rect 219788 201318 223087 201320
rect 223021 201315 223087 201318
rect 297909 201242 297975 201245
rect 297909 201240 300196 201242
rect 297909 201184 297914 201240
rect 297970 201184 300196 201240
rect 297909 201182 300196 201184
rect 297909 201179 297975 201182
rect 57329 201106 57395 201109
rect 57329 201104 60076 201106
rect 57329 201048 57334 201104
rect 57390 201048 60076 201104
rect 57329 201046 60076 201048
rect 57329 201043 57395 201046
rect 297909 199746 297975 199749
rect 297909 199744 300196 199746
rect 297909 199688 297914 199744
rect 297970 199688 300196 199744
rect 297909 199686 300196 199688
rect 297909 199683 297975 199686
rect 222929 198522 222995 198525
rect 219788 198520 222995 198522
rect 219788 198464 222934 198520
rect 222990 198464 222995 198520
rect 219788 198462 222995 198464
rect 222929 198459 222995 198462
rect 297909 198250 297975 198253
rect 297909 198248 300196 198250
rect 297909 198192 297914 198248
rect 297970 198192 300196 198248
rect 297909 198190 300196 198192
rect 297909 198187 297975 198190
rect 57329 197026 57395 197029
rect 57329 197024 60076 197026
rect 57329 196968 57334 197024
rect 57390 196968 60076 197024
rect 57329 196966 60076 196968
rect 57329 196963 57395 196966
rect 297909 196754 297975 196757
rect 297909 196752 300196 196754
rect 297909 196696 297914 196752
rect 297970 196696 300196 196752
rect 297909 196694 300196 196696
rect 297909 196691 297975 196694
rect 223481 195666 223547 195669
rect 219788 195664 223547 195666
rect 219788 195608 223486 195664
rect 223542 195608 223547 195664
rect 219788 195606 223547 195608
rect 223481 195603 223547 195606
rect 297909 195258 297975 195261
rect 297909 195256 300196 195258
rect 297909 195200 297914 195256
rect 297970 195200 300196 195256
rect 297909 195198 300196 195200
rect 297909 195195 297975 195198
rect 297909 193762 297975 193765
rect 297909 193760 300196 193762
rect 297909 193704 297914 193760
rect 297970 193704 300196 193760
rect 297909 193702 300196 193704
rect 297909 193699 297975 193702
rect 57329 192946 57395 192949
rect 57329 192944 60076 192946
rect 57329 192888 57334 192944
rect 57390 192888 60076 192944
rect 57329 192886 60076 192888
rect 57329 192883 57395 192886
rect 223481 192810 223547 192813
rect 219788 192808 223547 192810
rect 219788 192752 223486 192808
rect 223542 192752 223547 192808
rect 219788 192750 223547 192752
rect 223481 192747 223547 192750
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 297725 192266 297791 192269
rect 297725 192264 300196 192266
rect 297725 192208 297730 192264
rect 297786 192208 300196 192264
rect 297725 192206 300196 192208
rect 297725 192203 297791 192206
rect 297909 190770 297975 190773
rect 297909 190768 300196 190770
rect 297909 190712 297914 190768
rect 297970 190712 300196 190768
rect 297909 190710 300196 190712
rect 297909 190707 297975 190710
rect 223481 189954 223547 189957
rect 219788 189952 223547 189954
rect 219788 189896 223486 189952
rect 223542 189896 223547 189952
rect 219788 189894 223547 189896
rect 223481 189891 223547 189894
rect 297725 189274 297791 189277
rect 297725 189272 300196 189274
rect 297725 189216 297730 189272
rect 297786 189216 300196 189272
rect 297725 189214 300196 189216
rect 297725 189211 297791 189214
rect -960 188866 480 188956
rect 3785 188866 3851 188869
rect -960 188864 3851 188866
rect -960 188808 3790 188864
rect 3846 188808 3851 188864
rect -960 188806 3851 188808
rect -960 188716 480 188806
rect 3785 188803 3851 188806
rect 57329 188866 57395 188869
rect 57329 188864 60076 188866
rect 57329 188808 57334 188864
rect 57390 188808 60076 188864
rect 57329 188806 60076 188808
rect 57329 188803 57395 188806
rect 297909 187778 297975 187781
rect 297909 187776 300196 187778
rect 297909 187720 297914 187776
rect 297970 187720 300196 187776
rect 297909 187718 300196 187720
rect 297909 187715 297975 187718
rect 223481 187098 223547 187101
rect 219788 187096 223547 187098
rect 219788 187040 223486 187096
rect 223542 187040 223547 187096
rect 219788 187038 223547 187040
rect 223481 187035 223547 187038
rect 296805 186282 296871 186285
rect 296805 186280 300196 186282
rect 296805 186224 296810 186280
rect 296866 186224 300196 186280
rect 296805 186222 300196 186224
rect 296805 186219 296871 186222
rect 56685 184786 56751 184789
rect 297909 184786 297975 184789
rect 56685 184784 60076 184786
rect 56685 184728 56690 184784
rect 56746 184728 60076 184784
rect 56685 184726 60076 184728
rect 297909 184784 300196 184786
rect 297909 184728 297914 184784
rect 297970 184728 300196 184784
rect 297909 184726 300196 184728
rect 56685 184723 56751 184726
rect 297909 184723 297975 184726
rect 222285 184242 222351 184245
rect 219788 184240 222351 184242
rect 219788 184184 222290 184240
rect 222346 184184 222351 184240
rect 219788 184182 222351 184184
rect 222285 184179 222351 184182
rect 297909 183290 297975 183293
rect 297909 183288 300196 183290
rect 297909 183232 297914 183288
rect 297970 183232 300196 183288
rect 297909 183230 300196 183232
rect 297909 183227 297975 183230
rect 297909 181794 297975 181797
rect 297909 181792 300196 181794
rect 297909 181736 297914 181792
rect 297970 181736 300196 181792
rect 297909 181734 300196 181736
rect 297909 181731 297975 181734
rect 223481 181386 223547 181389
rect 219788 181384 223547 181386
rect 219788 181328 223486 181384
rect 223542 181328 223547 181384
rect 219788 181326 223547 181328
rect 223481 181323 223547 181326
rect 56685 180706 56751 180709
rect 56685 180704 60076 180706
rect 56685 180648 56690 180704
rect 56746 180648 60076 180704
rect 56685 180646 60076 180648
rect 56685 180643 56751 180646
rect 295977 180298 296043 180301
rect 295977 180296 300196 180298
rect 295977 180240 295982 180296
rect 296038 180240 300196 180296
rect 295977 180238 300196 180240
rect 295977 180235 296043 180238
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 297909 178802 297975 178805
rect 297909 178800 300196 178802
rect 297909 178744 297914 178800
rect 297970 178744 300196 178800
rect 297909 178742 300196 178744
rect 297909 178739 297975 178742
rect 222653 178530 222719 178533
rect 219788 178528 222719 178530
rect 219788 178472 222658 178528
rect 222714 178472 222719 178528
rect 219788 178470 222719 178472
rect 222653 178467 222719 178470
rect 297909 177306 297975 177309
rect 297909 177304 300196 177306
rect 297909 177248 297914 177304
rect 297970 177248 300196 177304
rect 297909 177246 300196 177248
rect 297909 177243 297975 177246
rect 57329 176626 57395 176629
rect 57329 176624 60076 176626
rect 57329 176568 57334 176624
rect 57390 176568 60076 176624
rect 57329 176566 60076 176568
rect 57329 176563 57395 176566
rect -960 175796 480 176036
rect 297909 175810 297975 175813
rect 297909 175808 300196 175810
rect 297909 175752 297914 175808
rect 297970 175752 300196 175808
rect 297909 175750 300196 175752
rect 297909 175747 297975 175750
rect 222653 175674 222719 175677
rect 219788 175672 222719 175674
rect 219788 175616 222658 175672
rect 222714 175616 222719 175672
rect 219788 175614 222719 175616
rect 222653 175611 222719 175614
rect 297909 174314 297975 174317
rect 297909 174312 300196 174314
rect 297909 174256 297914 174312
rect 297970 174256 300196 174312
rect 297909 174254 300196 174256
rect 297909 174251 297975 174254
rect 222377 172818 222443 172821
rect 219788 172816 222443 172818
rect 219788 172760 222382 172816
rect 222438 172760 222443 172816
rect 219788 172758 222443 172760
rect 222377 172755 222443 172758
rect 297909 172818 297975 172821
rect 297909 172816 300196 172818
rect 297909 172760 297914 172816
rect 297970 172760 300196 172816
rect 297909 172758 300196 172760
rect 297909 172755 297975 172758
rect 57237 172546 57303 172549
rect 57237 172544 60076 172546
rect 57237 172488 57242 172544
rect 57298 172488 60076 172544
rect 57237 172486 60076 172488
rect 57237 172483 57303 172486
rect 297909 171322 297975 171325
rect 297909 171320 300196 171322
rect 297909 171264 297914 171320
rect 297970 171264 300196 171320
rect 297909 171262 300196 171264
rect 297909 171259 297975 171262
rect 222469 169962 222535 169965
rect 219788 169960 222535 169962
rect 219788 169904 222474 169960
rect 222530 169904 222535 169960
rect 219788 169902 222535 169904
rect 222469 169899 222535 169902
rect 296805 169826 296871 169829
rect 296805 169824 300196 169826
rect 296805 169768 296810 169824
rect 296866 169768 300196 169824
rect 296805 169766 300196 169768
rect 296805 169763 296871 169766
rect 57329 168466 57395 168469
rect 57329 168464 60076 168466
rect 57329 168408 57334 168464
rect 57390 168408 60076 168464
rect 57329 168406 60076 168408
rect 57329 168403 57395 168406
rect 297909 168330 297975 168333
rect 297909 168328 300196 168330
rect 297909 168272 297914 168328
rect 297970 168272 300196 168328
rect 297909 168270 300196 168272
rect 297909 168267 297975 168270
rect 222929 167106 222995 167109
rect 219788 167104 222995 167106
rect 219788 167048 222934 167104
rect 222990 167048 222995 167104
rect 219788 167046 222995 167048
rect 222929 167043 222995 167046
rect 297909 166834 297975 166837
rect 297909 166832 300196 166834
rect 297909 166776 297914 166832
rect 297970 166776 300196 166832
rect 297909 166774 300196 166776
rect 297909 166771 297975 166774
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 297909 165338 297975 165341
rect 297909 165336 300196 165338
rect 297909 165280 297914 165336
rect 297970 165280 300196 165336
rect 297909 165278 300196 165280
rect 297909 165275 297975 165278
rect 55857 164386 55923 164389
rect 55857 164384 60076 164386
rect 55857 164328 55862 164384
rect 55918 164328 60076 164384
rect 55857 164326 60076 164328
rect 55857 164323 55923 164326
rect 223481 164250 223547 164253
rect 219788 164248 223547 164250
rect 219788 164192 223486 164248
rect 223542 164192 223547 164248
rect 219788 164190 223547 164192
rect 223481 164187 223547 164190
rect 297909 163842 297975 163845
rect 297909 163840 300196 163842
rect 297909 163784 297914 163840
rect 297970 163784 300196 163840
rect 297909 163782 300196 163784
rect 297909 163779 297975 163782
rect -960 162740 480 162980
rect 297909 162346 297975 162349
rect 297909 162344 300196 162346
rect 297909 162288 297914 162344
rect 297970 162288 300196 162344
rect 297909 162286 300196 162288
rect 297909 162283 297975 162286
rect 223021 161394 223087 161397
rect 219788 161392 223087 161394
rect 219788 161336 223026 161392
rect 223082 161336 223087 161392
rect 219788 161334 223087 161336
rect 223021 161331 223087 161334
rect 295977 160850 296043 160853
rect 295977 160848 300196 160850
rect 295977 160792 295982 160848
rect 296038 160792 300196 160848
rect 295977 160790 300196 160792
rect 295977 160787 296043 160790
rect 57053 160306 57119 160309
rect 57053 160304 60076 160306
rect 57053 160248 57058 160304
rect 57114 160248 60076 160304
rect 57053 160246 60076 160248
rect 57053 160243 57119 160246
rect 297909 159354 297975 159357
rect 297909 159352 300196 159354
rect 297909 159296 297914 159352
rect 297970 159296 300196 159352
rect 297909 159294 300196 159296
rect 297909 159291 297975 159294
rect 222929 158538 222995 158541
rect 219788 158536 222995 158538
rect 219788 158480 222934 158536
rect 222990 158480 222995 158536
rect 219788 158478 222995 158480
rect 222929 158475 222995 158478
rect 297909 157858 297975 157861
rect 297909 157856 300196 157858
rect 297909 157800 297914 157856
rect 297970 157800 300196 157856
rect 297909 157798 300196 157800
rect 297909 157795 297975 157798
rect 297909 156362 297975 156365
rect 297909 156360 300196 156362
rect 297909 156304 297914 156360
rect 297970 156304 300196 156360
rect 297909 156302 300196 156304
rect 297909 156299 297975 156302
rect 57053 156226 57119 156229
rect 57053 156224 60076 156226
rect 57053 156168 57058 156224
rect 57114 156168 60076 156224
rect 57053 156166 60076 156168
rect 57053 156163 57119 156166
rect 223481 155682 223547 155685
rect 219788 155680 223547 155682
rect 219788 155624 223486 155680
rect 223542 155624 223547 155680
rect 219788 155622 223547 155624
rect 223481 155619 223547 155622
rect 297909 154866 297975 154869
rect 297909 154864 300196 154866
rect 297909 154808 297914 154864
rect 297970 154808 300196 154864
rect 297909 154806 300196 154808
rect 297909 154803 297975 154806
rect 297909 153370 297975 153373
rect 297909 153368 300196 153370
rect 297909 153312 297914 153368
rect 297970 153312 300196 153368
rect 297909 153310 300196 153312
rect 297909 153307 297975 153310
rect 222653 152826 222719 152829
rect 219788 152824 222719 152826
rect 219788 152768 222658 152824
rect 222714 152768 222719 152824
rect 219788 152766 222719 152768
rect 222653 152763 222719 152766
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 57329 152146 57395 152149
rect 57329 152144 60076 152146
rect 57329 152088 57334 152144
rect 57390 152088 60076 152144
rect 57329 152086 60076 152088
rect 57329 152083 57395 152086
rect 296805 151874 296871 151877
rect 296805 151872 300196 151874
rect 296805 151816 296810 151872
rect 296866 151816 300196 151872
rect 296805 151814 300196 151816
rect 296805 151811 296871 151814
rect 297909 150378 297975 150381
rect 297909 150376 300196 150378
rect 297909 150320 297914 150376
rect 297970 150320 300196 150376
rect 297909 150318 300196 150320
rect 297909 150315 297975 150318
rect 223205 149970 223271 149973
rect 219788 149968 223271 149970
rect -960 149834 480 149924
rect 219788 149912 223210 149968
rect 223266 149912 223271 149968
rect 219788 149910 223271 149912
rect 223205 149907 223271 149910
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 296069 148882 296135 148885
rect 296069 148880 300196 148882
rect 296069 148824 296074 148880
rect 296130 148824 300196 148880
rect 296069 148822 300196 148824
rect 296069 148819 296135 148822
rect 57329 148066 57395 148069
rect 57329 148064 60076 148066
rect 57329 148008 57334 148064
rect 57390 148008 60076 148064
rect 57329 148006 60076 148008
rect 57329 148003 57395 148006
rect 341057 147522 341123 147525
rect 339940 147520 341123 147522
rect 339940 147464 341062 147520
rect 341118 147464 341123 147520
rect 339940 147462 341123 147464
rect 341057 147459 341123 147462
rect 297909 147386 297975 147389
rect 297909 147384 300196 147386
rect 297909 147328 297914 147384
rect 297970 147328 300196 147384
rect 297909 147326 300196 147328
rect 297909 147323 297975 147326
rect 222561 147114 222627 147117
rect 219788 147112 222627 147114
rect 219788 147056 222566 147112
rect 222622 147056 222627 147112
rect 219788 147054 222627 147056
rect 222561 147051 222627 147054
rect 297909 145890 297975 145893
rect 297909 145888 300196 145890
rect 297909 145832 297914 145888
rect 297970 145832 300196 145888
rect 297909 145830 300196 145832
rect 297909 145827 297975 145830
rect 340137 145346 340203 145349
rect 339940 145344 340203 145346
rect 339940 145288 340142 145344
rect 340198 145288 340203 145344
rect 339940 145286 340203 145288
rect 340137 145283 340203 145286
rect 297909 144394 297975 144397
rect 297909 144392 300196 144394
rect 297909 144336 297914 144392
rect 297970 144336 300196 144392
rect 297909 144334 300196 144336
rect 297909 144331 297975 144334
rect 223481 144258 223547 144261
rect 219788 144256 223547 144258
rect 219788 144200 223486 144256
rect 223542 144200 223547 144256
rect 219788 144198 223547 144200
rect 223481 144195 223547 144198
rect 57329 143986 57395 143989
rect 57329 143984 60076 143986
rect 57329 143928 57334 143984
rect 57390 143928 60076 143984
rect 57329 143926 60076 143928
rect 57329 143923 57395 143926
rect 343081 143170 343147 143173
rect 339940 143168 343147 143170
rect 339940 143112 343086 143168
rect 343142 143112 343147 143168
rect 339940 143110 343147 143112
rect 343081 143107 343147 143110
rect 295977 142898 296043 142901
rect 295977 142896 300196 142898
rect 295977 142840 295982 142896
rect 296038 142840 300196 142896
rect 295977 142838 300196 142840
rect 295977 142835 296043 142838
rect 223481 141402 223547 141405
rect 219788 141400 223547 141402
rect 219788 141344 223486 141400
rect 223542 141344 223547 141400
rect 219788 141342 223547 141344
rect 223481 141339 223547 141342
rect 297909 141402 297975 141405
rect 297909 141400 300196 141402
rect 297909 141344 297914 141400
rect 297970 141344 300196 141400
rect 297909 141342 300196 141344
rect 297909 141339 297975 141342
rect 340873 140994 340939 140997
rect 339940 140992 340939 140994
rect 339940 140936 340878 140992
rect 340934 140936 340939 140992
rect 339940 140934 340939 140936
rect 340873 140931 340939 140934
rect 57421 139906 57487 139909
rect 297909 139906 297975 139909
rect 57421 139904 60076 139906
rect 57421 139848 57426 139904
rect 57482 139848 60076 139904
rect 57421 139846 60076 139848
rect 297909 139904 300196 139906
rect 297909 139848 297914 139904
rect 297970 139848 300196 139904
rect 297909 139846 300196 139848
rect 57421 139843 57487 139846
rect 297909 139843 297975 139846
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 340229 138818 340295 138821
rect 339940 138816 340295 138818
rect 339940 138760 340234 138816
rect 340290 138760 340295 138816
rect 339940 138758 340295 138760
rect 340229 138755 340295 138758
rect 222929 138546 222995 138549
rect 219788 138544 222995 138546
rect 219788 138488 222934 138544
rect 222990 138488 222995 138544
rect 219788 138486 222995 138488
rect 222929 138483 222995 138486
rect 297909 138410 297975 138413
rect 297909 138408 300196 138410
rect 297909 138352 297914 138408
rect 297970 138352 300196 138408
rect 297909 138350 300196 138352
rect 297909 138347 297975 138350
rect 297909 136914 297975 136917
rect 297909 136912 300196 136914
rect -960 136778 480 136868
rect 297909 136856 297914 136912
rect 297970 136856 300196 136912
rect 297909 136854 300196 136856
rect 297909 136851 297975 136854
rect 3601 136778 3667 136781
rect -960 136776 3667 136778
rect -960 136720 3606 136776
rect 3662 136720 3667 136776
rect -960 136718 3667 136720
rect -960 136628 480 136718
rect 3601 136715 3667 136718
rect 342437 136642 342503 136645
rect 339940 136640 342503 136642
rect 339940 136584 342442 136640
rect 342498 136584 342503 136640
rect 339940 136582 342503 136584
rect 342437 136579 342503 136582
rect 57329 135826 57395 135829
rect 57329 135824 60076 135826
rect 57329 135768 57334 135824
rect 57390 135768 60076 135824
rect 57329 135766 60076 135768
rect 57329 135763 57395 135766
rect 222837 135690 222903 135693
rect 219788 135688 222903 135690
rect 219788 135632 222842 135688
rect 222898 135632 222903 135688
rect 219788 135630 222903 135632
rect 222837 135627 222903 135630
rect 297909 135418 297975 135421
rect 297909 135416 300196 135418
rect 297909 135360 297914 135416
rect 297970 135360 300196 135416
rect 297909 135358 300196 135360
rect 297909 135355 297975 135358
rect 342253 134466 342319 134469
rect 339940 134464 342319 134466
rect 339940 134408 342258 134464
rect 342314 134408 342319 134464
rect 339940 134406 342319 134408
rect 342253 134403 342319 134406
rect 297909 133922 297975 133925
rect 297909 133920 300196 133922
rect 297909 133864 297914 133920
rect 297970 133864 300196 133920
rect 297909 133862 300196 133864
rect 297909 133859 297975 133862
rect 222653 132834 222719 132837
rect 219788 132832 222719 132834
rect 219788 132776 222658 132832
rect 222714 132776 222719 132832
rect 219788 132774 222719 132776
rect 222653 132771 222719 132774
rect 296805 132426 296871 132429
rect 296805 132424 300196 132426
rect 296805 132368 296810 132424
rect 296866 132368 300196 132424
rect 296805 132366 300196 132368
rect 296805 132363 296871 132366
rect 341149 132290 341215 132293
rect 339940 132288 341215 132290
rect 339940 132232 341154 132288
rect 341210 132232 341215 132288
rect 339940 132230 341215 132232
rect 341149 132227 341215 132230
rect 57830 131684 57836 131748
rect 57900 131746 57906 131748
rect 57900 131686 60076 131746
rect 57900 131684 57906 131686
rect 297909 130930 297975 130933
rect 297909 130928 300196 130930
rect 297909 130872 297914 130928
rect 297970 130872 300196 130928
rect 297909 130870 300196 130872
rect 297909 130867 297975 130870
rect 339940 130054 340154 130114
rect 340094 129981 340154 130054
rect 223021 129978 223087 129981
rect 219788 129976 223087 129978
rect 219788 129920 223026 129976
rect 223082 129920 223087 129976
rect 219788 129918 223087 129920
rect 223021 129915 223087 129918
rect 340045 129976 340154 129981
rect 340045 129920 340050 129976
rect 340106 129920 340154 129976
rect 340045 129918 340154 129920
rect 340045 129915 340111 129918
rect 296805 129434 296871 129437
rect 296805 129432 300196 129434
rect 296805 129376 296810 129432
rect 296866 129376 300196 129432
rect 296805 129374 300196 129376
rect 296805 129371 296871 129374
rect 297909 127938 297975 127941
rect 342529 127938 342595 127941
rect 297909 127936 300196 127938
rect 297909 127880 297914 127936
rect 297970 127880 300196 127936
rect 297909 127878 300196 127880
rect 339940 127936 342595 127938
rect 339940 127880 342534 127936
rect 342590 127880 342595 127936
rect 339940 127878 342595 127880
rect 297909 127875 297975 127878
rect 342529 127875 342595 127878
rect 58893 127666 58959 127669
rect 58893 127664 60076 127666
rect 58893 127608 58898 127664
rect 58954 127608 60076 127664
rect 58893 127606 60076 127608
rect 58893 127603 58959 127606
rect 222837 127122 222903 127125
rect 219788 127120 222903 127122
rect 219788 127064 222842 127120
rect 222898 127064 222903 127120
rect 219788 127062 222903 127064
rect 222837 127059 222903 127062
rect 297909 126442 297975 126445
rect 297909 126440 300196 126442
rect 297909 126384 297914 126440
rect 297970 126384 300196 126440
rect 297909 126382 300196 126384
rect 297909 126379 297975 126382
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 342621 125762 342687 125765
rect 339940 125760 342687 125762
rect 339940 125704 342626 125760
rect 342682 125704 342687 125760
rect 339940 125702 342687 125704
rect 342621 125699 342687 125702
rect 297909 124946 297975 124949
rect 297909 124944 300196 124946
rect 297909 124888 297914 124944
rect 297970 124888 300196 124944
rect 297909 124886 300196 124888
rect 297909 124883 297975 124886
rect 222285 124266 222351 124269
rect 219788 124264 222351 124266
rect 219788 124208 222290 124264
rect 222346 124208 222351 124264
rect 219788 124206 222351 124208
rect 222285 124203 222351 124206
rect -960 123572 480 123812
rect 57513 123586 57579 123589
rect 342713 123586 342779 123589
rect 57513 123584 60076 123586
rect 57513 123528 57518 123584
rect 57574 123528 60076 123584
rect 57513 123526 60076 123528
rect 339940 123584 342779 123586
rect 339940 123528 342718 123584
rect 342774 123528 342779 123584
rect 339940 123526 342779 123528
rect 57513 123523 57579 123526
rect 342713 123523 342779 123526
rect 297909 123450 297975 123453
rect 297909 123448 300196 123450
rect 297909 123392 297914 123448
rect 297970 123392 300196 123448
rect 297909 123390 300196 123392
rect 297909 123387 297975 123390
rect 297909 121954 297975 121957
rect 297909 121952 300196 121954
rect 297909 121896 297914 121952
rect 297970 121896 300196 121952
rect 297909 121894 300196 121896
rect 297909 121891 297975 121894
rect 223481 121410 223547 121413
rect 340965 121410 341031 121413
rect 219788 121408 223547 121410
rect 219788 121352 223486 121408
rect 223542 121352 223547 121408
rect 219788 121350 223547 121352
rect 339940 121408 341031 121410
rect 339940 121352 340970 121408
rect 341026 121352 341031 121408
rect 339940 121350 341031 121352
rect 223481 121347 223547 121350
rect 340965 121347 341031 121350
rect 297909 120458 297975 120461
rect 297909 120456 300196 120458
rect 297909 120400 297914 120456
rect 297970 120400 300196 120456
rect 297909 120398 300196 120400
rect 297909 120395 297975 120398
rect 58801 119506 58867 119509
rect 58801 119504 60076 119506
rect 58801 119448 58806 119504
rect 58862 119448 60076 119504
rect 58801 119446 60076 119448
rect 58801 119443 58867 119446
rect 340321 119234 340387 119237
rect 339940 119232 340387 119234
rect 339940 119176 340326 119232
rect 340382 119176 340387 119232
rect 339940 119174 340387 119176
rect 340321 119171 340387 119174
rect 297909 118962 297975 118965
rect 297909 118960 300196 118962
rect 297909 118904 297914 118960
rect 297970 118904 300196 118960
rect 297909 118902 300196 118904
rect 297909 118899 297975 118902
rect 223481 118554 223547 118557
rect 219788 118552 223547 118554
rect 219788 118496 223486 118552
rect 223542 118496 223547 118552
rect 219788 118494 223547 118496
rect 223481 118491 223547 118494
rect 297909 117466 297975 117469
rect 297909 117464 300196 117466
rect 297909 117408 297914 117464
rect 297970 117408 300196 117464
rect 297909 117406 300196 117408
rect 297909 117403 297975 117406
rect 342345 117058 342411 117061
rect 339940 117056 342411 117058
rect 339940 117000 342350 117056
rect 342406 117000 342411 117056
rect 339940 116998 342411 117000
rect 342345 116995 342411 116998
rect 297909 115970 297975 115973
rect 297909 115968 300196 115970
rect 297909 115912 297914 115968
rect 297970 115912 300196 115968
rect 297909 115910 300196 115912
rect 297909 115907 297975 115910
rect 223481 115698 223547 115701
rect 219788 115696 223547 115698
rect 219788 115640 223486 115696
rect 223542 115640 223547 115696
rect 219788 115638 223547 115640
rect 223481 115635 223547 115638
rect 59445 115426 59511 115429
rect 59445 115424 60076 115426
rect 59445 115368 59450 115424
rect 59506 115368 60076 115424
rect 59445 115366 60076 115368
rect 59445 115363 59511 115366
rect 341333 114882 341399 114885
rect 339940 114880 341399 114882
rect 339940 114824 341338 114880
rect 341394 114824 341399 114880
rect 339940 114822 341399 114824
rect 341333 114819 341399 114822
rect 296805 114474 296871 114477
rect 296805 114472 300196 114474
rect 296805 114416 296810 114472
rect 296866 114416 300196 114472
rect 296805 114414 300196 114416
rect 296805 114411 296871 114414
rect 297909 112978 297975 112981
rect 297909 112976 300196 112978
rect 297909 112920 297914 112976
rect 297970 112920 300196 112976
rect 297909 112918 300196 112920
rect 297909 112915 297975 112918
rect 222193 112842 222259 112845
rect 219788 112840 222259 112842
rect 219788 112784 222198 112840
rect 222254 112784 222259 112840
rect 219788 112782 222259 112784
rect 222193 112779 222259 112782
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 341241 112706 341307 112709
rect 339940 112704 341307 112706
rect 339940 112648 341246 112704
rect 341302 112648 341307 112704
rect 583520 112692 584960 112782
rect 339940 112646 341307 112648
rect 341241 112643 341307 112646
rect 298921 111482 298987 111485
rect 298921 111480 300196 111482
rect 298921 111424 298926 111480
rect 298982 111424 300196 111480
rect 298921 111422 300196 111424
rect 298921 111419 298987 111422
rect 58709 111346 58775 111349
rect 58709 111344 60076 111346
rect 58709 111288 58714 111344
rect 58770 111288 60076 111344
rect 58709 111286 60076 111288
rect 58709 111283 58775 111286
rect -960 110516 480 110756
rect 340413 110530 340479 110533
rect 339940 110528 340479 110530
rect 339940 110472 340418 110528
rect 340474 110472 340479 110528
rect 339940 110470 340479 110472
rect 340413 110467 340479 110470
rect 223481 109986 223547 109989
rect 219788 109984 223547 109986
rect 219788 109928 223486 109984
rect 223542 109928 223547 109984
rect 219788 109926 223547 109928
rect 223481 109923 223547 109926
rect 297357 109986 297423 109989
rect 297357 109984 300196 109986
rect 297357 109928 297362 109984
rect 297418 109928 300196 109984
rect 297357 109926 300196 109928
rect 297357 109923 297423 109926
rect 299013 108490 299079 108493
rect 299013 108488 300196 108490
rect 299013 108432 299018 108488
rect 299074 108432 300196 108488
rect 299013 108430 300196 108432
rect 299013 108427 299079 108430
rect 340822 108354 340828 108356
rect 339940 108294 340828 108354
rect 340822 108292 340828 108294
rect 340892 108354 340898 108356
rect 342345 108354 342411 108357
rect 340892 108352 342411 108354
rect 340892 108296 342350 108352
rect 342406 108296 342411 108352
rect 340892 108294 342411 108296
rect 340892 108292 340898 108294
rect 342345 108291 342411 108294
rect 57605 107266 57671 107269
rect 57605 107264 60076 107266
rect 57605 107208 57610 107264
rect 57666 107208 60076 107264
rect 57605 107206 60076 107208
rect 57605 107203 57671 107206
rect 222653 107130 222719 107133
rect 219788 107128 222719 107130
rect 219788 107072 222658 107128
rect 222714 107072 222719 107128
rect 219788 107070 222719 107072
rect 222653 107067 222719 107070
rect 299105 106994 299171 106997
rect 299105 106992 300196 106994
rect 299105 106936 299110 106992
rect 299166 106936 300196 106992
rect 299105 106934 300196 106936
rect 299105 106931 299171 106934
rect 342345 106180 342411 106181
rect 342294 106178 342300 106180
rect 339940 106118 342300 106178
rect 342364 106176 342411 106180
rect 342406 106120 342411 106176
rect 342294 106116 342300 106118
rect 342364 106116 342411 106120
rect 342345 106115 342411 106116
rect 299197 105498 299263 105501
rect 299197 105496 300196 105498
rect 299197 105440 299202 105496
rect 299258 105440 300196 105496
rect 299197 105438 300196 105440
rect 299197 105435 299263 105438
rect 222837 104274 222903 104277
rect 219788 104272 222903 104274
rect 219788 104216 222842 104272
rect 222898 104216 222903 104272
rect 219788 104214 222903 104216
rect 222837 104211 222903 104214
rect 297449 104002 297515 104005
rect 341425 104002 341491 104005
rect 297449 104000 300196 104002
rect 297449 103944 297454 104000
rect 297510 103944 300196 104000
rect 297449 103942 300196 103944
rect 339940 104000 341491 104002
rect 339940 103944 341430 104000
rect 341486 103944 341491 104000
rect 339940 103942 341491 103944
rect 297449 103939 297515 103942
rect 341425 103939 341491 103942
rect 57697 103186 57763 103189
rect 57697 103184 60076 103186
rect 57697 103128 57702 103184
rect 57758 103128 60076 103184
rect 57697 103126 60076 103128
rect 57697 103123 57763 103126
rect 296989 102506 297055 102509
rect 296989 102504 300196 102506
rect 296989 102448 296994 102504
rect 297050 102448 300196 102504
rect 296989 102446 300196 102448
rect 296989 102443 297055 102446
rect 341517 101826 341583 101829
rect 339940 101824 341583 101826
rect 339940 101768 341522 101824
rect 341578 101768 341583 101824
rect 339940 101766 341583 101768
rect 341517 101763 341583 101766
rect 223481 101418 223547 101421
rect 219788 101416 223547 101418
rect 219788 101360 223486 101416
rect 223542 101360 223547 101416
rect 219788 101358 223547 101360
rect 223481 101355 223547 101358
rect 299289 101010 299355 101013
rect 299289 101008 300196 101010
rect 299289 100952 299294 101008
rect 299350 100952 300196 101008
rect 299289 100950 300196 100952
rect 299289 100947 299355 100950
rect 341609 99650 341675 99653
rect 339940 99648 341675 99650
rect 339940 99592 341614 99648
rect 341670 99592 341675 99648
rect 339940 99590 341675 99592
rect 341609 99587 341675 99590
rect 297541 99514 297607 99517
rect 297541 99512 300196 99514
rect 297541 99456 297546 99512
rect 297602 99456 300196 99512
rect 297541 99454 300196 99456
rect 297541 99451 297607 99454
rect 355174 99452 355180 99516
rect 355244 99514 355250 99516
rect 583520 99514 584960 99604
rect 355244 99454 584960 99514
rect 355244 99452 355250 99454
rect 583520 99364 584960 99454
rect 59261 99106 59327 99109
rect 59261 99104 60076 99106
rect 59261 99048 59266 99104
rect 59322 99048 60076 99104
rect 59261 99046 60076 99048
rect 59261 99043 59327 99046
rect 223021 98562 223087 98565
rect 219788 98560 223087 98562
rect 219788 98504 223026 98560
rect 223082 98504 223087 98560
rect 219788 98502 223087 98504
rect 223021 98499 223087 98502
rect 298737 98018 298803 98021
rect 298737 98016 300196 98018
rect 298737 97960 298742 98016
rect 298798 97960 300196 98016
rect 298737 97958 300196 97960
rect 298737 97955 298803 97958
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 341701 97474 341767 97477
rect 339940 97472 341767 97474
rect 339940 97416 341706 97472
rect 341762 97416 341767 97472
rect 339940 97414 341767 97416
rect 341701 97411 341767 97414
rect 297817 96522 297883 96525
rect 297817 96520 300196 96522
rect 297817 96464 297822 96520
rect 297878 96464 300196 96520
rect 297817 96462 300196 96464
rect 297817 96459 297883 96462
rect 223113 95706 223179 95709
rect 219788 95704 223179 95706
rect 219788 95648 223118 95704
rect 223174 95648 223179 95704
rect 219788 95646 223179 95648
rect 223113 95643 223179 95646
rect 341006 95298 341012 95300
rect 339940 95238 341012 95298
rect 341006 95236 341012 95238
rect 341076 95236 341082 95300
rect 59721 95026 59787 95029
rect 297633 95026 297699 95029
rect 59721 95024 60076 95026
rect 59721 94968 59726 95024
rect 59782 94968 60076 95024
rect 59721 94966 60076 94968
rect 297633 95024 300196 95026
rect 297633 94968 297638 95024
rect 297694 94968 300196 95024
rect 297633 94966 300196 94968
rect 59721 94963 59787 94966
rect 297633 94963 297699 94966
rect 298829 93530 298895 93533
rect 298829 93528 300196 93530
rect 298829 93472 298834 93528
rect 298890 93472 300196 93528
rect 298829 93470 300196 93472
rect 298829 93467 298895 93470
rect 342345 93122 342411 93125
rect 339940 93120 342411 93122
rect 339940 93064 342350 93120
rect 342406 93064 342411 93120
rect 339940 93062 342411 93064
rect 342345 93059 342411 93062
rect 223481 92850 223547 92853
rect 219788 92848 223547 92850
rect 219788 92792 223486 92848
rect 223542 92792 223547 92848
rect 219788 92790 223547 92792
rect 223481 92787 223547 92790
rect 297081 92034 297147 92037
rect 297081 92032 300196 92034
rect 297081 91976 297086 92032
rect 297142 91976 300196 92032
rect 297081 91974 300196 91976
rect 297081 91971 297147 91974
rect 59077 90946 59143 90949
rect 342805 90946 342871 90949
rect 59077 90944 60076 90946
rect 59077 90888 59082 90944
rect 59138 90888 60076 90944
rect 59077 90886 60076 90888
rect 339940 90944 342871 90946
rect 339940 90888 342810 90944
rect 342866 90888 342871 90944
rect 339940 90886 342871 90888
rect 59077 90883 59143 90886
rect 342805 90883 342871 90886
rect 298001 90538 298067 90541
rect 298001 90536 300196 90538
rect 298001 90480 298006 90536
rect 298062 90480 300196 90536
rect 298001 90478 300196 90480
rect 298001 90475 298067 90478
rect 223481 89994 223547 89997
rect 219788 89992 223547 89994
rect 219788 89936 223486 89992
rect 223542 89936 223547 89992
rect 219788 89934 223547 89936
rect 223481 89931 223547 89934
rect 299381 89042 299447 89045
rect 299381 89040 300196 89042
rect 299381 88984 299386 89040
rect 299442 88984 300196 89040
rect 299381 88982 300196 88984
rect 299381 88979 299447 88982
rect 342897 88770 342963 88773
rect 339940 88768 342963 88770
rect 339940 88712 342902 88768
rect 342958 88712 342963 88768
rect 339940 88710 342963 88712
rect 342897 88707 342963 88710
rect 298001 87546 298067 87549
rect 298001 87544 300196 87546
rect 298001 87488 298006 87544
rect 298062 87488 300196 87544
rect 298001 87486 300196 87488
rect 298001 87483 298067 87486
rect 223205 87138 223271 87141
rect 219788 87136 223271 87138
rect 219788 87080 223210 87136
rect 223266 87080 223271 87136
rect 219788 87078 223271 87080
rect 223205 87075 223271 87078
rect 57789 86866 57855 86869
rect 57789 86864 60076 86866
rect 57789 86808 57794 86864
rect 57850 86808 60076 86864
rect 57789 86806 60076 86808
rect 57789 86803 57855 86806
rect 343173 86594 343239 86597
rect 339940 86592 343239 86594
rect 339940 86536 343178 86592
rect 343234 86536 343239 86592
rect 339940 86534 343239 86536
rect 343173 86531 343239 86534
rect 580257 86186 580323 86189
rect 583520 86186 584960 86276
rect 580257 86184 584960 86186
rect 580257 86128 580262 86184
rect 580318 86128 584960 86184
rect 580257 86126 584960 86128
rect 580257 86123 580323 86126
rect 297173 86050 297239 86053
rect 297173 86048 300196 86050
rect 297173 85992 297178 86048
rect 297234 85992 300196 86048
rect 583520 86036 584960 86126
rect 297173 85990 300196 85992
rect 297173 85987 297239 85990
rect 340086 85444 340092 85508
rect 340156 85506 340162 85508
rect 342294 85506 342300 85508
rect 340156 85446 342300 85506
rect 340156 85444 340162 85446
rect 342294 85444 342300 85446
rect 342364 85444 342370 85508
rect -960 84690 480 84780
rect 3417 84690 3483 84693
rect -960 84688 3483 84690
rect -960 84632 3422 84688
rect 3478 84632 3483 84688
rect -960 84630 3483 84632
rect -960 84540 480 84630
rect 3417 84627 3483 84630
rect 296805 84554 296871 84557
rect 296805 84552 300196 84554
rect 296805 84496 296810 84552
rect 296866 84496 300196 84552
rect 296805 84494 300196 84496
rect 296805 84491 296871 84494
rect 342478 84418 342484 84420
rect 339940 84358 342484 84418
rect 342478 84356 342484 84358
rect 342548 84356 342554 84420
rect 223205 84282 223271 84285
rect 219788 84280 223271 84282
rect 219788 84224 223210 84280
rect 223266 84224 223271 84280
rect 219788 84222 223271 84224
rect 223205 84219 223271 84222
rect 297909 83058 297975 83061
rect 297909 83056 300196 83058
rect 297909 83000 297914 83056
rect 297970 83000 300196 83056
rect 297909 82998 300196 83000
rect 297909 82995 297975 82998
rect 58985 82786 59051 82789
rect 58985 82784 60076 82786
rect 58985 82728 58990 82784
rect 59046 82728 60076 82784
rect 58985 82726 60076 82728
rect 58985 82723 59051 82726
rect 342294 82242 342300 82244
rect 339940 82182 342300 82242
rect 342294 82180 342300 82182
rect 342364 82180 342370 82244
rect 297909 81562 297975 81565
rect 297909 81560 300196 81562
rect 297909 81504 297914 81560
rect 297970 81504 300196 81560
rect 297909 81502 300196 81504
rect 297909 81499 297975 81502
rect 223481 81426 223547 81429
rect 219788 81424 223547 81426
rect 219788 81368 223486 81424
rect 223542 81368 223547 81424
rect 219788 81366 223547 81368
rect 223481 81363 223547 81366
rect 298001 80066 298067 80069
rect 298001 80064 300196 80066
rect 298001 80008 298006 80064
rect 298062 80008 300196 80064
rect 298001 80006 300196 80008
rect 339940 80006 340890 80066
rect 298001 80003 298067 80006
rect 340830 79250 340890 80006
rect 341374 79324 341380 79388
rect 341444 79386 341450 79388
rect 342345 79386 342411 79389
rect 341444 79384 342411 79386
rect 341444 79328 342350 79384
rect 342406 79328 342411 79384
rect 341444 79326 342411 79328
rect 341444 79324 341450 79326
rect 342345 79323 342411 79326
rect 342345 79250 342411 79253
rect 340830 79248 342411 79250
rect 340830 79192 342350 79248
rect 342406 79192 342411 79248
rect 340830 79190 342411 79192
rect 342345 79187 342411 79190
rect 57881 78706 57947 78709
rect 57881 78704 60076 78706
rect 57881 78648 57886 78704
rect 57942 78648 60076 78704
rect 57881 78646 60076 78648
rect 57881 78643 57947 78646
rect 222469 78570 222535 78573
rect 219788 78568 222535 78570
rect 219788 78512 222474 78568
rect 222530 78512 222535 78568
rect 219788 78510 222535 78512
rect 222469 78507 222535 78510
rect 297541 78570 297607 78573
rect 297541 78568 300196 78570
rect 297541 78512 297546 78568
rect 297602 78512 300196 78568
rect 297541 78510 300196 78512
rect 297541 78507 297607 78510
rect 342662 77890 342668 77892
rect 339940 77830 342668 77890
rect 342662 77828 342668 77830
rect 342732 77828 342738 77892
rect 297173 77074 297239 77077
rect 297173 77072 300196 77074
rect 297173 77016 297178 77072
rect 297234 77016 300196 77072
rect 297173 77014 300196 77016
rect 297173 77011 297239 77014
rect 222193 75714 222259 75717
rect 340505 75714 340571 75717
rect 219788 75712 222259 75714
rect 219788 75656 222198 75712
rect 222254 75656 222259 75712
rect 219788 75654 222259 75656
rect 339940 75712 340571 75714
rect 339940 75656 340510 75712
rect 340566 75656 340571 75712
rect 339940 75654 340571 75656
rect 222193 75651 222259 75654
rect 340505 75651 340571 75654
rect 298001 75578 298067 75581
rect 298001 75576 300196 75578
rect 298001 75520 298006 75576
rect 298062 75520 300196 75576
rect 298001 75518 300196 75520
rect 298001 75515 298067 75518
rect 59629 74626 59695 74629
rect 59629 74624 60076 74626
rect 59629 74568 59634 74624
rect 59690 74568 60076 74624
rect 59629 74566 60076 74568
rect 59629 74563 59695 74566
rect 298001 74082 298067 74085
rect 298001 74080 300196 74082
rect 298001 74024 298006 74080
rect 298062 74024 300196 74080
rect 298001 74022 300196 74024
rect 298001 74019 298067 74022
rect 340270 73538 340276 73540
rect 339940 73478 340276 73538
rect 340270 73476 340276 73478
rect 340340 73476 340346 73540
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 222193 72858 222259 72861
rect 219788 72856 222259 72858
rect 219788 72800 222198 72856
rect 222254 72800 222259 72856
rect 583520 72844 584960 72934
rect 219788 72798 222259 72800
rect 222193 72795 222259 72798
rect 296805 72586 296871 72589
rect 296805 72584 300196 72586
rect 296805 72528 296810 72584
rect 296866 72528 300196 72584
rect 296805 72526 300196 72528
rect 296805 72523 296871 72526
rect -960 71484 480 71724
rect 341190 71362 341196 71364
rect 339940 71302 341196 71362
rect 341190 71300 341196 71302
rect 341260 71300 341266 71364
rect 297725 71090 297791 71093
rect 297725 71088 300196 71090
rect 297725 71032 297730 71088
rect 297786 71032 300196 71088
rect 297725 71030 300196 71032
rect 297725 71027 297791 71030
rect 59353 70546 59419 70549
rect 59353 70544 60076 70546
rect 59353 70488 59358 70544
rect 59414 70488 60076 70544
rect 59353 70486 60076 70488
rect 59353 70483 59419 70486
rect 223481 70002 223547 70005
rect 219788 70000 223547 70002
rect 219788 69944 223486 70000
rect 223542 69944 223547 70000
rect 219788 69942 223547 69944
rect 223481 69939 223547 69942
rect 298001 69594 298067 69597
rect 298001 69592 300196 69594
rect 298001 69536 298006 69592
rect 298062 69536 300196 69592
rect 298001 69534 300196 69536
rect 298001 69531 298067 69534
rect 342989 69186 343055 69189
rect 339940 69184 343055 69186
rect 339940 69128 342994 69184
rect 343050 69128 343055 69184
rect 339940 69126 343055 69128
rect 342989 69123 343055 69126
rect 297173 68098 297239 68101
rect 297173 68096 300196 68098
rect 297173 68040 297178 68096
rect 297234 68040 300196 68096
rect 297173 68038 300196 68040
rect 297173 68035 297239 68038
rect 223481 67146 223547 67149
rect 219788 67144 223547 67146
rect 219788 67088 223486 67144
rect 223542 67088 223547 67144
rect 219788 67086 223547 67088
rect 223481 67083 223547 67086
rect 342989 67010 343055 67013
rect 339940 67008 343055 67010
rect 339940 66952 342994 67008
rect 343050 66952 343055 67008
rect 339940 66950 343055 66952
rect 342989 66947 343055 66950
rect 297541 66602 297607 66605
rect 297541 66600 300196 66602
rect 297541 66544 297546 66600
rect 297602 66544 300196 66600
rect 297541 66542 300196 66544
rect 297541 66539 297607 66542
rect 59537 66466 59603 66469
rect 59537 66464 60076 66466
rect 59537 66408 59542 66464
rect 59598 66408 60076 66464
rect 59537 66406 60076 66408
rect 59537 66403 59603 66406
rect 297357 65106 297423 65109
rect 297357 65104 300196 65106
rect 297357 65048 297362 65104
rect 297418 65048 300196 65104
rect 297357 65046 300196 65048
rect 297357 65043 297423 65046
rect 342989 64834 343055 64837
rect 339940 64832 343055 64834
rect 339940 64776 342994 64832
rect 343050 64776 343055 64832
rect 339940 64774 343055 64776
rect 342989 64771 343055 64774
rect 222837 64290 222903 64293
rect 219788 64288 222903 64290
rect 219788 64232 222842 64288
rect 222898 64232 222903 64288
rect 219788 64230 222903 64232
rect 222837 64227 222903 64230
rect 297909 63610 297975 63613
rect 297909 63608 300196 63610
rect 297909 63552 297914 63608
rect 297970 63552 300196 63608
rect 297909 63550 300196 63552
rect 297909 63547 297975 63550
rect 342345 62658 342411 62661
rect 339940 62656 342411 62658
rect 339940 62600 342350 62656
rect 342406 62600 342411 62656
rect 339940 62598 342411 62600
rect 342345 62595 342411 62598
rect 59169 62386 59235 62389
rect 59169 62384 60076 62386
rect 59169 62328 59174 62384
rect 59230 62328 60076 62384
rect 59169 62326 60076 62328
rect 59169 62323 59235 62326
rect 298001 62114 298067 62117
rect 298001 62112 300196 62114
rect 298001 62056 298006 62112
rect 298062 62056 300196 62112
rect 298001 62054 300196 62056
rect 298001 62051 298067 62054
rect 165613 61570 165679 61573
rect 341006 61570 341012 61572
rect 165613 61568 341012 61570
rect 165613 61512 165618 61568
rect 165674 61512 341012 61568
rect 165613 61510 341012 61512
rect 165613 61507 165679 61510
rect 341006 61508 341012 61510
rect 341076 61508 341082 61572
rect 126973 61434 127039 61437
rect 341190 61434 341196 61436
rect 126973 61432 341196 61434
rect 126973 61376 126978 61432
rect 127034 61376 341196 61432
rect 126973 61374 341196 61376
rect 126973 61371 127039 61374
rect 341190 61372 341196 61374
rect 341260 61372 341266 61436
rect 317413 60074 317479 60077
rect 349286 60074 349292 60076
rect 317413 60072 349292 60074
rect 317413 60016 317418 60072
rect 317474 60016 349292 60072
rect 317413 60014 349292 60016
rect 317413 60011 317479 60014
rect 349286 60012 349292 60014
rect 349356 60012 349362 60076
rect 136633 59938 136699 59941
rect 342662 59938 342668 59940
rect 136633 59936 342668 59938
rect 136633 59880 136638 59936
rect 136694 59880 342668 59936
rect 136633 59878 342668 59880
rect 136633 59875 136699 59878
rect 342662 59876 342668 59878
rect 342732 59876 342738 59940
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 147673 57218 147739 57221
rect 342478 57218 342484 57220
rect 147673 57216 342484 57218
rect 147673 57160 147678 57216
rect 147734 57160 342484 57216
rect 147673 57158 342484 57160
rect 147673 57155 147739 57158
rect 342478 57156 342484 57158
rect 342548 57156 342554 57220
rect 129733 55858 129799 55861
rect 340270 55858 340276 55860
rect 129733 55856 340276 55858
rect 129733 55800 129738 55856
rect 129794 55800 340276 55856
rect 129733 55798 340276 55800
rect 129733 55795 129799 55798
rect 340270 55796 340276 55798
rect 340340 55796 340346 55860
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 403566 44780 403572 44844
rect 403636 44842 403642 44844
rect 444373 44842 444439 44845
rect 403636 44840 444439 44842
rect 403636 44784 444378 44840
rect 444434 44784 444439 44840
rect 403636 44782 444439 44784
rect 403636 44780 403642 44782
rect 444373 44779 444439 44782
rect 186313 39266 186379 39269
rect 340822 39266 340828 39268
rect 186313 39264 340828 39266
rect 186313 39208 186318 39264
rect 186374 39208 340828 39264
rect 186313 39206 340828 39208
rect 186313 39203 186379 39206
rect 340822 39204 340828 39206
rect 340892 39204 340898 39268
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 92473 24170 92539 24173
rect 404854 24170 404860 24172
rect 92473 24168 404860 24170
rect 92473 24112 92478 24168
rect 92534 24112 404860 24168
rect 92473 24110 404860 24112
rect 92473 24107 92539 24110
rect 404854 24108 404860 24110
rect 404924 24108 404930 24172
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 24209 8938 24275 8941
rect 521694 8938 521700 8940
rect 24209 8936 521700 8938
rect 24209 8880 24214 8936
rect 24270 8880 521700 8936
rect 24209 8878 521700 8880
rect 24209 8875 24275 8878
rect 521694 8876 521700 8878
rect 521764 8876 521770 8940
rect 71497 7578 71563 7581
rect 494646 7578 494652 7580
rect 71497 7576 494652 7578
rect 71497 7520 71502 7576
rect 71558 7520 494652 7576
rect 71497 7518 494652 7520
rect 71497 7515 71563 7518
rect 494646 7516 494652 7518
rect 494716 7516 494722 7580
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 67909 6218 67975 6221
rect 512494 6218 512500 6220
rect 67909 6216 512500 6218
rect 67909 6160 67914 6216
rect 67970 6160 512500 6216
rect 67909 6158 512500 6160
rect 67909 6155 67975 6158
rect 512494 6156 512500 6158
rect 512564 6156 512570 6220
rect 144729 5130 144795 5133
rect 342294 5130 342300 5132
rect 144729 5128 342300 5130
rect 144729 5072 144734 5128
rect 144790 5072 342300 5128
rect 144729 5070 342300 5072
rect 144729 5067 144795 5070
rect 342294 5068 342300 5070
rect 342364 5068 342370 5132
rect 254669 4994 254735 4997
rect 484342 4994 484348 4996
rect 254669 4992 484348 4994
rect 254669 4936 254674 4992
rect 254730 4936 484348 4992
rect 254669 4934 484348 4936
rect 254669 4931 254735 4934
rect 484342 4932 484348 4934
rect 484412 4932 484418 4996
rect 53741 4858 53807 4861
rect 518934 4858 518940 4860
rect 53741 4856 518940 4858
rect 53741 4800 53746 4856
rect 53802 4800 518940 4856
rect 53741 4798 518940 4800
rect 53741 4795 53807 4798
rect 518934 4796 518940 4798
rect 519004 4796 519010 4860
rect 505502 3980 505508 4044
rect 505572 4042 505578 4044
rect 510061 4042 510127 4045
rect 505572 4040 510127 4042
rect 505572 3984 510066 4040
rect 510122 3984 510127 4040
rect 505572 3982 510127 3984
rect 505572 3980 505578 3982
rect 510061 3979 510127 3982
rect 297265 3634 297331 3637
rect 298502 3634 298508 3636
rect 297265 3632 298508 3634
rect 297265 3576 297270 3632
rect 297326 3576 298508 3632
rect 297265 3574 298508 3576
rect 297265 3571 297331 3574
rect 298502 3572 298508 3574
rect 298572 3572 298578 3636
rect 299790 3572 299796 3636
rect 299860 3634 299866 3636
rect 300761 3634 300827 3637
rect 299860 3632 300827 3634
rect 299860 3576 300766 3632
rect 300822 3576 300827 3632
rect 299860 3574 300827 3576
rect 299860 3572 299866 3574
rect 300761 3571 300827 3574
rect 329189 3634 329255 3637
rect 349102 3634 349108 3636
rect 329189 3632 349108 3634
rect 329189 3576 329194 3632
rect 329250 3576 349108 3632
rect 329189 3574 349108 3576
rect 329189 3571 329255 3574
rect 349102 3572 349108 3574
rect 349172 3572 349178 3636
rect 183737 3498 183803 3501
rect 340086 3498 340092 3500
rect 183737 3496 340092 3498
rect 183737 3440 183742 3496
rect 183798 3440 340092 3496
rect 183737 3438 340092 3440
rect 183737 3435 183803 3438
rect 340086 3436 340092 3438
rect 340156 3436 340162 3500
rect 502190 3436 502196 3500
rect 502260 3498 502266 3500
rect 502977 3498 503043 3501
rect 502260 3496 503043 3498
rect 502260 3440 502982 3496
rect 503038 3440 503043 3496
rect 502260 3438 503043 3440
rect 502260 3436 502266 3438
rect 502977 3435 503043 3438
rect 513557 3498 513623 3501
rect 516358 3498 516364 3500
rect 513557 3496 516364 3498
rect 513557 3440 513562 3496
rect 513618 3440 516364 3496
rect 513557 3438 516364 3440
rect 513557 3435 513623 3438
rect 516358 3436 516364 3438
rect 516428 3436 516434 3500
rect 162485 3362 162551 3365
rect 341374 3362 341380 3364
rect 162485 3360 341380 3362
rect 162485 3304 162490 3360
rect 162546 3304 341380 3360
rect 162485 3302 341380 3304
rect 162485 3299 162551 3302
rect 341374 3300 341380 3302
rect 341444 3300 341450 3364
rect 495893 3362 495959 3365
rect 511206 3362 511212 3364
rect 495893 3360 511212 3362
rect 495893 3304 495898 3360
rect 495954 3304 511212 3360
rect 495893 3302 511212 3304
rect 495893 3299 495959 3302
rect 511206 3300 511212 3302
rect 511276 3300 511282 3364
<< via3 >>
rect 360700 700300 360764 700364
rect 283420 663172 283484 663236
rect 405044 663036 405108 663100
rect 286180 662900 286244 662964
rect 317644 662764 317708 662828
rect 51028 662628 51092 662692
rect 401548 662628 401612 662692
rect 51580 662492 51644 662556
rect 403020 662492 403084 662556
rect 282316 661812 282380 661876
rect 295012 661676 295076 661740
rect 295932 661540 295996 661604
rect 297220 661404 297284 661468
rect 311020 661404 311084 661468
rect 308628 661268 308692 661332
rect 359964 661268 360028 661332
rect 401732 661268 401796 661332
rect 49004 661132 49068 661196
rect 309364 661132 309428 661196
rect 309180 660996 309244 661060
rect 279372 660588 279436 660652
rect 49372 660452 49436 660516
rect 308812 660316 308876 660380
rect 49188 660180 49252 660244
rect 310468 660180 310532 660244
rect 502932 660180 502996 660244
rect 508452 660180 508516 660244
rect 311940 660044 312004 660108
rect 489684 659908 489748 659972
rect 49924 659772 49988 659836
rect 49740 659636 49804 659700
rect 50108 659636 50172 659700
rect 398604 642092 398668 642156
rect 358860 641956 358924 642020
rect 363460 641684 363524 641748
rect 304764 641004 304828 641068
rect 306236 640868 306300 640932
rect 351132 640596 351196 640660
rect 355180 640460 355244 640524
rect 301452 640324 301516 640388
rect 358676 639644 358740 639708
rect 362724 639508 362788 639572
rect 355364 639372 355428 639436
rect 362356 639372 362420 639436
rect 362540 639432 362604 639436
rect 362540 639376 362590 639432
rect 362590 639376 362604 639432
rect 362540 639372 362604 639376
rect 364012 639432 364076 639436
rect 364012 639376 364062 639432
rect 364062 639376 364076 639432
rect 364012 639372 364076 639376
rect 377260 639644 377324 639708
rect 381124 639508 381188 639572
rect 285444 639296 285508 639300
rect 285444 639240 285458 639296
rect 285458 639240 285508 639296
rect 285444 639236 285508 639240
rect 288204 639296 288268 639300
rect 288204 639240 288254 639296
rect 288254 639240 288268 639296
rect 288204 639236 288268 639240
rect 289492 639236 289556 639300
rect 290964 639296 291028 639300
rect 290964 639240 290978 639296
rect 290978 639240 291028 639296
rect 290964 639236 291028 639240
rect 292436 639236 292500 639300
rect 293724 639236 293788 639300
rect 298508 639296 298572 639300
rect 298508 639240 298522 639296
rect 298522 639240 298572 639296
rect 298508 639236 298572 639240
rect 306972 639236 307036 639300
rect 300716 639100 300780 639164
rect 377260 639100 377324 639164
rect 303476 638964 303540 639028
rect 381124 638964 381188 639028
rect 49372 637604 49436 637668
rect 49372 637468 49436 637532
rect 50108 618292 50172 618356
rect 49188 614212 49252 614276
rect 49556 612716 49620 612780
rect 49556 608364 49620 608428
rect 49556 607140 49620 607204
rect 49924 605916 49988 605980
rect 49004 602516 49068 602580
rect 49188 601020 49252 601084
rect 51580 601020 51644 601084
rect 303476 600672 303540 600676
rect 303476 600616 303490 600672
rect 303490 600616 303540 600672
rect 303476 600612 303540 600616
rect 304764 600672 304828 600676
rect 304764 600616 304778 600672
rect 304778 600616 304828 600672
rect 304764 600612 304828 600616
rect 306236 600672 306300 600676
rect 306236 600616 306250 600672
rect 306250 600616 306300 600672
rect 306236 600612 306300 600616
rect 306972 600476 307036 600540
rect 300716 600128 300780 600132
rect 300716 600072 300730 600128
rect 300730 600072 300780 600128
rect 300716 600068 300780 600072
rect 369900 599524 369964 599588
rect 301452 598844 301516 598908
rect 382228 598164 382292 598228
rect 306972 597680 307036 597684
rect 306972 597624 307022 597680
rect 307022 597624 307036 597680
rect 306972 597620 307036 597624
rect 368980 597620 369044 597684
rect 362356 595444 362420 595508
rect 362908 593268 362972 593332
rect 363460 593132 363524 593196
rect 380940 589868 381004 589932
rect 376156 587148 376220 587212
rect 384068 582932 384132 582996
rect 364012 581708 364076 581772
rect 292436 581572 292500 581636
rect 373212 581572 373276 581636
rect 394740 580348 394804 580412
rect 389588 580212 389652 580276
rect 385540 579532 385604 579596
rect 376892 578852 376956 578916
rect 391980 577492 392044 577556
rect 394004 575452 394068 575516
rect 391060 573276 391124 573340
rect 361620 571916 361684 571980
rect 377260 569332 377324 569396
rect 290964 569196 291028 569260
rect 380572 569196 380636 569260
rect 366220 568516 366284 568580
rect 378732 565796 378796 565860
rect 362540 564980 362604 565044
rect 385724 564436 385788 564500
rect 364748 563620 364812 563684
rect 368244 563620 368308 563684
rect 382780 563620 382844 563684
rect 371556 563076 371620 563140
rect 386460 562396 386524 562460
rect 289492 562260 289556 562324
rect 400628 562260 400692 562324
rect 376340 561172 376404 561236
rect 298508 561036 298572 561100
rect 400444 561036 400508 561100
rect 285444 560900 285508 560964
rect 399156 560900 399220 560964
rect 358308 559676 358372 559740
rect 398788 559540 398852 559604
rect 361436 558316 361500 558380
rect 288204 558180 288268 558244
rect 400260 556684 400324 556748
rect 358124 555460 358188 555524
rect 399340 555324 399404 555388
rect 358492 554100 358556 554164
rect 359044 553964 359108 554028
rect 359964 552604 360028 552668
rect 403572 552060 403636 552124
rect 359228 551924 359292 551988
rect 359412 551652 359476 551716
rect 362724 551516 362788 551580
rect 400812 551380 400876 551444
rect 293724 551244 293788 551308
rect 398972 551244 399036 551308
rect 401916 550020 401980 550084
rect 401732 549204 401796 549268
rect 358124 547300 358188 547364
rect 295932 543628 295996 543692
rect 317644 543628 317708 543692
rect 401916 543628 401980 543692
rect 489868 543628 489932 543692
rect 295012 543492 295076 543556
rect 508452 543492 508516 543556
rect 286180 543356 286244 543420
rect 297220 543356 297284 543420
rect 283420 543220 283484 543284
rect 279372 543084 279436 543148
rect 311940 543084 312004 543148
rect 282316 542948 282380 543012
rect 282132 542676 282196 542740
rect 308812 542540 308876 542604
rect 309364 542540 309428 542604
rect 310468 542540 310532 542604
rect 308628 542464 308692 542468
rect 308628 542408 308678 542464
rect 308678 542408 308692 542464
rect 308628 542404 308692 542408
rect 309180 542404 309244 542468
rect 311020 542464 311084 542468
rect 311020 542408 311070 542464
rect 311070 542408 311084 542464
rect 311020 542404 311084 542408
rect 359412 541996 359476 542060
rect 495940 541044 496004 541108
rect 511212 541044 511276 541108
rect 358308 540636 358372 540700
rect 485636 539820 485700 539884
rect 512500 539820 512564 539884
rect 287284 539684 287348 539748
rect 288572 539684 288636 539748
rect 290596 539684 290660 539748
rect 486372 539684 486436 539748
rect 494652 539684 494716 539748
rect 502196 539744 502260 539748
rect 502196 539688 502210 539744
rect 502210 539688 502260 539744
rect 502196 539684 502260 539688
rect 505508 539744 505572 539748
rect 505508 539688 505558 539744
rect 505558 539688 505572 539744
rect 505508 539684 505572 539688
rect 516364 539744 516428 539748
rect 516364 539688 516414 539744
rect 516414 539688 516428 539744
rect 516364 539684 516428 539688
rect 284892 539548 284956 539612
rect 285996 539548 286060 539612
rect 287652 539608 287716 539612
rect 287652 539552 287666 539608
rect 287666 539552 287716 539608
rect 287652 539548 287716 539552
rect 288388 539548 288452 539612
rect 290780 539608 290844 539612
rect 290780 539552 290794 539608
rect 290794 539552 290844 539608
rect 290780 539548 290844 539552
rect 291148 539548 291212 539612
rect 292620 539548 292684 539612
rect 293908 539548 293972 539612
rect 295380 539548 295444 539612
rect 401548 539548 401612 539612
rect 521884 538460 521948 538524
rect 404860 538188 404924 538252
rect 400628 537780 400692 537844
rect 519308 533836 519372 533900
rect 522068 532748 522132 532812
rect 49188 532340 49252 532404
rect 400812 531796 400876 531860
rect 405044 531524 405108 531588
rect 359228 530572 359292 530636
rect 358676 527716 358740 527780
rect 399340 527716 399404 527780
rect 519308 523364 519372 523428
rect 400444 523160 400508 523224
rect 349108 518876 349172 518940
rect 399340 518604 399404 518668
rect 358492 516836 358556 516900
rect 403020 513300 403084 513364
rect 399340 507724 399404 507788
rect 399524 505956 399588 506020
rect 359044 505004 359108 505068
rect 49556 503160 49620 503164
rect 49556 503104 49606 503160
rect 49606 503104 49620 503160
rect 49556 503100 49620 503104
rect 521700 502964 521764 503028
rect 358860 502284 358924 502348
rect 400260 501400 400324 501464
rect 49740 500924 49804 500988
rect 361436 499836 361500 499900
rect 362908 499896 362972 499900
rect 362908 499840 362958 499896
rect 362958 499840 362972 499896
rect 362908 499836 362972 499840
rect 364748 499836 364812 499900
rect 368244 499836 368308 499900
rect 369900 499836 369964 499900
rect 371556 499896 371620 499900
rect 371556 499840 371606 499896
rect 371606 499840 371620 499896
rect 371556 499836 371620 499840
rect 376156 499836 376220 499900
rect 376892 499836 376956 499900
rect 380572 499896 380636 499900
rect 380572 499840 380622 499896
rect 380622 499840 380636 499896
rect 380572 499836 380636 499840
rect 380940 499836 381004 499900
rect 382780 499836 382844 499900
rect 385540 499836 385604 499900
rect 386460 499836 386524 499900
rect 389588 499836 389652 499900
rect 391980 499836 392044 499900
rect 394740 499836 394804 499900
rect 398604 499836 398668 499900
rect 502932 499836 502996 499900
rect 361620 499700 361684 499764
rect 385724 499700 385788 499764
rect 495940 499564 496004 499628
rect 366220 499428 366284 499492
rect 368980 499428 369044 499492
rect 376340 499428 376404 499492
rect 360700 499292 360764 499356
rect 298324 498748 298388 498812
rect 373212 498068 373276 498132
rect 377260 498068 377324 498132
rect 384068 498068 384132 498132
rect 378732 497932 378796 497996
rect 391060 497932 391124 497996
rect 394004 497524 394068 497588
rect 382228 497388 382292 497452
rect 349292 496844 349356 496908
rect 484348 496844 484412 496908
rect 485636 496844 485700 496908
rect 51028 485556 51092 485620
rect 49556 484392 49620 484396
rect 49556 484336 49606 484392
rect 49606 484336 49620 484392
rect 49556 484332 49620 484336
rect 49372 479708 49436 479772
rect 298508 349692 298572 349756
rect 299796 335956 299860 336020
rect 299612 331196 299676 331260
rect 351868 320180 351932 320244
rect 297220 309980 297284 310044
rect 284892 292572 284956 292636
rect 298324 282372 298388 282436
rect 291148 281964 291212 282028
rect 285996 281828 286060 281892
rect 288572 281420 288636 281484
rect 486372 281420 486436 281484
rect 290780 281284 290844 281348
rect 290596 281148 290660 281212
rect 287284 281012 287348 281076
rect 288388 280876 288452 280940
rect 287652 280740 287716 280804
rect 282132 280604 282196 280668
rect 292620 280468 292684 280532
rect 295380 280060 295444 280124
rect 293908 279924 293972 279988
rect 297220 279380 297284 279444
rect 49372 278700 49436 278764
rect 355364 258028 355428 258092
rect 57836 227020 57900 227084
rect 522068 226884 522132 226948
rect 351868 225524 351932 225588
rect 521884 224300 521948 224364
rect 519124 224164 519188 224228
rect 49556 223484 49620 223548
rect 351132 218044 351196 218108
rect 299612 216684 299676 216748
rect 57836 131684 57900 131748
rect 340828 108292 340892 108356
rect 342300 106176 342364 106180
rect 342300 106120 342350 106176
rect 342350 106120 342364 106176
rect 342300 106116 342364 106120
rect 355180 99452 355244 99516
rect 341012 95236 341076 95300
rect 340092 85444 340156 85508
rect 342300 85444 342364 85508
rect 342484 84356 342548 84420
rect 342300 82180 342364 82244
rect 341380 79324 341444 79388
rect 342668 77828 342732 77892
rect 340276 73476 340340 73540
rect 341196 71300 341260 71364
rect 341012 61508 341076 61572
rect 341196 61372 341260 61436
rect 349292 60012 349356 60076
rect 342668 59876 342732 59940
rect 342484 57156 342548 57220
rect 340276 55796 340340 55860
rect 403572 44780 403636 44844
rect 340828 39204 340892 39268
rect 404860 24108 404924 24172
rect 521700 8876 521764 8940
rect 494652 7516 494716 7580
rect 512500 6156 512564 6220
rect 342300 5068 342364 5132
rect 484348 4932 484412 4996
rect 518940 4796 519004 4860
rect 505508 3980 505572 4044
rect 298508 3572 298572 3636
rect 299796 3572 299860 3636
rect 349108 3572 349172 3636
rect 340092 3436 340156 3500
rect 502196 3436 502260 3500
rect 516364 3436 516428 3500
rect 341380 3300 341444 3364
rect 511212 3300 511276 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 682954 -8106 711002
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 -8106 682954
rect -8726 682634 -8106 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 -8106 682634
rect -8726 646954 -8106 682398
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 -8106 646954
rect -8726 646634 -8106 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 -8106 646634
rect -8726 610954 -8106 646398
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 -8106 610954
rect -8726 610634 -8106 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 -8106 610634
rect -8726 574954 -8106 610398
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 -8106 574954
rect -8726 574634 -8106 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 -8106 574634
rect -8726 538954 -8106 574398
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 -8106 538954
rect -8726 538634 -8106 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 -8106 538634
rect -8726 502954 -8106 538398
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 -8106 502954
rect -8726 502634 -8106 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 -8106 502634
rect -8726 466954 -8106 502398
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 -8106 466954
rect -8726 466634 -8106 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 -8106 466634
rect -8726 430954 -8106 466398
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 -8106 430954
rect -8726 430634 -8106 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 -8106 430634
rect -8726 394954 -8106 430398
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 -8106 394954
rect -8726 394634 -8106 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 -8106 394634
rect -8726 358954 -8106 394398
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 -8106 358954
rect -8726 358634 -8106 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 -8106 358634
rect -8726 322954 -8106 358398
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 -8106 322954
rect -8726 322634 -8106 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 -8106 322634
rect -8726 286954 -8106 322398
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 -8106 286954
rect -8726 286634 -8106 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 -8106 286634
rect -8726 250954 -8106 286398
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 -8106 250954
rect -8726 250634 -8106 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 -8106 250634
rect -8726 214954 -8106 250398
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 -8106 214954
rect -8726 214634 -8106 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 -8106 214634
rect -8726 178954 -8106 214398
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 -8106 178954
rect -8726 178634 -8106 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 -8106 178634
rect -8726 142954 -8106 178398
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 -8106 142954
rect -8726 142634 -8106 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 -8106 142634
rect -8726 106954 -8106 142398
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 -8106 106954
rect -8726 106634 -8106 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 -8106 106634
rect -8726 70954 -8106 106398
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 -8106 70954
rect -8726 70634 -8106 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 -8106 70634
rect -8726 34954 -8106 70398
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 -8106 34954
rect -8726 34634 -8106 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 -8106 34634
rect -8726 -7066 -8106 34398
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 678454 -7146 710042
rect -7766 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 -7146 678454
rect -7766 678134 -7146 678218
rect -7766 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 -7146 678134
rect -7766 642454 -7146 677898
rect -7766 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 -7146 642454
rect -7766 642134 -7146 642218
rect -7766 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 -7146 642134
rect -7766 606454 -7146 641898
rect -7766 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 -7146 606454
rect -7766 606134 -7146 606218
rect -7766 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 -7146 606134
rect -7766 570454 -7146 605898
rect -7766 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 -7146 570454
rect -7766 570134 -7146 570218
rect -7766 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 -7146 570134
rect -7766 534454 -7146 569898
rect -7766 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 -7146 534454
rect -7766 534134 -7146 534218
rect -7766 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 -7146 534134
rect -7766 498454 -7146 533898
rect -7766 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 -7146 498454
rect -7766 498134 -7146 498218
rect -7766 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 -7146 498134
rect -7766 462454 -7146 497898
rect -7766 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 -7146 462454
rect -7766 462134 -7146 462218
rect -7766 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 -7146 462134
rect -7766 426454 -7146 461898
rect -7766 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 -7146 426454
rect -7766 426134 -7146 426218
rect -7766 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 -7146 426134
rect -7766 390454 -7146 425898
rect -7766 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 -7146 390454
rect -7766 390134 -7146 390218
rect -7766 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 -7146 390134
rect -7766 354454 -7146 389898
rect -7766 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 -7146 354454
rect -7766 354134 -7146 354218
rect -7766 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 -7146 354134
rect -7766 318454 -7146 353898
rect -7766 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 -7146 318454
rect -7766 318134 -7146 318218
rect -7766 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 -7146 318134
rect -7766 282454 -7146 317898
rect -7766 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 -7146 282454
rect -7766 282134 -7146 282218
rect -7766 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 -7146 282134
rect -7766 246454 -7146 281898
rect -7766 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 -7146 246454
rect -7766 246134 -7146 246218
rect -7766 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 -7146 246134
rect -7766 210454 -7146 245898
rect -7766 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 -7146 210454
rect -7766 210134 -7146 210218
rect -7766 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 -7146 210134
rect -7766 174454 -7146 209898
rect -7766 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 -7146 174454
rect -7766 174134 -7146 174218
rect -7766 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 -7146 174134
rect -7766 138454 -7146 173898
rect -7766 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 -7146 138454
rect -7766 138134 -7146 138218
rect -7766 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 -7146 138134
rect -7766 102454 -7146 137898
rect -7766 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 -7146 102454
rect -7766 102134 -7146 102218
rect -7766 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 -7146 102134
rect -7766 66454 -7146 101898
rect -7766 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 -7146 66454
rect -7766 66134 -7146 66218
rect -7766 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 -7146 66134
rect -7766 30454 -7146 65898
rect -7766 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 -7146 30454
rect -7766 30134 -7146 30218
rect -7766 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 -7146 30134
rect -7766 -6106 -7146 29898
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 673954 -6186 709082
rect -6806 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 -6186 673954
rect -6806 673634 -6186 673718
rect -6806 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 -6186 673634
rect -6806 637954 -6186 673398
rect -6806 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 -6186 637954
rect -6806 637634 -6186 637718
rect -6806 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 -6186 637634
rect -6806 601954 -6186 637398
rect -6806 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 -6186 601954
rect -6806 601634 -6186 601718
rect -6806 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 -6186 601634
rect -6806 565954 -6186 601398
rect -6806 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 -6186 565954
rect -6806 565634 -6186 565718
rect -6806 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 -6186 565634
rect -6806 529954 -6186 565398
rect -6806 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 -6186 529954
rect -6806 529634 -6186 529718
rect -6806 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 -6186 529634
rect -6806 493954 -6186 529398
rect -6806 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 -6186 493954
rect -6806 493634 -6186 493718
rect -6806 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 -6186 493634
rect -6806 457954 -6186 493398
rect -6806 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 -6186 457954
rect -6806 457634 -6186 457718
rect -6806 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 -6186 457634
rect -6806 421954 -6186 457398
rect -6806 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 -6186 421954
rect -6806 421634 -6186 421718
rect -6806 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 -6186 421634
rect -6806 385954 -6186 421398
rect -6806 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 -6186 385954
rect -6806 385634 -6186 385718
rect -6806 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 -6186 385634
rect -6806 349954 -6186 385398
rect -6806 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 -6186 349954
rect -6806 349634 -6186 349718
rect -6806 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 -6186 349634
rect -6806 313954 -6186 349398
rect -6806 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 -6186 313954
rect -6806 313634 -6186 313718
rect -6806 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 -6186 313634
rect -6806 277954 -6186 313398
rect -6806 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 -6186 277954
rect -6806 277634 -6186 277718
rect -6806 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 -6186 277634
rect -6806 241954 -6186 277398
rect -6806 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 -6186 241954
rect -6806 241634 -6186 241718
rect -6806 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 -6186 241634
rect -6806 205954 -6186 241398
rect -6806 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 -6186 205954
rect -6806 205634 -6186 205718
rect -6806 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 -6186 205634
rect -6806 169954 -6186 205398
rect -6806 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 -6186 169954
rect -6806 169634 -6186 169718
rect -6806 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 -6186 169634
rect -6806 133954 -6186 169398
rect -6806 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 -6186 133954
rect -6806 133634 -6186 133718
rect -6806 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 -6186 133634
rect -6806 97954 -6186 133398
rect -6806 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 -6186 97954
rect -6806 97634 -6186 97718
rect -6806 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 -6186 97634
rect -6806 61954 -6186 97398
rect -6806 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 -6186 61954
rect -6806 61634 -6186 61718
rect -6806 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 -6186 61634
rect -6806 25954 -6186 61398
rect -6806 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 -6186 25954
rect -6806 25634 -6186 25718
rect -6806 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 -6186 25634
rect -6806 -5146 -6186 25398
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 669454 -5226 708122
rect -5846 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 -5226 669454
rect -5846 669134 -5226 669218
rect -5846 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 -5226 669134
rect -5846 633454 -5226 668898
rect -5846 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 -5226 633454
rect -5846 633134 -5226 633218
rect -5846 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 -5226 633134
rect -5846 597454 -5226 632898
rect -5846 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 -5226 597454
rect -5846 597134 -5226 597218
rect -5846 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 -5226 597134
rect -5846 561454 -5226 596898
rect -5846 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 -5226 561454
rect -5846 561134 -5226 561218
rect -5846 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 -5226 561134
rect -5846 525454 -5226 560898
rect -5846 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 -5226 525454
rect -5846 525134 -5226 525218
rect -5846 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 -5226 525134
rect -5846 489454 -5226 524898
rect -5846 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 -5226 489454
rect -5846 489134 -5226 489218
rect -5846 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 -5226 489134
rect -5846 453454 -5226 488898
rect -5846 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 -5226 453454
rect -5846 453134 -5226 453218
rect -5846 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 -5226 453134
rect -5846 417454 -5226 452898
rect -5846 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 -5226 417454
rect -5846 417134 -5226 417218
rect -5846 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 -5226 417134
rect -5846 381454 -5226 416898
rect -5846 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 -5226 381454
rect -5846 381134 -5226 381218
rect -5846 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 -5226 381134
rect -5846 345454 -5226 380898
rect -5846 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 -5226 345454
rect -5846 345134 -5226 345218
rect -5846 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 -5226 345134
rect -5846 309454 -5226 344898
rect -5846 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 -5226 309454
rect -5846 309134 -5226 309218
rect -5846 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 -5226 309134
rect -5846 273454 -5226 308898
rect -5846 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 -5226 273454
rect -5846 273134 -5226 273218
rect -5846 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 -5226 273134
rect -5846 237454 -5226 272898
rect -5846 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 -5226 237454
rect -5846 237134 -5226 237218
rect -5846 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 -5226 237134
rect -5846 201454 -5226 236898
rect -5846 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 -5226 201454
rect -5846 201134 -5226 201218
rect -5846 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 -5226 201134
rect -5846 165454 -5226 200898
rect -5846 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 -5226 165454
rect -5846 165134 -5226 165218
rect -5846 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 -5226 165134
rect -5846 129454 -5226 164898
rect -5846 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 -5226 129454
rect -5846 129134 -5226 129218
rect -5846 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 -5226 129134
rect -5846 93454 -5226 128898
rect -5846 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 -5226 93454
rect -5846 93134 -5226 93218
rect -5846 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 -5226 93134
rect -5846 57454 -5226 92898
rect -5846 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 -5226 57454
rect -5846 57134 -5226 57218
rect -5846 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 -5226 57134
rect -5846 21454 -5226 56898
rect -5846 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 -5226 21454
rect -5846 21134 -5226 21218
rect -5846 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 -5226 21134
rect -5846 -4186 -5226 20898
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 700954 -4266 707162
rect -4886 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 -4266 700954
rect -4886 700634 -4266 700718
rect -4886 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 -4266 700634
rect -4886 664954 -4266 700398
rect -4886 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 -4266 664954
rect -4886 664634 -4266 664718
rect -4886 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 -4266 664634
rect -4886 628954 -4266 664398
rect -4886 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 -4266 628954
rect -4886 628634 -4266 628718
rect -4886 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 -4266 628634
rect -4886 592954 -4266 628398
rect -4886 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 -4266 592954
rect -4886 592634 -4266 592718
rect -4886 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 -4266 592634
rect -4886 556954 -4266 592398
rect -4886 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 -4266 556954
rect -4886 556634 -4266 556718
rect -4886 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 -4266 556634
rect -4886 520954 -4266 556398
rect -4886 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 -4266 520954
rect -4886 520634 -4266 520718
rect -4886 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 -4266 520634
rect -4886 484954 -4266 520398
rect -4886 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 -4266 484954
rect -4886 484634 -4266 484718
rect -4886 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 -4266 484634
rect -4886 448954 -4266 484398
rect -4886 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 -4266 448954
rect -4886 448634 -4266 448718
rect -4886 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 -4266 448634
rect -4886 412954 -4266 448398
rect -4886 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 -4266 412954
rect -4886 412634 -4266 412718
rect -4886 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 -4266 412634
rect -4886 376954 -4266 412398
rect -4886 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 -4266 376954
rect -4886 376634 -4266 376718
rect -4886 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 -4266 376634
rect -4886 340954 -4266 376398
rect -4886 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 -4266 340954
rect -4886 340634 -4266 340718
rect -4886 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 -4266 340634
rect -4886 304954 -4266 340398
rect -4886 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 -4266 304954
rect -4886 304634 -4266 304718
rect -4886 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 -4266 304634
rect -4886 268954 -4266 304398
rect -4886 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 -4266 268954
rect -4886 268634 -4266 268718
rect -4886 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 -4266 268634
rect -4886 232954 -4266 268398
rect -4886 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 -4266 232954
rect -4886 232634 -4266 232718
rect -4886 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 -4266 232634
rect -4886 196954 -4266 232398
rect -4886 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 -4266 196954
rect -4886 196634 -4266 196718
rect -4886 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 -4266 196634
rect -4886 160954 -4266 196398
rect -4886 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 -4266 160954
rect -4886 160634 -4266 160718
rect -4886 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 -4266 160634
rect -4886 124954 -4266 160398
rect -4886 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 -4266 124954
rect -4886 124634 -4266 124718
rect -4886 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 -4266 124634
rect -4886 88954 -4266 124398
rect -4886 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 -4266 88954
rect -4886 88634 -4266 88718
rect -4886 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 -4266 88634
rect -4886 52954 -4266 88398
rect -4886 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 -4266 52954
rect -4886 52634 -4266 52718
rect -4886 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 -4266 52634
rect -4886 16954 -4266 52398
rect -4886 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 -4266 16954
rect -4886 16634 -4266 16718
rect -4886 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 -4266 16634
rect -4886 -3226 -4266 16398
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 696454 -3306 706202
rect -3926 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 -3306 696454
rect -3926 696134 -3306 696218
rect -3926 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 -3306 696134
rect -3926 660454 -3306 695898
rect -3926 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 -3306 660454
rect -3926 660134 -3306 660218
rect -3926 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 -3306 660134
rect -3926 624454 -3306 659898
rect -3926 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 -3306 624454
rect -3926 624134 -3306 624218
rect -3926 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 -3306 624134
rect -3926 588454 -3306 623898
rect -3926 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 -3306 588454
rect -3926 588134 -3306 588218
rect -3926 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 -3306 588134
rect -3926 552454 -3306 587898
rect -3926 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 -3306 552454
rect -3926 552134 -3306 552218
rect -3926 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 -3306 552134
rect -3926 516454 -3306 551898
rect -3926 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 -3306 516454
rect -3926 516134 -3306 516218
rect -3926 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 -3306 516134
rect -3926 480454 -3306 515898
rect -3926 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 -3306 480454
rect -3926 480134 -3306 480218
rect -3926 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 -3306 480134
rect -3926 444454 -3306 479898
rect -3926 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 -3306 444454
rect -3926 444134 -3306 444218
rect -3926 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 -3306 444134
rect -3926 408454 -3306 443898
rect -3926 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 -3306 408454
rect -3926 408134 -3306 408218
rect -3926 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 -3306 408134
rect -3926 372454 -3306 407898
rect -3926 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 -3306 372454
rect -3926 372134 -3306 372218
rect -3926 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 -3306 372134
rect -3926 336454 -3306 371898
rect -3926 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 -3306 336454
rect -3926 336134 -3306 336218
rect -3926 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 -3306 336134
rect -3926 300454 -3306 335898
rect -3926 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 -3306 300454
rect -3926 300134 -3306 300218
rect -3926 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 -3306 300134
rect -3926 264454 -3306 299898
rect -3926 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 -3306 264454
rect -3926 264134 -3306 264218
rect -3926 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 -3306 264134
rect -3926 228454 -3306 263898
rect -3926 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 -3306 228454
rect -3926 228134 -3306 228218
rect -3926 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 -3306 228134
rect -3926 192454 -3306 227898
rect -3926 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 -3306 192454
rect -3926 192134 -3306 192218
rect -3926 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 -3306 192134
rect -3926 156454 -3306 191898
rect -3926 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 -3306 156454
rect -3926 156134 -3306 156218
rect -3926 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 -3306 156134
rect -3926 120454 -3306 155898
rect -3926 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 -3306 120454
rect -3926 120134 -3306 120218
rect -3926 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 -3306 120134
rect -3926 84454 -3306 119898
rect -3926 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 -3306 84454
rect -3926 84134 -3306 84218
rect -3926 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 -3306 84134
rect -3926 48454 -3306 83898
rect -3926 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 -3306 48454
rect -3926 48134 -3306 48218
rect -3926 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 -3306 48134
rect -3926 12454 -3306 47898
rect -3926 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 -3306 12454
rect -3926 12134 -3306 12218
rect -3926 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 -3306 12134
rect -3926 -2266 -3306 11898
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691954 -2346 705242
rect -2966 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 -2346 691954
rect -2966 691634 -2346 691718
rect -2966 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 -2346 691634
rect -2966 655954 -2346 691398
rect -2966 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 -2346 655954
rect -2966 655634 -2346 655718
rect -2966 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 -2346 655634
rect -2966 619954 -2346 655398
rect -2966 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 -2346 619954
rect -2966 619634 -2346 619718
rect -2966 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 -2346 619634
rect -2966 583954 -2346 619398
rect -2966 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 -2346 583954
rect -2966 583634 -2346 583718
rect -2966 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 -2346 583634
rect -2966 547954 -2346 583398
rect -2966 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 -2346 547954
rect -2966 547634 -2346 547718
rect -2966 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 -2346 547634
rect -2966 511954 -2346 547398
rect -2966 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 -2346 511954
rect -2966 511634 -2346 511718
rect -2966 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 -2346 511634
rect -2966 475954 -2346 511398
rect -2966 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 -2346 475954
rect -2966 475634 -2346 475718
rect -2966 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 -2346 475634
rect -2966 439954 -2346 475398
rect -2966 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 -2346 439954
rect -2966 439634 -2346 439718
rect -2966 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 -2346 439634
rect -2966 403954 -2346 439398
rect -2966 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 -2346 403954
rect -2966 403634 -2346 403718
rect -2966 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 -2346 403634
rect -2966 367954 -2346 403398
rect -2966 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 -2346 367954
rect -2966 367634 -2346 367718
rect -2966 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 -2346 367634
rect -2966 331954 -2346 367398
rect -2966 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 -2346 331954
rect -2966 331634 -2346 331718
rect -2966 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 -2346 331634
rect -2966 295954 -2346 331398
rect -2966 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 -2346 295954
rect -2966 295634 -2346 295718
rect -2966 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 -2346 295634
rect -2966 259954 -2346 295398
rect -2966 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 -2346 259954
rect -2966 259634 -2346 259718
rect -2966 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 -2346 259634
rect -2966 223954 -2346 259398
rect -2966 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 -2346 223954
rect -2966 223634 -2346 223718
rect -2966 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 -2346 223634
rect -2966 187954 -2346 223398
rect -2966 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 -2346 187954
rect -2966 187634 -2346 187718
rect -2966 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 -2346 187634
rect -2966 151954 -2346 187398
rect -2966 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 -2346 151954
rect -2966 151634 -2346 151718
rect -2966 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 -2346 151634
rect -2966 115954 -2346 151398
rect -2966 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 -2346 115954
rect -2966 115634 -2346 115718
rect -2966 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 -2346 115634
rect -2966 79954 -2346 115398
rect -2966 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 -2346 79954
rect -2966 79634 -2346 79718
rect -2966 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 -2346 79634
rect -2966 43954 -2346 79398
rect -2966 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 -2346 43954
rect -2966 43634 -2346 43718
rect -2966 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 -2346 43634
rect -2966 7954 -2346 43398
rect -2966 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 -2346 7954
rect -2966 7634 -2346 7718
rect -2966 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 -2346 7634
rect -2966 -1306 -2346 7398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 6294 705798 6914 711590
rect 6294 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 6914 705798
rect 6294 705478 6914 705562
rect 6294 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 6914 705478
rect 6294 691954 6914 705242
rect 6294 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 6914 691954
rect 6294 691634 6914 691718
rect 6294 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 6914 691634
rect 6294 655954 6914 691398
rect 6294 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 6914 655954
rect 6294 655634 6914 655718
rect 6294 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 6914 655634
rect 6294 619954 6914 655398
rect 6294 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 6914 619954
rect 6294 619634 6914 619718
rect 6294 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 6914 619634
rect 6294 583954 6914 619398
rect 6294 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 6914 583954
rect 6294 583634 6914 583718
rect 6294 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 6914 583634
rect 6294 547954 6914 583398
rect 6294 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 6914 547954
rect 6294 547634 6914 547718
rect 6294 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 6914 547634
rect 6294 511954 6914 547398
rect 6294 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 6914 511954
rect 6294 511634 6914 511718
rect 6294 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 6914 511634
rect 6294 475954 6914 511398
rect 6294 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 6914 475954
rect 6294 475634 6914 475718
rect 6294 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 6914 475634
rect 6294 439954 6914 475398
rect 6294 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 6914 439954
rect 6294 439634 6914 439718
rect 6294 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 6914 439634
rect 6294 403954 6914 439398
rect 6294 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 6914 403954
rect 6294 403634 6914 403718
rect 6294 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 6914 403634
rect 6294 367954 6914 403398
rect 6294 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 6914 367954
rect 6294 367634 6914 367718
rect 6294 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 6914 367634
rect 6294 331954 6914 367398
rect 6294 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 6914 331954
rect 6294 331634 6914 331718
rect 6294 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 6914 331634
rect 6294 295954 6914 331398
rect 6294 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 6914 295954
rect 6294 295634 6914 295718
rect 6294 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 6914 295634
rect 6294 259954 6914 295398
rect 6294 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 6914 259954
rect 6294 259634 6914 259718
rect 6294 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 6914 259634
rect 6294 223954 6914 259398
rect 6294 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 6914 223954
rect 6294 223634 6914 223718
rect 6294 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 6914 223634
rect 6294 187954 6914 223398
rect 6294 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 6914 187954
rect 6294 187634 6914 187718
rect 6294 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 6914 187634
rect 6294 151954 6914 187398
rect 6294 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 6914 151954
rect 6294 151634 6914 151718
rect 6294 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 6914 151634
rect 6294 115954 6914 151398
rect 6294 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 6914 115954
rect 6294 115634 6914 115718
rect 6294 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 6914 115634
rect 6294 79954 6914 115398
rect 6294 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 6914 79954
rect 6294 79634 6914 79718
rect 6294 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 6914 79634
rect 6294 43954 6914 79398
rect 6294 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 6914 43954
rect 6294 43634 6914 43718
rect 6294 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 6914 43634
rect 6294 7954 6914 43398
rect 6294 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 6914 7954
rect 6294 7634 6914 7718
rect 6294 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 6914 7634
rect 6294 -1306 6914 7398
rect 6294 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 6914 -1306
rect 6294 -1626 6914 -1542
rect 6294 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 6914 -1626
rect 6294 -7654 6914 -1862
rect 10794 706758 11414 711590
rect 10794 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 11414 706758
rect 10794 706438 11414 706522
rect 10794 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 11414 706438
rect 10794 696454 11414 706202
rect 10794 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 11414 696454
rect 10794 696134 11414 696218
rect 10794 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 11414 696134
rect 10794 660454 11414 695898
rect 10794 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 11414 660454
rect 10794 660134 11414 660218
rect 10794 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 11414 660134
rect 10794 624454 11414 659898
rect 10794 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 11414 624454
rect 10794 624134 11414 624218
rect 10794 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 11414 624134
rect 10794 588454 11414 623898
rect 10794 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 11414 588454
rect 10794 588134 11414 588218
rect 10794 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 11414 588134
rect 10794 552454 11414 587898
rect 10794 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 11414 552454
rect 10794 552134 11414 552218
rect 10794 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 11414 552134
rect 10794 516454 11414 551898
rect 10794 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 11414 516454
rect 10794 516134 11414 516218
rect 10794 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 11414 516134
rect 10794 480454 11414 515898
rect 10794 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 11414 480454
rect 10794 480134 11414 480218
rect 10794 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 11414 480134
rect 10794 444454 11414 479898
rect 10794 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 11414 444454
rect 10794 444134 11414 444218
rect 10794 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 11414 444134
rect 10794 408454 11414 443898
rect 10794 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 11414 408454
rect 10794 408134 11414 408218
rect 10794 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 11414 408134
rect 10794 372454 11414 407898
rect 10794 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 11414 372454
rect 10794 372134 11414 372218
rect 10794 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 11414 372134
rect 10794 336454 11414 371898
rect 10794 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 11414 336454
rect 10794 336134 11414 336218
rect 10794 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 11414 336134
rect 10794 300454 11414 335898
rect 10794 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 11414 300454
rect 10794 300134 11414 300218
rect 10794 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 11414 300134
rect 10794 264454 11414 299898
rect 10794 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 11414 264454
rect 10794 264134 11414 264218
rect 10794 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 11414 264134
rect 10794 228454 11414 263898
rect 10794 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 11414 228454
rect 10794 228134 11414 228218
rect 10794 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 11414 228134
rect 10794 192454 11414 227898
rect 10794 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 11414 192454
rect 10794 192134 11414 192218
rect 10794 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 11414 192134
rect 10794 156454 11414 191898
rect 10794 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 11414 156454
rect 10794 156134 11414 156218
rect 10794 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 11414 156134
rect 10794 120454 11414 155898
rect 10794 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 11414 120454
rect 10794 120134 11414 120218
rect 10794 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 11414 120134
rect 10794 84454 11414 119898
rect 10794 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 11414 84454
rect 10794 84134 11414 84218
rect 10794 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 11414 84134
rect 10794 48454 11414 83898
rect 10794 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 11414 48454
rect 10794 48134 11414 48218
rect 10794 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 11414 48134
rect 10794 12454 11414 47898
rect 10794 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 11414 12454
rect 10794 12134 11414 12218
rect 10794 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 11414 12134
rect 10794 -2266 11414 11898
rect 10794 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 11414 -2266
rect 10794 -2586 11414 -2502
rect 10794 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 11414 -2586
rect 10794 -7654 11414 -2822
rect 15294 707718 15914 711590
rect 15294 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 15914 707718
rect 15294 707398 15914 707482
rect 15294 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 15914 707398
rect 15294 700954 15914 707162
rect 15294 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 15914 700954
rect 15294 700634 15914 700718
rect 15294 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 15914 700634
rect 15294 664954 15914 700398
rect 15294 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 15914 664954
rect 15294 664634 15914 664718
rect 15294 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 15914 664634
rect 15294 628954 15914 664398
rect 15294 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 15914 628954
rect 15294 628634 15914 628718
rect 15294 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 15914 628634
rect 15294 592954 15914 628398
rect 15294 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 15914 592954
rect 15294 592634 15914 592718
rect 15294 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 15914 592634
rect 15294 556954 15914 592398
rect 15294 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 15914 556954
rect 15294 556634 15914 556718
rect 15294 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 15914 556634
rect 15294 520954 15914 556398
rect 15294 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 15914 520954
rect 15294 520634 15914 520718
rect 15294 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 15914 520634
rect 15294 484954 15914 520398
rect 15294 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 15914 484954
rect 15294 484634 15914 484718
rect 15294 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 15914 484634
rect 15294 448954 15914 484398
rect 15294 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 15914 448954
rect 15294 448634 15914 448718
rect 15294 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 15914 448634
rect 15294 412954 15914 448398
rect 15294 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 15914 412954
rect 15294 412634 15914 412718
rect 15294 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 15914 412634
rect 15294 376954 15914 412398
rect 15294 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 15914 376954
rect 15294 376634 15914 376718
rect 15294 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 15914 376634
rect 15294 340954 15914 376398
rect 15294 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 15914 340954
rect 15294 340634 15914 340718
rect 15294 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 15914 340634
rect 15294 304954 15914 340398
rect 15294 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 15914 304954
rect 15294 304634 15914 304718
rect 15294 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 15914 304634
rect 15294 268954 15914 304398
rect 15294 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 15914 268954
rect 15294 268634 15914 268718
rect 15294 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 15914 268634
rect 15294 232954 15914 268398
rect 15294 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 15914 232954
rect 15294 232634 15914 232718
rect 15294 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 15914 232634
rect 15294 196954 15914 232398
rect 15294 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 15914 196954
rect 15294 196634 15914 196718
rect 15294 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 15914 196634
rect 15294 160954 15914 196398
rect 15294 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 15914 160954
rect 15294 160634 15914 160718
rect 15294 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 15914 160634
rect 15294 124954 15914 160398
rect 15294 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 15914 124954
rect 15294 124634 15914 124718
rect 15294 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 15914 124634
rect 15294 88954 15914 124398
rect 15294 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 15914 88954
rect 15294 88634 15914 88718
rect 15294 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 15914 88634
rect 15294 52954 15914 88398
rect 15294 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 15914 52954
rect 15294 52634 15914 52718
rect 15294 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 15914 52634
rect 15294 16954 15914 52398
rect 15294 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 15914 16954
rect 15294 16634 15914 16718
rect 15294 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 15914 16634
rect 15294 -3226 15914 16398
rect 15294 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 15914 -3226
rect 15294 -3546 15914 -3462
rect 15294 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 15914 -3546
rect 15294 -7654 15914 -3782
rect 19794 708678 20414 711590
rect 19794 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 20414 708678
rect 19794 708358 20414 708442
rect 19794 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 20414 708358
rect 19794 669454 20414 708122
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -4186 20414 20898
rect 19794 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 20414 -4186
rect 19794 -4506 20414 -4422
rect 19794 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 20414 -4506
rect 19794 -7654 20414 -4742
rect 24294 709638 24914 711590
rect 24294 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 24914 709638
rect 24294 709318 24914 709402
rect 24294 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 24914 709318
rect 24294 673954 24914 709082
rect 24294 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 24914 673954
rect 24294 673634 24914 673718
rect 24294 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 24914 673634
rect 24294 637954 24914 673398
rect 24294 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 24914 637954
rect 24294 637634 24914 637718
rect 24294 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 24914 637634
rect 24294 601954 24914 637398
rect 24294 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 24914 601954
rect 24294 601634 24914 601718
rect 24294 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 24914 601634
rect 24294 565954 24914 601398
rect 24294 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 24914 565954
rect 24294 565634 24914 565718
rect 24294 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 24914 565634
rect 24294 529954 24914 565398
rect 24294 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 24914 529954
rect 24294 529634 24914 529718
rect 24294 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 24914 529634
rect 24294 493954 24914 529398
rect 24294 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 24914 493954
rect 24294 493634 24914 493718
rect 24294 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 24914 493634
rect 24294 457954 24914 493398
rect 24294 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 24914 457954
rect 24294 457634 24914 457718
rect 24294 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 24914 457634
rect 24294 421954 24914 457398
rect 24294 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 24914 421954
rect 24294 421634 24914 421718
rect 24294 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 24914 421634
rect 24294 385954 24914 421398
rect 24294 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 24914 385954
rect 24294 385634 24914 385718
rect 24294 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 24914 385634
rect 24294 349954 24914 385398
rect 24294 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 24914 349954
rect 24294 349634 24914 349718
rect 24294 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 24914 349634
rect 24294 313954 24914 349398
rect 24294 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 24914 313954
rect 24294 313634 24914 313718
rect 24294 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 24914 313634
rect 24294 277954 24914 313398
rect 24294 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 24914 277954
rect 24294 277634 24914 277718
rect 24294 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 24914 277634
rect 24294 241954 24914 277398
rect 24294 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 24914 241954
rect 24294 241634 24914 241718
rect 24294 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 24914 241634
rect 24294 205954 24914 241398
rect 24294 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 24914 205954
rect 24294 205634 24914 205718
rect 24294 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 24914 205634
rect 24294 169954 24914 205398
rect 24294 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 24914 169954
rect 24294 169634 24914 169718
rect 24294 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 24914 169634
rect 24294 133954 24914 169398
rect 24294 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 24914 133954
rect 24294 133634 24914 133718
rect 24294 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 24914 133634
rect 24294 97954 24914 133398
rect 24294 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 24914 97954
rect 24294 97634 24914 97718
rect 24294 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 24914 97634
rect 24294 61954 24914 97398
rect 24294 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 24914 61954
rect 24294 61634 24914 61718
rect 24294 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 24914 61634
rect 24294 25954 24914 61398
rect 24294 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 24914 25954
rect 24294 25634 24914 25718
rect 24294 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 24914 25634
rect 24294 -5146 24914 25398
rect 24294 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 24914 -5146
rect 24294 -5466 24914 -5382
rect 24294 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 24914 -5466
rect 24294 -7654 24914 -5702
rect 28794 710598 29414 711590
rect 28794 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 29414 710598
rect 28794 710278 29414 710362
rect 28794 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 29414 710278
rect 28794 678454 29414 710042
rect 28794 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 29414 678454
rect 28794 678134 29414 678218
rect 28794 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 29414 678134
rect 28794 642454 29414 677898
rect 28794 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642218 29414 642454
rect 28794 642134 29414 642218
rect 28794 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 641898 29414 642134
rect 28794 606454 29414 641898
rect 28794 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 29414 606454
rect 28794 606134 29414 606218
rect 28794 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 29414 606134
rect 28794 570454 29414 605898
rect 28794 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 29414 570454
rect 28794 570134 29414 570218
rect 28794 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 29414 570134
rect 28794 534454 29414 569898
rect 28794 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 29414 534454
rect 28794 534134 29414 534218
rect 28794 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 29414 534134
rect 28794 498454 29414 533898
rect 28794 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 29414 498454
rect 28794 498134 29414 498218
rect 28794 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 29414 498134
rect 28794 462454 29414 497898
rect 28794 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 29414 462454
rect 28794 462134 29414 462218
rect 28794 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 29414 462134
rect 28794 426454 29414 461898
rect 28794 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 29414 426454
rect 28794 426134 29414 426218
rect 28794 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 29414 426134
rect 28794 390454 29414 425898
rect 28794 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 29414 390454
rect 28794 390134 29414 390218
rect 28794 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 29414 390134
rect 28794 354454 29414 389898
rect 28794 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 29414 354454
rect 28794 354134 29414 354218
rect 28794 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 29414 354134
rect 28794 318454 29414 353898
rect 28794 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 29414 318454
rect 28794 318134 29414 318218
rect 28794 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 29414 318134
rect 28794 282454 29414 317898
rect 28794 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 29414 282454
rect 28794 282134 29414 282218
rect 28794 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 29414 282134
rect 28794 246454 29414 281898
rect 28794 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 29414 246454
rect 28794 246134 29414 246218
rect 28794 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 29414 246134
rect 28794 210454 29414 245898
rect 28794 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 29414 210454
rect 28794 210134 29414 210218
rect 28794 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 29414 210134
rect 28794 174454 29414 209898
rect 28794 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 29414 174454
rect 28794 174134 29414 174218
rect 28794 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 29414 174134
rect 28794 138454 29414 173898
rect 28794 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 29414 138454
rect 28794 138134 29414 138218
rect 28794 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 29414 138134
rect 28794 102454 29414 137898
rect 28794 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 29414 102454
rect 28794 102134 29414 102218
rect 28794 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 29414 102134
rect 28794 66454 29414 101898
rect 28794 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 29414 66454
rect 28794 66134 29414 66218
rect 28794 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 29414 66134
rect 28794 30454 29414 65898
rect 28794 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 29414 30454
rect 28794 30134 29414 30218
rect 28794 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 29414 30134
rect 28794 -6106 29414 29898
rect 28794 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 29414 -6106
rect 28794 -6426 29414 -6342
rect 28794 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 29414 -6426
rect 28794 -7654 29414 -6662
rect 33294 711558 33914 711590
rect 33294 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 33914 711558
rect 33294 711238 33914 711322
rect 33294 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 33914 711238
rect 33294 682954 33914 711002
rect 33294 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 33914 682954
rect 33294 682634 33914 682718
rect 33294 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 33914 682634
rect 33294 646954 33914 682398
rect 33294 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 33914 646954
rect 33294 646634 33914 646718
rect 33294 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 33914 646634
rect 33294 610954 33914 646398
rect 33294 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 33914 610954
rect 33294 610634 33914 610718
rect 33294 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 33914 610634
rect 33294 574954 33914 610398
rect 33294 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 33914 574954
rect 33294 574634 33914 574718
rect 33294 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 33914 574634
rect 33294 538954 33914 574398
rect 33294 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 33914 538954
rect 33294 538634 33914 538718
rect 33294 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 33914 538634
rect 33294 502954 33914 538398
rect 33294 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 33914 502954
rect 33294 502634 33914 502718
rect 33294 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 33914 502634
rect 33294 466954 33914 502398
rect 33294 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 33914 466954
rect 33294 466634 33914 466718
rect 33294 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 33914 466634
rect 33294 430954 33914 466398
rect 33294 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 33914 430954
rect 33294 430634 33914 430718
rect 33294 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 33914 430634
rect 33294 394954 33914 430398
rect 33294 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 33914 394954
rect 33294 394634 33914 394718
rect 33294 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 33914 394634
rect 33294 358954 33914 394398
rect 33294 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 33914 358954
rect 33294 358634 33914 358718
rect 33294 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 33914 358634
rect 33294 322954 33914 358398
rect 33294 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 33914 322954
rect 33294 322634 33914 322718
rect 33294 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 33914 322634
rect 33294 286954 33914 322398
rect 33294 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 33914 286954
rect 33294 286634 33914 286718
rect 33294 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 33914 286634
rect 33294 250954 33914 286398
rect 33294 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 33914 250954
rect 33294 250634 33914 250718
rect 33294 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 33914 250634
rect 33294 214954 33914 250398
rect 33294 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 33914 214954
rect 33294 214634 33914 214718
rect 33294 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 33914 214634
rect 33294 178954 33914 214398
rect 33294 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 33914 178954
rect 33294 178634 33914 178718
rect 33294 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 33914 178634
rect 33294 142954 33914 178398
rect 33294 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 33914 142954
rect 33294 142634 33914 142718
rect 33294 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 33914 142634
rect 33294 106954 33914 142398
rect 33294 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 33914 106954
rect 33294 106634 33914 106718
rect 33294 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 33914 106634
rect 33294 70954 33914 106398
rect 33294 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 33914 70954
rect 33294 70634 33914 70718
rect 33294 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 33914 70634
rect 33294 34954 33914 70398
rect 33294 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 33914 34954
rect 33294 34634 33914 34718
rect 33294 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 33914 34634
rect 33294 -7066 33914 34398
rect 33294 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 33914 -7066
rect 33294 -7386 33914 -7302
rect 33294 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 33914 -7386
rect 33294 -7654 33914 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 42294 705798 42914 711590
rect 42294 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 42914 705798
rect 42294 705478 42914 705562
rect 42294 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 42914 705478
rect 42294 691954 42914 705242
rect 42294 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 42914 691954
rect 42294 691634 42914 691718
rect 42294 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 42914 691634
rect 42294 655954 42914 691398
rect 42294 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 42914 655954
rect 42294 655634 42914 655718
rect 42294 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 42914 655634
rect 42294 619954 42914 655398
rect 42294 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 42914 619954
rect 42294 619634 42914 619718
rect 42294 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 42914 619634
rect 42294 583954 42914 619398
rect 42294 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 42914 583954
rect 42294 583634 42914 583718
rect 42294 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 42914 583634
rect 42294 547954 42914 583398
rect 42294 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 42914 547954
rect 42294 547634 42914 547718
rect 42294 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 42914 547634
rect 42294 511954 42914 547398
rect 42294 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 42914 511954
rect 42294 511634 42914 511718
rect 42294 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 42914 511634
rect 42294 475954 42914 511398
rect 42294 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 42914 475954
rect 42294 475634 42914 475718
rect 42294 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 42914 475634
rect 42294 439954 42914 475398
rect 42294 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 42914 439954
rect 42294 439634 42914 439718
rect 42294 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 42914 439634
rect 42294 403954 42914 439398
rect 42294 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 42914 403954
rect 42294 403634 42914 403718
rect 42294 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 42914 403634
rect 42294 367954 42914 403398
rect 42294 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 42914 367954
rect 42294 367634 42914 367718
rect 42294 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 42914 367634
rect 42294 331954 42914 367398
rect 42294 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 42914 331954
rect 42294 331634 42914 331718
rect 42294 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 42914 331634
rect 42294 295954 42914 331398
rect 42294 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 42914 295954
rect 42294 295634 42914 295718
rect 42294 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 42914 295634
rect 42294 259954 42914 295398
rect 42294 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 42914 259954
rect 42294 259634 42914 259718
rect 42294 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 42914 259634
rect 42294 223954 42914 259398
rect 42294 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 42914 223954
rect 42294 223634 42914 223718
rect 42294 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 42914 223634
rect 42294 187954 42914 223398
rect 42294 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 42914 187954
rect 42294 187634 42914 187718
rect 42294 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 42914 187634
rect 42294 151954 42914 187398
rect 42294 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 42914 151954
rect 42294 151634 42914 151718
rect 42294 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 42914 151634
rect 42294 115954 42914 151398
rect 42294 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 42914 115954
rect 42294 115634 42914 115718
rect 42294 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 42914 115634
rect 42294 79954 42914 115398
rect 42294 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 42914 79954
rect 42294 79634 42914 79718
rect 42294 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 42914 79634
rect 42294 43954 42914 79398
rect 42294 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 42914 43954
rect 42294 43634 42914 43718
rect 42294 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 42914 43634
rect 42294 7954 42914 43398
rect 42294 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 42914 7954
rect 42294 7634 42914 7718
rect 42294 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 42914 7634
rect 42294 -1306 42914 7398
rect 42294 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 42914 -1306
rect 42294 -1626 42914 -1542
rect 42294 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 42914 -1626
rect 42294 -7654 42914 -1862
rect 46794 706758 47414 711590
rect 46794 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 47414 706758
rect 46794 706438 47414 706522
rect 46794 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 47414 706438
rect 46794 696454 47414 706202
rect 46794 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 47414 696454
rect 46794 696134 47414 696218
rect 46794 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 47414 696134
rect 46794 660454 47414 695898
rect 51294 707718 51914 711590
rect 51294 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 51914 707718
rect 51294 707398 51914 707482
rect 51294 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 51914 707398
rect 51294 700954 51914 707162
rect 51294 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 51914 700954
rect 51294 700634 51914 700718
rect 51294 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 51914 700634
rect 51294 664954 51914 700398
rect 51294 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 51914 664954
rect 51294 664634 51914 664718
rect 51294 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 51914 664634
rect 51294 664000 51914 664398
rect 55794 708678 56414 711590
rect 55794 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 56414 708678
rect 55794 708358 56414 708442
rect 55794 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 56414 708358
rect 55794 669454 56414 708122
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 664000 56414 668898
rect 60294 709638 60914 711590
rect 60294 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 60914 709638
rect 60294 709318 60914 709402
rect 60294 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 60914 709318
rect 60294 673954 60914 709082
rect 60294 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 60914 673954
rect 60294 673634 60914 673718
rect 60294 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 60914 673634
rect 60294 664000 60914 673398
rect 64794 710598 65414 711590
rect 64794 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 65414 710598
rect 64794 710278 65414 710362
rect 64794 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 65414 710278
rect 64794 678454 65414 710042
rect 64794 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 65414 678454
rect 64794 678134 65414 678218
rect 64794 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 65414 678134
rect 64794 664000 65414 677898
rect 69294 711558 69914 711590
rect 69294 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 69914 711558
rect 69294 711238 69914 711322
rect 69294 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 69914 711238
rect 69294 682954 69914 711002
rect 69294 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 69914 682954
rect 69294 682634 69914 682718
rect 69294 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 69914 682634
rect 69294 664000 69914 682398
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 664000 74414 686898
rect 78294 705798 78914 711590
rect 78294 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 78914 705798
rect 78294 705478 78914 705562
rect 78294 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 78914 705478
rect 78294 691954 78914 705242
rect 78294 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 78914 691954
rect 78294 691634 78914 691718
rect 78294 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 78914 691634
rect 78294 664000 78914 691398
rect 82794 706758 83414 711590
rect 82794 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 83414 706758
rect 82794 706438 83414 706522
rect 82794 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 83414 706438
rect 82794 696454 83414 706202
rect 82794 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 83414 696454
rect 82794 696134 83414 696218
rect 82794 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 83414 696134
rect 82794 664000 83414 695898
rect 87294 707718 87914 711590
rect 87294 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 87914 707718
rect 87294 707398 87914 707482
rect 87294 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 87914 707398
rect 87294 700954 87914 707162
rect 87294 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 87914 700954
rect 87294 700634 87914 700718
rect 87294 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 87914 700634
rect 87294 664954 87914 700398
rect 87294 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 87914 664954
rect 87294 664634 87914 664718
rect 87294 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 87914 664634
rect 87294 664000 87914 664398
rect 91794 708678 92414 711590
rect 91794 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 92414 708678
rect 91794 708358 92414 708442
rect 91794 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 92414 708358
rect 91794 669454 92414 708122
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 664000 92414 668898
rect 96294 709638 96914 711590
rect 96294 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 96914 709638
rect 96294 709318 96914 709402
rect 96294 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 96914 709318
rect 96294 673954 96914 709082
rect 96294 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 96914 673954
rect 96294 673634 96914 673718
rect 96294 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 96914 673634
rect 96294 664000 96914 673398
rect 100794 710598 101414 711590
rect 100794 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 101414 710598
rect 100794 710278 101414 710362
rect 100794 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 101414 710278
rect 100794 678454 101414 710042
rect 100794 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 101414 678454
rect 100794 678134 101414 678218
rect 100794 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 101414 678134
rect 100794 664000 101414 677898
rect 105294 711558 105914 711590
rect 105294 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 105914 711558
rect 105294 711238 105914 711322
rect 105294 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 105914 711238
rect 105294 682954 105914 711002
rect 105294 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 105914 682954
rect 105294 682634 105914 682718
rect 105294 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 105914 682634
rect 105294 664000 105914 682398
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 664000 110414 686898
rect 114294 705798 114914 711590
rect 114294 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 114914 705798
rect 114294 705478 114914 705562
rect 114294 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 114914 705478
rect 114294 691954 114914 705242
rect 114294 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 114914 691954
rect 114294 691634 114914 691718
rect 114294 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 114914 691634
rect 114294 664000 114914 691398
rect 118794 706758 119414 711590
rect 118794 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 119414 706758
rect 118794 706438 119414 706522
rect 118794 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 119414 706438
rect 118794 696454 119414 706202
rect 118794 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 119414 696454
rect 118794 696134 119414 696218
rect 118794 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 119414 696134
rect 118794 664000 119414 695898
rect 123294 707718 123914 711590
rect 123294 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 123914 707718
rect 123294 707398 123914 707482
rect 123294 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 123914 707398
rect 123294 700954 123914 707162
rect 123294 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 123914 700954
rect 123294 700634 123914 700718
rect 123294 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 123914 700634
rect 123294 664954 123914 700398
rect 123294 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 123914 664954
rect 123294 664634 123914 664718
rect 123294 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 123914 664634
rect 123294 664000 123914 664398
rect 127794 708678 128414 711590
rect 127794 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 128414 708678
rect 127794 708358 128414 708442
rect 127794 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 128414 708358
rect 127794 669454 128414 708122
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 664000 128414 668898
rect 132294 709638 132914 711590
rect 132294 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 132914 709638
rect 132294 709318 132914 709402
rect 132294 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 132914 709318
rect 132294 673954 132914 709082
rect 132294 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 132914 673954
rect 132294 673634 132914 673718
rect 132294 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 132914 673634
rect 132294 664000 132914 673398
rect 136794 710598 137414 711590
rect 136794 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 137414 710598
rect 136794 710278 137414 710362
rect 136794 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 137414 710278
rect 136794 678454 137414 710042
rect 136794 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 137414 678454
rect 136794 678134 137414 678218
rect 136794 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 137414 678134
rect 136794 664000 137414 677898
rect 141294 711558 141914 711590
rect 141294 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 141914 711558
rect 141294 711238 141914 711322
rect 141294 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 141914 711238
rect 141294 682954 141914 711002
rect 141294 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 141914 682954
rect 141294 682634 141914 682718
rect 141294 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 141914 682634
rect 141294 664000 141914 682398
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 664000 146414 686898
rect 150294 705798 150914 711590
rect 150294 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 150914 705798
rect 150294 705478 150914 705562
rect 150294 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 150914 705478
rect 150294 691954 150914 705242
rect 150294 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 150914 691954
rect 150294 691634 150914 691718
rect 150294 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 150914 691634
rect 150294 664000 150914 691398
rect 154794 706758 155414 711590
rect 154794 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 155414 706758
rect 154794 706438 155414 706522
rect 154794 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 155414 706438
rect 154794 696454 155414 706202
rect 154794 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 155414 696454
rect 154794 696134 155414 696218
rect 154794 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 155414 696134
rect 154794 664000 155414 695898
rect 159294 707718 159914 711590
rect 159294 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 159914 707718
rect 159294 707398 159914 707482
rect 159294 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 159914 707398
rect 159294 700954 159914 707162
rect 159294 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 159914 700954
rect 159294 700634 159914 700718
rect 159294 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 159914 700634
rect 159294 664954 159914 700398
rect 159294 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 159914 664954
rect 159294 664634 159914 664718
rect 159294 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 159914 664634
rect 159294 664000 159914 664398
rect 163794 708678 164414 711590
rect 163794 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 164414 708678
rect 163794 708358 164414 708442
rect 163794 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 164414 708358
rect 163794 669454 164414 708122
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 664000 164414 668898
rect 168294 709638 168914 711590
rect 168294 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 168914 709638
rect 168294 709318 168914 709402
rect 168294 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 168914 709318
rect 168294 673954 168914 709082
rect 168294 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 168914 673954
rect 168294 673634 168914 673718
rect 168294 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 168914 673634
rect 168294 664000 168914 673398
rect 172794 710598 173414 711590
rect 172794 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 173414 710598
rect 172794 710278 173414 710362
rect 172794 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 173414 710278
rect 172794 678454 173414 710042
rect 172794 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 173414 678454
rect 172794 678134 173414 678218
rect 172794 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 173414 678134
rect 172794 664000 173414 677898
rect 177294 711558 177914 711590
rect 177294 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 177914 711558
rect 177294 711238 177914 711322
rect 177294 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 177914 711238
rect 177294 682954 177914 711002
rect 177294 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 177914 682954
rect 177294 682634 177914 682718
rect 177294 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 177914 682634
rect 177294 664000 177914 682398
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 664000 182414 686898
rect 186294 705798 186914 711590
rect 186294 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 186914 705798
rect 186294 705478 186914 705562
rect 186294 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 186914 705478
rect 186294 691954 186914 705242
rect 186294 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 186914 691954
rect 186294 691634 186914 691718
rect 186294 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 186914 691634
rect 186294 664000 186914 691398
rect 190794 706758 191414 711590
rect 190794 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 191414 706758
rect 190794 706438 191414 706522
rect 190794 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 191414 706438
rect 190794 696454 191414 706202
rect 190794 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 191414 696454
rect 190794 696134 191414 696218
rect 190794 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 191414 696134
rect 190794 664000 191414 695898
rect 195294 707718 195914 711590
rect 195294 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 195914 707718
rect 195294 707398 195914 707482
rect 195294 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 195914 707398
rect 195294 700954 195914 707162
rect 195294 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 195914 700954
rect 195294 700634 195914 700718
rect 195294 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 195914 700634
rect 195294 664954 195914 700398
rect 195294 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 195914 664954
rect 195294 664634 195914 664718
rect 195294 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 195914 664634
rect 195294 664000 195914 664398
rect 199794 708678 200414 711590
rect 199794 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 200414 708678
rect 199794 708358 200414 708442
rect 199794 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 200414 708358
rect 199794 669454 200414 708122
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 664000 200414 668898
rect 204294 709638 204914 711590
rect 204294 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 204914 709638
rect 204294 709318 204914 709402
rect 204294 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 204914 709318
rect 204294 673954 204914 709082
rect 204294 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 204914 673954
rect 204294 673634 204914 673718
rect 204294 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 204914 673634
rect 204294 664000 204914 673398
rect 208794 710598 209414 711590
rect 208794 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 209414 710598
rect 208794 710278 209414 710362
rect 208794 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 209414 710278
rect 208794 678454 209414 710042
rect 208794 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 209414 678454
rect 208794 678134 209414 678218
rect 208794 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 209414 678134
rect 208794 664000 209414 677898
rect 213294 711558 213914 711590
rect 213294 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 213914 711558
rect 213294 711238 213914 711322
rect 213294 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 213914 711238
rect 213294 682954 213914 711002
rect 213294 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 213914 682954
rect 213294 682634 213914 682718
rect 213294 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 213914 682634
rect 213294 664000 213914 682398
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 664000 218414 686898
rect 222294 705798 222914 711590
rect 222294 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 222914 705798
rect 222294 705478 222914 705562
rect 222294 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 222914 705478
rect 222294 691954 222914 705242
rect 222294 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 222914 691954
rect 222294 691634 222914 691718
rect 222294 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 222914 691634
rect 222294 664000 222914 691398
rect 226794 706758 227414 711590
rect 226794 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 227414 706758
rect 226794 706438 227414 706522
rect 226794 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 227414 706438
rect 226794 696454 227414 706202
rect 226794 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 227414 696454
rect 226794 696134 227414 696218
rect 226794 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 227414 696134
rect 226794 664000 227414 695898
rect 231294 707718 231914 711590
rect 231294 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 231914 707718
rect 231294 707398 231914 707482
rect 231294 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 231914 707398
rect 231294 700954 231914 707162
rect 231294 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 231914 700954
rect 231294 700634 231914 700718
rect 231294 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 231914 700634
rect 231294 664954 231914 700398
rect 231294 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 231914 664954
rect 231294 664634 231914 664718
rect 231294 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 231914 664634
rect 231294 664000 231914 664398
rect 235794 708678 236414 711590
rect 235794 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 236414 708678
rect 235794 708358 236414 708442
rect 235794 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 236414 708358
rect 235794 669454 236414 708122
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 664000 236414 668898
rect 240294 709638 240914 711590
rect 240294 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 240914 709638
rect 240294 709318 240914 709402
rect 240294 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 240914 709318
rect 240294 673954 240914 709082
rect 240294 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 240914 673954
rect 240294 673634 240914 673718
rect 240294 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 240914 673634
rect 240294 664000 240914 673398
rect 244794 710598 245414 711590
rect 244794 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 245414 710598
rect 244794 710278 245414 710362
rect 244794 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 245414 710278
rect 244794 678454 245414 710042
rect 244794 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 245414 678454
rect 244794 678134 245414 678218
rect 244794 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 245414 678134
rect 244794 664000 245414 677898
rect 249294 711558 249914 711590
rect 249294 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 249914 711558
rect 249294 711238 249914 711322
rect 249294 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 249914 711238
rect 249294 682954 249914 711002
rect 249294 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 249914 682954
rect 249294 682634 249914 682718
rect 249294 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 249914 682634
rect 249294 664000 249914 682398
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 664000 254414 686898
rect 258294 705798 258914 711590
rect 258294 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 258914 705798
rect 258294 705478 258914 705562
rect 258294 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 258914 705478
rect 258294 691954 258914 705242
rect 258294 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 258914 691954
rect 258294 691634 258914 691718
rect 258294 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 258914 691634
rect 51027 662692 51093 662693
rect 51027 662628 51028 662692
rect 51092 662628 51093 662692
rect 51027 662627 51093 662628
rect 49003 661196 49069 661197
rect 49003 661132 49004 661196
rect 49068 661132 49069 661196
rect 49003 661131 49069 661132
rect 46794 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 47414 660454
rect 46794 660134 47414 660218
rect 46794 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 47414 660134
rect 46794 624454 47414 659898
rect 46794 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 47414 624454
rect 46794 624134 47414 624218
rect 46794 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 47414 624134
rect 46794 588454 47414 623898
rect 49006 602581 49066 661131
rect 49371 660516 49437 660517
rect 49371 660452 49372 660516
rect 49436 660452 49437 660516
rect 49371 660451 49437 660452
rect 49187 660244 49253 660245
rect 49187 660180 49188 660244
rect 49252 660180 49253 660244
rect 49187 660179 49253 660180
rect 49190 614277 49250 660179
rect 49374 637669 49434 660451
rect 49923 659836 49989 659837
rect 49923 659772 49924 659836
rect 49988 659772 49989 659836
rect 49923 659771 49989 659772
rect 49739 659700 49805 659701
rect 49739 659636 49740 659700
rect 49804 659636 49805 659700
rect 49739 659635 49805 659636
rect 49371 637668 49437 637669
rect 49371 637604 49372 637668
rect 49436 637604 49437 637668
rect 49371 637603 49437 637604
rect 49371 637532 49437 637533
rect 49371 637468 49372 637532
rect 49436 637468 49437 637532
rect 49371 637467 49437 637468
rect 49187 614276 49253 614277
rect 49187 614212 49188 614276
rect 49252 614212 49253 614276
rect 49187 614211 49253 614212
rect 49003 602580 49069 602581
rect 49003 602516 49004 602580
rect 49068 602516 49069 602580
rect 49003 602515 49069 602516
rect 49187 601084 49253 601085
rect 49187 601020 49188 601084
rect 49252 601020 49253 601084
rect 49187 601019 49253 601020
rect 46794 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 47414 588454
rect 46794 588134 47414 588218
rect 46794 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 47414 588134
rect 46794 552454 47414 587898
rect 46794 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 47414 552454
rect 46794 552134 47414 552218
rect 46794 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 47414 552134
rect 46794 516454 47414 551898
rect 49190 532405 49250 601019
rect 49187 532404 49253 532405
rect 49187 532340 49188 532404
rect 49252 532340 49253 532404
rect 49187 532339 49253 532340
rect 46794 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 47414 516454
rect 46794 516134 47414 516218
rect 46794 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 47414 516134
rect 46794 480454 47414 515898
rect 46794 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 47414 480454
rect 46794 480134 47414 480218
rect 46794 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 47414 480134
rect 46794 444454 47414 479898
rect 49374 479773 49434 637467
rect 49555 612780 49621 612781
rect 49555 612716 49556 612780
rect 49620 612716 49621 612780
rect 49555 612715 49621 612716
rect 49558 608429 49618 612715
rect 49555 608428 49621 608429
rect 49555 608364 49556 608428
rect 49620 608364 49621 608428
rect 49555 608363 49621 608364
rect 49555 607204 49621 607205
rect 49555 607140 49556 607204
rect 49620 607140 49621 607204
rect 49555 607139 49621 607140
rect 49558 503165 49618 607139
rect 49555 503164 49621 503165
rect 49555 503100 49556 503164
rect 49620 503100 49621 503164
rect 49555 503099 49621 503100
rect 49742 500989 49802 659635
rect 49926 605981 49986 659771
rect 50107 659700 50173 659701
rect 50107 659636 50108 659700
rect 50172 659636 50173 659700
rect 50107 659635 50173 659636
rect 50110 618357 50170 659635
rect 50107 618356 50173 618357
rect 50107 618292 50108 618356
rect 50172 618292 50173 618356
rect 50107 618291 50173 618292
rect 49923 605980 49989 605981
rect 49923 605916 49924 605980
rect 49988 605916 49989 605980
rect 49923 605915 49989 605916
rect 49739 500988 49805 500989
rect 49739 500924 49740 500988
rect 49804 500924 49805 500988
rect 49739 500923 49805 500924
rect 51030 485621 51090 662627
rect 51579 662556 51645 662557
rect 51579 662492 51580 662556
rect 51644 662492 51645 662556
rect 51579 662491 51645 662492
rect 51582 601085 51642 662491
rect 71568 655954 71888 655986
rect 71568 655718 71610 655954
rect 71846 655718 71888 655954
rect 71568 655634 71888 655718
rect 71568 655398 71610 655634
rect 71846 655398 71888 655634
rect 71568 655366 71888 655398
rect 102288 655954 102608 655986
rect 102288 655718 102330 655954
rect 102566 655718 102608 655954
rect 102288 655634 102608 655718
rect 102288 655398 102330 655634
rect 102566 655398 102608 655634
rect 102288 655366 102608 655398
rect 133008 655954 133328 655986
rect 133008 655718 133050 655954
rect 133286 655718 133328 655954
rect 133008 655634 133328 655718
rect 133008 655398 133050 655634
rect 133286 655398 133328 655634
rect 133008 655366 133328 655398
rect 163728 655954 164048 655986
rect 163728 655718 163770 655954
rect 164006 655718 164048 655954
rect 163728 655634 164048 655718
rect 163728 655398 163770 655634
rect 164006 655398 164048 655634
rect 163728 655366 164048 655398
rect 194448 655954 194768 655986
rect 194448 655718 194490 655954
rect 194726 655718 194768 655954
rect 194448 655634 194768 655718
rect 194448 655398 194490 655634
rect 194726 655398 194768 655634
rect 194448 655366 194768 655398
rect 225168 655954 225488 655986
rect 225168 655718 225210 655954
rect 225446 655718 225488 655954
rect 225168 655634 225488 655718
rect 225168 655398 225210 655634
rect 225446 655398 225488 655634
rect 225168 655366 225488 655398
rect 258294 655954 258914 691398
rect 258294 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 258914 655954
rect 258294 655634 258914 655718
rect 258294 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 258914 655634
rect 56208 651454 56528 651486
rect 56208 651218 56250 651454
rect 56486 651218 56528 651454
rect 56208 651134 56528 651218
rect 56208 650898 56250 651134
rect 56486 650898 56528 651134
rect 56208 650866 56528 650898
rect 86928 651454 87248 651486
rect 86928 651218 86970 651454
rect 87206 651218 87248 651454
rect 86928 651134 87248 651218
rect 86928 650898 86970 651134
rect 87206 650898 87248 651134
rect 86928 650866 87248 650898
rect 117648 651454 117968 651486
rect 117648 651218 117690 651454
rect 117926 651218 117968 651454
rect 117648 651134 117968 651218
rect 117648 650898 117690 651134
rect 117926 650898 117968 651134
rect 117648 650866 117968 650898
rect 148368 651454 148688 651486
rect 148368 651218 148410 651454
rect 148646 651218 148688 651454
rect 148368 651134 148688 651218
rect 148368 650898 148410 651134
rect 148646 650898 148688 651134
rect 148368 650866 148688 650898
rect 179088 651454 179408 651486
rect 179088 651218 179130 651454
rect 179366 651218 179408 651454
rect 179088 651134 179408 651218
rect 179088 650898 179130 651134
rect 179366 650898 179408 651134
rect 179088 650866 179408 650898
rect 209808 651454 210128 651486
rect 209808 651218 209850 651454
rect 210086 651218 210128 651454
rect 209808 651134 210128 651218
rect 209808 650898 209850 651134
rect 210086 650898 210128 651134
rect 209808 650866 210128 650898
rect 240528 651454 240848 651486
rect 240528 651218 240570 651454
rect 240806 651218 240848 651454
rect 240528 651134 240848 651218
rect 240528 650898 240570 651134
rect 240806 650898 240848 651134
rect 240528 650866 240848 650898
rect 71568 619954 71888 619986
rect 71568 619718 71610 619954
rect 71846 619718 71888 619954
rect 71568 619634 71888 619718
rect 71568 619398 71610 619634
rect 71846 619398 71888 619634
rect 71568 619366 71888 619398
rect 102288 619954 102608 619986
rect 102288 619718 102330 619954
rect 102566 619718 102608 619954
rect 102288 619634 102608 619718
rect 102288 619398 102330 619634
rect 102566 619398 102608 619634
rect 102288 619366 102608 619398
rect 133008 619954 133328 619986
rect 133008 619718 133050 619954
rect 133286 619718 133328 619954
rect 133008 619634 133328 619718
rect 133008 619398 133050 619634
rect 133286 619398 133328 619634
rect 133008 619366 133328 619398
rect 163728 619954 164048 619986
rect 163728 619718 163770 619954
rect 164006 619718 164048 619954
rect 163728 619634 164048 619718
rect 163728 619398 163770 619634
rect 164006 619398 164048 619634
rect 163728 619366 164048 619398
rect 194448 619954 194768 619986
rect 194448 619718 194490 619954
rect 194726 619718 194768 619954
rect 194448 619634 194768 619718
rect 194448 619398 194490 619634
rect 194726 619398 194768 619634
rect 194448 619366 194768 619398
rect 225168 619954 225488 619986
rect 225168 619718 225210 619954
rect 225446 619718 225488 619954
rect 225168 619634 225488 619718
rect 225168 619398 225210 619634
rect 225446 619398 225488 619634
rect 225168 619366 225488 619398
rect 258294 619954 258914 655398
rect 258294 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 258914 619954
rect 258294 619634 258914 619718
rect 258294 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 258914 619634
rect 56208 615454 56528 615486
rect 56208 615218 56250 615454
rect 56486 615218 56528 615454
rect 56208 615134 56528 615218
rect 56208 614898 56250 615134
rect 56486 614898 56528 615134
rect 56208 614866 56528 614898
rect 86928 615454 87248 615486
rect 86928 615218 86970 615454
rect 87206 615218 87248 615454
rect 86928 615134 87248 615218
rect 86928 614898 86970 615134
rect 87206 614898 87248 615134
rect 86928 614866 87248 614898
rect 117648 615454 117968 615486
rect 117648 615218 117690 615454
rect 117926 615218 117968 615454
rect 117648 615134 117968 615218
rect 117648 614898 117690 615134
rect 117926 614898 117968 615134
rect 117648 614866 117968 614898
rect 148368 615454 148688 615486
rect 148368 615218 148410 615454
rect 148646 615218 148688 615454
rect 148368 615134 148688 615218
rect 148368 614898 148410 615134
rect 148646 614898 148688 615134
rect 148368 614866 148688 614898
rect 179088 615454 179408 615486
rect 179088 615218 179130 615454
rect 179366 615218 179408 615454
rect 179088 615134 179408 615218
rect 179088 614898 179130 615134
rect 179366 614898 179408 615134
rect 179088 614866 179408 614898
rect 209808 615454 210128 615486
rect 209808 615218 209850 615454
rect 210086 615218 210128 615454
rect 209808 615134 210128 615218
rect 209808 614898 209850 615134
rect 210086 614898 210128 615134
rect 209808 614866 210128 614898
rect 240528 615454 240848 615486
rect 240528 615218 240570 615454
rect 240806 615218 240848 615454
rect 240528 615134 240848 615218
rect 240528 614898 240570 615134
rect 240806 614898 240848 615134
rect 240528 614866 240848 614898
rect 51579 601084 51645 601085
rect 51579 601020 51580 601084
rect 51644 601020 51645 601084
rect 51579 601019 51645 601020
rect 71568 583954 71888 583986
rect 71568 583718 71610 583954
rect 71846 583718 71888 583954
rect 71568 583634 71888 583718
rect 71568 583398 71610 583634
rect 71846 583398 71888 583634
rect 71568 583366 71888 583398
rect 102288 583954 102608 583986
rect 102288 583718 102330 583954
rect 102566 583718 102608 583954
rect 102288 583634 102608 583718
rect 102288 583398 102330 583634
rect 102566 583398 102608 583634
rect 102288 583366 102608 583398
rect 133008 583954 133328 583986
rect 133008 583718 133050 583954
rect 133286 583718 133328 583954
rect 133008 583634 133328 583718
rect 133008 583398 133050 583634
rect 133286 583398 133328 583634
rect 133008 583366 133328 583398
rect 163728 583954 164048 583986
rect 163728 583718 163770 583954
rect 164006 583718 164048 583954
rect 163728 583634 164048 583718
rect 163728 583398 163770 583634
rect 164006 583398 164048 583634
rect 163728 583366 164048 583398
rect 194448 583954 194768 583986
rect 194448 583718 194490 583954
rect 194726 583718 194768 583954
rect 194448 583634 194768 583718
rect 194448 583398 194490 583634
rect 194726 583398 194768 583634
rect 194448 583366 194768 583398
rect 225168 583954 225488 583986
rect 225168 583718 225210 583954
rect 225446 583718 225488 583954
rect 225168 583634 225488 583718
rect 225168 583398 225210 583634
rect 225446 583398 225488 583634
rect 225168 583366 225488 583398
rect 258294 583954 258914 619398
rect 258294 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 258914 583954
rect 258294 583634 258914 583718
rect 258294 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 258914 583634
rect 56208 579454 56528 579486
rect 56208 579218 56250 579454
rect 56486 579218 56528 579454
rect 56208 579134 56528 579218
rect 56208 578898 56250 579134
rect 56486 578898 56528 579134
rect 56208 578866 56528 578898
rect 86928 579454 87248 579486
rect 86928 579218 86970 579454
rect 87206 579218 87248 579454
rect 86928 579134 87248 579218
rect 86928 578898 86970 579134
rect 87206 578898 87248 579134
rect 86928 578866 87248 578898
rect 117648 579454 117968 579486
rect 117648 579218 117690 579454
rect 117926 579218 117968 579454
rect 117648 579134 117968 579218
rect 117648 578898 117690 579134
rect 117926 578898 117968 579134
rect 117648 578866 117968 578898
rect 148368 579454 148688 579486
rect 148368 579218 148410 579454
rect 148646 579218 148688 579454
rect 148368 579134 148688 579218
rect 148368 578898 148410 579134
rect 148646 578898 148688 579134
rect 148368 578866 148688 578898
rect 179088 579454 179408 579486
rect 179088 579218 179130 579454
rect 179366 579218 179408 579454
rect 179088 579134 179408 579218
rect 179088 578898 179130 579134
rect 179366 578898 179408 579134
rect 179088 578866 179408 578898
rect 209808 579454 210128 579486
rect 209808 579218 209850 579454
rect 210086 579218 210128 579454
rect 209808 579134 210128 579218
rect 209808 578898 209850 579134
rect 210086 578898 210128 579134
rect 209808 578866 210128 578898
rect 240528 579454 240848 579486
rect 240528 579218 240570 579454
rect 240806 579218 240848 579454
rect 240528 579134 240848 579218
rect 240528 578898 240570 579134
rect 240806 578898 240848 579134
rect 240528 578866 240848 578898
rect 71568 547954 71888 547986
rect 71568 547718 71610 547954
rect 71846 547718 71888 547954
rect 71568 547634 71888 547718
rect 71568 547398 71610 547634
rect 71846 547398 71888 547634
rect 71568 547366 71888 547398
rect 102288 547954 102608 547986
rect 102288 547718 102330 547954
rect 102566 547718 102608 547954
rect 102288 547634 102608 547718
rect 102288 547398 102330 547634
rect 102566 547398 102608 547634
rect 102288 547366 102608 547398
rect 133008 547954 133328 547986
rect 133008 547718 133050 547954
rect 133286 547718 133328 547954
rect 133008 547634 133328 547718
rect 133008 547398 133050 547634
rect 133286 547398 133328 547634
rect 133008 547366 133328 547398
rect 163728 547954 164048 547986
rect 163728 547718 163770 547954
rect 164006 547718 164048 547954
rect 163728 547634 164048 547718
rect 163728 547398 163770 547634
rect 164006 547398 164048 547634
rect 163728 547366 164048 547398
rect 194448 547954 194768 547986
rect 194448 547718 194490 547954
rect 194726 547718 194768 547954
rect 194448 547634 194768 547718
rect 194448 547398 194490 547634
rect 194726 547398 194768 547634
rect 194448 547366 194768 547398
rect 225168 547954 225488 547986
rect 225168 547718 225210 547954
rect 225446 547718 225488 547954
rect 225168 547634 225488 547718
rect 225168 547398 225210 547634
rect 225446 547398 225488 547634
rect 225168 547366 225488 547398
rect 258294 547954 258914 583398
rect 258294 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 258914 547954
rect 258294 547634 258914 547718
rect 258294 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 258914 547634
rect 56208 543454 56528 543486
rect 56208 543218 56250 543454
rect 56486 543218 56528 543454
rect 56208 543134 56528 543218
rect 56208 542898 56250 543134
rect 56486 542898 56528 543134
rect 56208 542866 56528 542898
rect 86928 543454 87248 543486
rect 86928 543218 86970 543454
rect 87206 543218 87248 543454
rect 86928 543134 87248 543218
rect 86928 542898 86970 543134
rect 87206 542898 87248 543134
rect 86928 542866 87248 542898
rect 117648 543454 117968 543486
rect 117648 543218 117690 543454
rect 117926 543218 117968 543454
rect 117648 543134 117968 543218
rect 117648 542898 117690 543134
rect 117926 542898 117968 543134
rect 117648 542866 117968 542898
rect 148368 543454 148688 543486
rect 148368 543218 148410 543454
rect 148646 543218 148688 543454
rect 148368 543134 148688 543218
rect 148368 542898 148410 543134
rect 148646 542898 148688 543134
rect 148368 542866 148688 542898
rect 179088 543454 179408 543486
rect 179088 543218 179130 543454
rect 179366 543218 179408 543454
rect 179088 543134 179408 543218
rect 179088 542898 179130 543134
rect 179366 542898 179408 543134
rect 179088 542866 179408 542898
rect 209808 543454 210128 543486
rect 209808 543218 209850 543454
rect 210086 543218 210128 543454
rect 209808 543134 210128 543218
rect 209808 542898 209850 543134
rect 210086 542898 210128 543134
rect 209808 542866 210128 542898
rect 240528 543454 240848 543486
rect 240528 543218 240570 543454
rect 240806 543218 240848 543454
rect 240528 543134 240848 543218
rect 240528 542898 240570 543134
rect 240806 542898 240848 543134
rect 240528 542866 240848 542898
rect 71568 511954 71888 511986
rect 71568 511718 71610 511954
rect 71846 511718 71888 511954
rect 71568 511634 71888 511718
rect 71568 511398 71610 511634
rect 71846 511398 71888 511634
rect 71568 511366 71888 511398
rect 102288 511954 102608 511986
rect 102288 511718 102330 511954
rect 102566 511718 102608 511954
rect 102288 511634 102608 511718
rect 102288 511398 102330 511634
rect 102566 511398 102608 511634
rect 102288 511366 102608 511398
rect 133008 511954 133328 511986
rect 133008 511718 133050 511954
rect 133286 511718 133328 511954
rect 133008 511634 133328 511718
rect 133008 511398 133050 511634
rect 133286 511398 133328 511634
rect 133008 511366 133328 511398
rect 163728 511954 164048 511986
rect 163728 511718 163770 511954
rect 164006 511718 164048 511954
rect 163728 511634 164048 511718
rect 163728 511398 163770 511634
rect 164006 511398 164048 511634
rect 163728 511366 164048 511398
rect 194448 511954 194768 511986
rect 194448 511718 194490 511954
rect 194726 511718 194768 511954
rect 194448 511634 194768 511718
rect 194448 511398 194490 511634
rect 194726 511398 194768 511634
rect 194448 511366 194768 511398
rect 225168 511954 225488 511986
rect 225168 511718 225210 511954
rect 225446 511718 225488 511954
rect 225168 511634 225488 511718
rect 225168 511398 225210 511634
rect 225446 511398 225488 511634
rect 225168 511366 225488 511398
rect 258294 511954 258914 547398
rect 258294 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 258914 511954
rect 258294 511634 258914 511718
rect 258294 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 258914 511634
rect 56208 507454 56528 507486
rect 56208 507218 56250 507454
rect 56486 507218 56528 507454
rect 56208 507134 56528 507218
rect 56208 506898 56250 507134
rect 56486 506898 56528 507134
rect 56208 506866 56528 506898
rect 86928 507454 87248 507486
rect 86928 507218 86970 507454
rect 87206 507218 87248 507454
rect 86928 507134 87248 507218
rect 86928 506898 86970 507134
rect 87206 506898 87248 507134
rect 86928 506866 87248 506898
rect 117648 507454 117968 507486
rect 117648 507218 117690 507454
rect 117926 507218 117968 507454
rect 117648 507134 117968 507218
rect 117648 506898 117690 507134
rect 117926 506898 117968 507134
rect 117648 506866 117968 506898
rect 148368 507454 148688 507486
rect 148368 507218 148410 507454
rect 148646 507218 148688 507454
rect 148368 507134 148688 507218
rect 148368 506898 148410 507134
rect 148646 506898 148688 507134
rect 148368 506866 148688 506898
rect 179088 507454 179408 507486
rect 179088 507218 179130 507454
rect 179366 507218 179408 507454
rect 179088 507134 179408 507218
rect 179088 506898 179130 507134
rect 179366 506898 179408 507134
rect 179088 506866 179408 506898
rect 209808 507454 210128 507486
rect 209808 507218 209850 507454
rect 210086 507218 210128 507454
rect 209808 507134 210128 507218
rect 209808 506898 209850 507134
rect 210086 506898 210128 507134
rect 209808 506866 210128 506898
rect 240528 507454 240848 507486
rect 240528 507218 240570 507454
rect 240806 507218 240848 507454
rect 240528 507134 240848 507218
rect 240528 506898 240570 507134
rect 240806 506898 240848 507134
rect 240528 506866 240848 506898
rect 51027 485620 51093 485621
rect 51027 485556 51028 485620
rect 51092 485556 51093 485620
rect 51027 485555 51093 485556
rect 49555 484396 49621 484397
rect 49555 484332 49556 484396
rect 49620 484332 49621 484396
rect 49555 484331 49621 484332
rect 49371 479772 49437 479773
rect 49371 479708 49372 479772
rect 49436 479708 49437 479772
rect 49371 479707 49437 479708
rect 46794 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 47414 444454
rect 46794 444134 47414 444218
rect 46794 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 47414 444134
rect 46794 408454 47414 443898
rect 46794 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 47414 408454
rect 46794 408134 47414 408218
rect 46794 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 47414 408134
rect 46794 372454 47414 407898
rect 46794 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 47414 372454
rect 46794 372134 47414 372218
rect 46794 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 47414 372134
rect 46794 336454 47414 371898
rect 46794 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 47414 336454
rect 46794 336134 47414 336218
rect 46794 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 47414 336134
rect 46794 300454 47414 335898
rect 46794 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 47414 300454
rect 46794 300134 47414 300218
rect 46794 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 47414 300134
rect 46794 264454 47414 299898
rect 49374 278765 49434 479707
rect 49371 278764 49437 278765
rect 49371 278700 49372 278764
rect 49436 278700 49437 278764
rect 49371 278699 49437 278700
rect 46794 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 47414 264454
rect 46794 264134 47414 264218
rect 46794 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 47414 264134
rect 46794 228454 47414 263898
rect 46794 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 47414 228454
rect 46794 228134 47414 228218
rect 46794 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 47414 228134
rect 46794 192454 47414 227898
rect 49558 223549 49618 484331
rect 71568 475954 71888 475986
rect 71568 475718 71610 475954
rect 71846 475718 71888 475954
rect 71568 475634 71888 475718
rect 71568 475398 71610 475634
rect 71846 475398 71888 475634
rect 71568 475366 71888 475398
rect 102288 475954 102608 475986
rect 102288 475718 102330 475954
rect 102566 475718 102608 475954
rect 102288 475634 102608 475718
rect 102288 475398 102330 475634
rect 102566 475398 102608 475634
rect 102288 475366 102608 475398
rect 133008 475954 133328 475986
rect 133008 475718 133050 475954
rect 133286 475718 133328 475954
rect 133008 475634 133328 475718
rect 133008 475398 133050 475634
rect 133286 475398 133328 475634
rect 133008 475366 133328 475398
rect 163728 475954 164048 475986
rect 163728 475718 163770 475954
rect 164006 475718 164048 475954
rect 163728 475634 164048 475718
rect 163728 475398 163770 475634
rect 164006 475398 164048 475634
rect 163728 475366 164048 475398
rect 194448 475954 194768 475986
rect 194448 475718 194490 475954
rect 194726 475718 194768 475954
rect 194448 475634 194768 475718
rect 194448 475398 194490 475634
rect 194726 475398 194768 475634
rect 194448 475366 194768 475398
rect 225168 475954 225488 475986
rect 225168 475718 225210 475954
rect 225446 475718 225488 475954
rect 225168 475634 225488 475718
rect 225168 475398 225210 475634
rect 225446 475398 225488 475634
rect 225168 475366 225488 475398
rect 258294 475954 258914 511398
rect 258294 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 258914 475954
rect 258294 475634 258914 475718
rect 258294 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 258914 475634
rect 56208 471454 56528 471486
rect 56208 471218 56250 471454
rect 56486 471218 56528 471454
rect 56208 471134 56528 471218
rect 56208 470898 56250 471134
rect 56486 470898 56528 471134
rect 56208 470866 56528 470898
rect 86928 471454 87248 471486
rect 86928 471218 86970 471454
rect 87206 471218 87248 471454
rect 86928 471134 87248 471218
rect 86928 470898 86970 471134
rect 87206 470898 87248 471134
rect 86928 470866 87248 470898
rect 117648 471454 117968 471486
rect 117648 471218 117690 471454
rect 117926 471218 117968 471454
rect 117648 471134 117968 471218
rect 117648 470898 117690 471134
rect 117926 470898 117968 471134
rect 117648 470866 117968 470898
rect 148368 471454 148688 471486
rect 148368 471218 148410 471454
rect 148646 471218 148688 471454
rect 148368 471134 148688 471218
rect 148368 470898 148410 471134
rect 148646 470898 148688 471134
rect 148368 470866 148688 470898
rect 179088 471454 179408 471486
rect 179088 471218 179130 471454
rect 179366 471218 179408 471454
rect 179088 471134 179408 471218
rect 179088 470898 179130 471134
rect 179366 470898 179408 471134
rect 179088 470866 179408 470898
rect 209808 471454 210128 471486
rect 209808 471218 209850 471454
rect 210086 471218 210128 471454
rect 209808 471134 210128 471218
rect 209808 470898 209850 471134
rect 210086 470898 210128 471134
rect 209808 470866 210128 470898
rect 240528 471454 240848 471486
rect 240528 471218 240570 471454
rect 240806 471218 240848 471454
rect 240528 471134 240848 471218
rect 240528 470898 240570 471134
rect 240806 470898 240848 471134
rect 240528 470866 240848 470898
rect 71568 439954 71888 439986
rect 71568 439718 71610 439954
rect 71846 439718 71888 439954
rect 71568 439634 71888 439718
rect 71568 439398 71610 439634
rect 71846 439398 71888 439634
rect 71568 439366 71888 439398
rect 102288 439954 102608 439986
rect 102288 439718 102330 439954
rect 102566 439718 102608 439954
rect 102288 439634 102608 439718
rect 102288 439398 102330 439634
rect 102566 439398 102608 439634
rect 102288 439366 102608 439398
rect 133008 439954 133328 439986
rect 133008 439718 133050 439954
rect 133286 439718 133328 439954
rect 133008 439634 133328 439718
rect 133008 439398 133050 439634
rect 133286 439398 133328 439634
rect 133008 439366 133328 439398
rect 163728 439954 164048 439986
rect 163728 439718 163770 439954
rect 164006 439718 164048 439954
rect 163728 439634 164048 439718
rect 163728 439398 163770 439634
rect 164006 439398 164048 439634
rect 163728 439366 164048 439398
rect 194448 439954 194768 439986
rect 194448 439718 194490 439954
rect 194726 439718 194768 439954
rect 194448 439634 194768 439718
rect 194448 439398 194490 439634
rect 194726 439398 194768 439634
rect 194448 439366 194768 439398
rect 225168 439954 225488 439986
rect 225168 439718 225210 439954
rect 225446 439718 225488 439954
rect 225168 439634 225488 439718
rect 225168 439398 225210 439634
rect 225446 439398 225488 439634
rect 225168 439366 225488 439398
rect 258294 439954 258914 475398
rect 258294 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 258914 439954
rect 258294 439634 258914 439718
rect 258294 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 258914 439634
rect 56208 435454 56528 435486
rect 56208 435218 56250 435454
rect 56486 435218 56528 435454
rect 56208 435134 56528 435218
rect 56208 434898 56250 435134
rect 56486 434898 56528 435134
rect 56208 434866 56528 434898
rect 86928 435454 87248 435486
rect 86928 435218 86970 435454
rect 87206 435218 87248 435454
rect 86928 435134 87248 435218
rect 86928 434898 86970 435134
rect 87206 434898 87248 435134
rect 86928 434866 87248 434898
rect 117648 435454 117968 435486
rect 117648 435218 117690 435454
rect 117926 435218 117968 435454
rect 117648 435134 117968 435218
rect 117648 434898 117690 435134
rect 117926 434898 117968 435134
rect 117648 434866 117968 434898
rect 148368 435454 148688 435486
rect 148368 435218 148410 435454
rect 148646 435218 148688 435454
rect 148368 435134 148688 435218
rect 148368 434898 148410 435134
rect 148646 434898 148688 435134
rect 148368 434866 148688 434898
rect 179088 435454 179408 435486
rect 179088 435218 179130 435454
rect 179366 435218 179408 435454
rect 179088 435134 179408 435218
rect 179088 434898 179130 435134
rect 179366 434898 179408 435134
rect 179088 434866 179408 434898
rect 209808 435454 210128 435486
rect 209808 435218 209850 435454
rect 210086 435218 210128 435454
rect 209808 435134 210128 435218
rect 209808 434898 209850 435134
rect 210086 434898 210128 435134
rect 209808 434866 210128 434898
rect 240528 435454 240848 435486
rect 240528 435218 240570 435454
rect 240806 435218 240848 435454
rect 240528 435134 240848 435218
rect 240528 434898 240570 435134
rect 240806 434898 240848 435134
rect 240528 434866 240848 434898
rect 71568 403954 71888 403986
rect 71568 403718 71610 403954
rect 71846 403718 71888 403954
rect 71568 403634 71888 403718
rect 71568 403398 71610 403634
rect 71846 403398 71888 403634
rect 71568 403366 71888 403398
rect 102288 403954 102608 403986
rect 102288 403718 102330 403954
rect 102566 403718 102608 403954
rect 102288 403634 102608 403718
rect 102288 403398 102330 403634
rect 102566 403398 102608 403634
rect 102288 403366 102608 403398
rect 133008 403954 133328 403986
rect 133008 403718 133050 403954
rect 133286 403718 133328 403954
rect 133008 403634 133328 403718
rect 133008 403398 133050 403634
rect 133286 403398 133328 403634
rect 133008 403366 133328 403398
rect 163728 403954 164048 403986
rect 163728 403718 163770 403954
rect 164006 403718 164048 403954
rect 163728 403634 164048 403718
rect 163728 403398 163770 403634
rect 164006 403398 164048 403634
rect 163728 403366 164048 403398
rect 194448 403954 194768 403986
rect 194448 403718 194490 403954
rect 194726 403718 194768 403954
rect 194448 403634 194768 403718
rect 194448 403398 194490 403634
rect 194726 403398 194768 403634
rect 194448 403366 194768 403398
rect 225168 403954 225488 403986
rect 225168 403718 225210 403954
rect 225446 403718 225488 403954
rect 225168 403634 225488 403718
rect 225168 403398 225210 403634
rect 225446 403398 225488 403634
rect 225168 403366 225488 403398
rect 258294 403954 258914 439398
rect 258294 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 258914 403954
rect 258294 403634 258914 403718
rect 258294 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 258914 403634
rect 56208 399454 56528 399486
rect 56208 399218 56250 399454
rect 56486 399218 56528 399454
rect 56208 399134 56528 399218
rect 56208 398898 56250 399134
rect 56486 398898 56528 399134
rect 56208 398866 56528 398898
rect 86928 399454 87248 399486
rect 86928 399218 86970 399454
rect 87206 399218 87248 399454
rect 86928 399134 87248 399218
rect 86928 398898 86970 399134
rect 87206 398898 87248 399134
rect 86928 398866 87248 398898
rect 117648 399454 117968 399486
rect 117648 399218 117690 399454
rect 117926 399218 117968 399454
rect 117648 399134 117968 399218
rect 117648 398898 117690 399134
rect 117926 398898 117968 399134
rect 117648 398866 117968 398898
rect 148368 399454 148688 399486
rect 148368 399218 148410 399454
rect 148646 399218 148688 399454
rect 148368 399134 148688 399218
rect 148368 398898 148410 399134
rect 148646 398898 148688 399134
rect 148368 398866 148688 398898
rect 179088 399454 179408 399486
rect 179088 399218 179130 399454
rect 179366 399218 179408 399454
rect 179088 399134 179408 399218
rect 179088 398898 179130 399134
rect 179366 398898 179408 399134
rect 179088 398866 179408 398898
rect 209808 399454 210128 399486
rect 209808 399218 209850 399454
rect 210086 399218 210128 399454
rect 209808 399134 210128 399218
rect 209808 398898 209850 399134
rect 210086 398898 210128 399134
rect 209808 398866 210128 398898
rect 240528 399454 240848 399486
rect 240528 399218 240570 399454
rect 240806 399218 240848 399454
rect 240528 399134 240848 399218
rect 240528 398898 240570 399134
rect 240806 398898 240848 399134
rect 240528 398866 240848 398898
rect 71568 367954 71888 367986
rect 71568 367718 71610 367954
rect 71846 367718 71888 367954
rect 71568 367634 71888 367718
rect 71568 367398 71610 367634
rect 71846 367398 71888 367634
rect 71568 367366 71888 367398
rect 102288 367954 102608 367986
rect 102288 367718 102330 367954
rect 102566 367718 102608 367954
rect 102288 367634 102608 367718
rect 102288 367398 102330 367634
rect 102566 367398 102608 367634
rect 102288 367366 102608 367398
rect 133008 367954 133328 367986
rect 133008 367718 133050 367954
rect 133286 367718 133328 367954
rect 133008 367634 133328 367718
rect 133008 367398 133050 367634
rect 133286 367398 133328 367634
rect 133008 367366 133328 367398
rect 163728 367954 164048 367986
rect 163728 367718 163770 367954
rect 164006 367718 164048 367954
rect 163728 367634 164048 367718
rect 163728 367398 163770 367634
rect 164006 367398 164048 367634
rect 163728 367366 164048 367398
rect 194448 367954 194768 367986
rect 194448 367718 194490 367954
rect 194726 367718 194768 367954
rect 194448 367634 194768 367718
rect 194448 367398 194490 367634
rect 194726 367398 194768 367634
rect 194448 367366 194768 367398
rect 225168 367954 225488 367986
rect 225168 367718 225210 367954
rect 225446 367718 225488 367954
rect 225168 367634 225488 367718
rect 225168 367398 225210 367634
rect 225446 367398 225488 367634
rect 225168 367366 225488 367398
rect 258294 367954 258914 403398
rect 258294 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 258914 367954
rect 258294 367634 258914 367718
rect 258294 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 258914 367634
rect 56208 363454 56528 363486
rect 56208 363218 56250 363454
rect 56486 363218 56528 363454
rect 56208 363134 56528 363218
rect 56208 362898 56250 363134
rect 56486 362898 56528 363134
rect 56208 362866 56528 362898
rect 86928 363454 87248 363486
rect 86928 363218 86970 363454
rect 87206 363218 87248 363454
rect 86928 363134 87248 363218
rect 86928 362898 86970 363134
rect 87206 362898 87248 363134
rect 86928 362866 87248 362898
rect 117648 363454 117968 363486
rect 117648 363218 117690 363454
rect 117926 363218 117968 363454
rect 117648 363134 117968 363218
rect 117648 362898 117690 363134
rect 117926 362898 117968 363134
rect 117648 362866 117968 362898
rect 148368 363454 148688 363486
rect 148368 363218 148410 363454
rect 148646 363218 148688 363454
rect 148368 363134 148688 363218
rect 148368 362898 148410 363134
rect 148646 362898 148688 363134
rect 148368 362866 148688 362898
rect 179088 363454 179408 363486
rect 179088 363218 179130 363454
rect 179366 363218 179408 363454
rect 179088 363134 179408 363218
rect 179088 362898 179130 363134
rect 179366 362898 179408 363134
rect 179088 362866 179408 362898
rect 209808 363454 210128 363486
rect 209808 363218 209850 363454
rect 210086 363218 210128 363454
rect 209808 363134 210128 363218
rect 209808 362898 209850 363134
rect 210086 362898 210128 363134
rect 209808 362866 210128 362898
rect 240528 363454 240848 363486
rect 240528 363218 240570 363454
rect 240806 363218 240848 363454
rect 240528 363134 240848 363218
rect 240528 362898 240570 363134
rect 240806 362898 240848 363134
rect 240528 362866 240848 362898
rect 71568 331954 71888 331986
rect 71568 331718 71610 331954
rect 71846 331718 71888 331954
rect 71568 331634 71888 331718
rect 71568 331398 71610 331634
rect 71846 331398 71888 331634
rect 71568 331366 71888 331398
rect 102288 331954 102608 331986
rect 102288 331718 102330 331954
rect 102566 331718 102608 331954
rect 102288 331634 102608 331718
rect 102288 331398 102330 331634
rect 102566 331398 102608 331634
rect 102288 331366 102608 331398
rect 133008 331954 133328 331986
rect 133008 331718 133050 331954
rect 133286 331718 133328 331954
rect 133008 331634 133328 331718
rect 133008 331398 133050 331634
rect 133286 331398 133328 331634
rect 133008 331366 133328 331398
rect 163728 331954 164048 331986
rect 163728 331718 163770 331954
rect 164006 331718 164048 331954
rect 163728 331634 164048 331718
rect 163728 331398 163770 331634
rect 164006 331398 164048 331634
rect 163728 331366 164048 331398
rect 194448 331954 194768 331986
rect 194448 331718 194490 331954
rect 194726 331718 194768 331954
rect 194448 331634 194768 331718
rect 194448 331398 194490 331634
rect 194726 331398 194768 331634
rect 194448 331366 194768 331398
rect 225168 331954 225488 331986
rect 225168 331718 225210 331954
rect 225446 331718 225488 331954
rect 225168 331634 225488 331718
rect 225168 331398 225210 331634
rect 225446 331398 225488 331634
rect 225168 331366 225488 331398
rect 258294 331954 258914 367398
rect 258294 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 258914 331954
rect 258294 331634 258914 331718
rect 258294 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 258914 331634
rect 56208 327454 56528 327486
rect 56208 327218 56250 327454
rect 56486 327218 56528 327454
rect 56208 327134 56528 327218
rect 56208 326898 56250 327134
rect 56486 326898 56528 327134
rect 56208 326866 56528 326898
rect 86928 327454 87248 327486
rect 86928 327218 86970 327454
rect 87206 327218 87248 327454
rect 86928 327134 87248 327218
rect 86928 326898 86970 327134
rect 87206 326898 87248 327134
rect 86928 326866 87248 326898
rect 117648 327454 117968 327486
rect 117648 327218 117690 327454
rect 117926 327218 117968 327454
rect 117648 327134 117968 327218
rect 117648 326898 117690 327134
rect 117926 326898 117968 327134
rect 117648 326866 117968 326898
rect 148368 327454 148688 327486
rect 148368 327218 148410 327454
rect 148646 327218 148688 327454
rect 148368 327134 148688 327218
rect 148368 326898 148410 327134
rect 148646 326898 148688 327134
rect 148368 326866 148688 326898
rect 179088 327454 179408 327486
rect 179088 327218 179130 327454
rect 179366 327218 179408 327454
rect 179088 327134 179408 327218
rect 179088 326898 179130 327134
rect 179366 326898 179408 327134
rect 179088 326866 179408 326898
rect 209808 327454 210128 327486
rect 209808 327218 209850 327454
rect 210086 327218 210128 327454
rect 209808 327134 210128 327218
rect 209808 326898 209850 327134
rect 210086 326898 210128 327134
rect 209808 326866 210128 326898
rect 240528 327454 240848 327486
rect 240528 327218 240570 327454
rect 240806 327218 240848 327454
rect 240528 327134 240848 327218
rect 240528 326898 240570 327134
rect 240806 326898 240848 327134
rect 240528 326866 240848 326898
rect 71568 295954 71888 295986
rect 71568 295718 71610 295954
rect 71846 295718 71888 295954
rect 71568 295634 71888 295718
rect 71568 295398 71610 295634
rect 71846 295398 71888 295634
rect 71568 295366 71888 295398
rect 102288 295954 102608 295986
rect 102288 295718 102330 295954
rect 102566 295718 102608 295954
rect 102288 295634 102608 295718
rect 102288 295398 102330 295634
rect 102566 295398 102608 295634
rect 102288 295366 102608 295398
rect 133008 295954 133328 295986
rect 133008 295718 133050 295954
rect 133286 295718 133328 295954
rect 133008 295634 133328 295718
rect 133008 295398 133050 295634
rect 133286 295398 133328 295634
rect 133008 295366 133328 295398
rect 163728 295954 164048 295986
rect 163728 295718 163770 295954
rect 164006 295718 164048 295954
rect 163728 295634 164048 295718
rect 163728 295398 163770 295634
rect 164006 295398 164048 295634
rect 163728 295366 164048 295398
rect 194448 295954 194768 295986
rect 194448 295718 194490 295954
rect 194726 295718 194768 295954
rect 194448 295634 194768 295718
rect 194448 295398 194490 295634
rect 194726 295398 194768 295634
rect 194448 295366 194768 295398
rect 225168 295954 225488 295986
rect 225168 295718 225210 295954
rect 225446 295718 225488 295954
rect 225168 295634 225488 295718
rect 225168 295398 225210 295634
rect 225446 295398 225488 295634
rect 225168 295366 225488 295398
rect 258294 295954 258914 331398
rect 258294 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 258914 295954
rect 258294 295634 258914 295718
rect 258294 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 258914 295634
rect 56208 291454 56528 291486
rect 56208 291218 56250 291454
rect 56486 291218 56528 291454
rect 56208 291134 56528 291218
rect 56208 290898 56250 291134
rect 56486 290898 56528 291134
rect 56208 290866 56528 290898
rect 86928 291454 87248 291486
rect 86928 291218 86970 291454
rect 87206 291218 87248 291454
rect 86928 291134 87248 291218
rect 86928 290898 86970 291134
rect 87206 290898 87248 291134
rect 86928 290866 87248 290898
rect 117648 291454 117968 291486
rect 117648 291218 117690 291454
rect 117926 291218 117968 291454
rect 117648 291134 117968 291218
rect 117648 290898 117690 291134
rect 117926 290898 117968 291134
rect 117648 290866 117968 290898
rect 148368 291454 148688 291486
rect 148368 291218 148410 291454
rect 148646 291218 148688 291454
rect 148368 291134 148688 291218
rect 148368 290898 148410 291134
rect 148646 290898 148688 291134
rect 148368 290866 148688 290898
rect 179088 291454 179408 291486
rect 179088 291218 179130 291454
rect 179366 291218 179408 291454
rect 179088 291134 179408 291218
rect 179088 290898 179130 291134
rect 179366 290898 179408 291134
rect 179088 290866 179408 290898
rect 209808 291454 210128 291486
rect 209808 291218 209850 291454
rect 210086 291218 210128 291454
rect 209808 291134 210128 291218
rect 209808 290898 209850 291134
rect 210086 290898 210128 291134
rect 209808 290866 210128 290898
rect 240528 291454 240848 291486
rect 240528 291218 240570 291454
rect 240806 291218 240848 291454
rect 240528 291134 240848 291218
rect 240528 290898 240570 291134
rect 240806 290898 240848 291134
rect 240528 290866 240848 290898
rect 51294 268954 51914 278000
rect 51294 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 51914 268954
rect 51294 268634 51914 268718
rect 51294 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 51914 268634
rect 51294 232954 51914 268398
rect 51294 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 51914 232954
rect 51294 232634 51914 232718
rect 51294 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 51914 232634
rect 49555 223548 49621 223549
rect 49555 223484 49556 223548
rect 49620 223484 49621 223548
rect 49555 223483 49621 223484
rect 46794 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 47414 192454
rect 46794 192134 47414 192218
rect 46794 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 47414 192134
rect 46794 156454 47414 191898
rect 46794 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 47414 156454
rect 46794 156134 47414 156218
rect 46794 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 47414 156134
rect 46794 120454 47414 155898
rect 46794 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 47414 120454
rect 46794 120134 47414 120218
rect 46794 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 47414 120134
rect 46794 84454 47414 119898
rect 46794 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 47414 84454
rect 46794 84134 47414 84218
rect 46794 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 47414 84134
rect 46794 48454 47414 83898
rect 46794 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 47414 48454
rect 46794 48134 47414 48218
rect 46794 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 47414 48134
rect 46794 12454 47414 47898
rect 46794 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 47414 12454
rect 46794 12134 47414 12218
rect 46794 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 47414 12134
rect 46794 -2266 47414 11898
rect 46794 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 47414 -2266
rect 46794 -2586 47414 -2502
rect 46794 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 47414 -2586
rect 46794 -7654 47414 -2822
rect 51294 196954 51914 232398
rect 55794 273454 56414 278000
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 222000 56414 236898
rect 60294 277954 60914 278000
rect 60294 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 60914 277954
rect 60294 277634 60914 277718
rect 60294 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 60914 277634
rect 60294 241954 60914 277398
rect 60294 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 60914 241954
rect 60294 241634 60914 241718
rect 60294 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 60914 241634
rect 57835 227084 57901 227085
rect 57835 227020 57836 227084
rect 57900 227020 57901 227084
rect 57835 227019 57901 227020
rect 51294 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 51914 196954
rect 51294 196634 51914 196718
rect 51294 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 51914 196634
rect 51294 160954 51914 196398
rect 51294 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 51914 160954
rect 51294 160634 51914 160718
rect 51294 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 51914 160634
rect 51294 124954 51914 160398
rect 57838 131749 57898 227019
rect 60294 222000 60914 241398
rect 78294 259954 78914 278000
rect 78294 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 78914 259954
rect 78294 259634 78914 259718
rect 78294 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 78914 259634
rect 78294 223954 78914 259398
rect 78294 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 78914 223954
rect 78294 223634 78914 223718
rect 78294 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 78914 223634
rect 78294 222000 78914 223398
rect 82794 264454 83414 278000
rect 82794 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 83414 264454
rect 82794 264134 83414 264218
rect 82794 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 83414 264134
rect 82794 228454 83414 263898
rect 82794 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 83414 228454
rect 82794 228134 83414 228218
rect 82794 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 83414 228134
rect 82794 222000 83414 227898
rect 87294 268954 87914 278000
rect 87294 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 87914 268954
rect 87294 268634 87914 268718
rect 87294 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 87914 268634
rect 87294 232954 87914 268398
rect 87294 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 87914 232954
rect 87294 232634 87914 232718
rect 87294 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 87914 232634
rect 87294 222000 87914 232398
rect 91794 273454 92414 278000
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 222000 92414 236898
rect 96294 277954 96914 278000
rect 96294 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 96914 277954
rect 96294 277634 96914 277718
rect 96294 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 96914 277634
rect 96294 241954 96914 277398
rect 96294 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 96914 241954
rect 96294 241634 96914 241718
rect 96294 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 96914 241634
rect 96294 222000 96914 241398
rect 114294 259954 114914 278000
rect 114294 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 114914 259954
rect 114294 259634 114914 259718
rect 114294 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 114914 259634
rect 114294 223954 114914 259398
rect 114294 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 114914 223954
rect 114294 223634 114914 223718
rect 114294 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 114914 223634
rect 114294 222000 114914 223398
rect 118794 264454 119414 278000
rect 118794 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 119414 264454
rect 118794 264134 119414 264218
rect 118794 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 119414 264134
rect 118794 228454 119414 263898
rect 118794 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 119414 228454
rect 118794 228134 119414 228218
rect 118794 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 119414 228134
rect 118794 222000 119414 227898
rect 123294 268954 123914 278000
rect 123294 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 123914 268954
rect 123294 268634 123914 268718
rect 123294 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 123914 268634
rect 123294 232954 123914 268398
rect 123294 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 123914 232954
rect 123294 232634 123914 232718
rect 123294 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 123914 232634
rect 123294 222000 123914 232398
rect 127794 273454 128414 278000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 222000 128414 236898
rect 132294 277954 132914 278000
rect 132294 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 132914 277954
rect 132294 277634 132914 277718
rect 132294 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 132914 277634
rect 132294 241954 132914 277398
rect 132294 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 132914 241954
rect 132294 241634 132914 241718
rect 132294 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 132914 241634
rect 132294 222000 132914 241398
rect 150294 259954 150914 278000
rect 150294 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 150914 259954
rect 150294 259634 150914 259718
rect 150294 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 150914 259634
rect 150294 223954 150914 259398
rect 150294 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 150914 223954
rect 150294 223634 150914 223718
rect 150294 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 150914 223634
rect 150294 222000 150914 223398
rect 154794 264454 155414 278000
rect 154794 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 155414 264454
rect 154794 264134 155414 264218
rect 154794 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 155414 264134
rect 154794 228454 155414 263898
rect 154794 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 155414 228454
rect 154794 228134 155414 228218
rect 154794 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 155414 228134
rect 154794 222000 155414 227898
rect 159294 268954 159914 278000
rect 159294 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 159914 268954
rect 159294 268634 159914 268718
rect 159294 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 159914 268634
rect 159294 232954 159914 268398
rect 159294 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 159914 232954
rect 159294 232634 159914 232718
rect 159294 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 159914 232634
rect 159294 222000 159914 232398
rect 163794 273454 164414 278000
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 222000 164414 236898
rect 168294 277954 168914 278000
rect 168294 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 168914 277954
rect 168294 277634 168914 277718
rect 168294 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 168914 277634
rect 168294 241954 168914 277398
rect 168294 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 168914 241954
rect 168294 241634 168914 241718
rect 168294 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 168914 241634
rect 168294 222000 168914 241398
rect 186294 259954 186914 278000
rect 186294 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 186914 259954
rect 186294 259634 186914 259718
rect 186294 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 186914 259634
rect 186294 223954 186914 259398
rect 186294 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 186914 223954
rect 186294 223634 186914 223718
rect 186294 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 186914 223634
rect 186294 222000 186914 223398
rect 190794 264454 191414 278000
rect 190794 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 191414 264454
rect 190794 264134 191414 264218
rect 190794 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 191414 264134
rect 190794 228454 191414 263898
rect 190794 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 191414 228454
rect 190794 228134 191414 228218
rect 190794 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 191414 228134
rect 190794 222000 191414 227898
rect 195294 268954 195914 278000
rect 195294 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 195914 268954
rect 195294 268634 195914 268718
rect 195294 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 195914 268634
rect 195294 232954 195914 268398
rect 195294 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 195914 232954
rect 195294 232634 195914 232718
rect 195294 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 195914 232634
rect 195294 222000 195914 232398
rect 199794 273454 200414 278000
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 222000 200414 236898
rect 204294 277954 204914 278000
rect 204294 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 204914 277954
rect 204294 277634 204914 277718
rect 204294 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 204914 277634
rect 204294 241954 204914 277398
rect 204294 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 204914 241954
rect 204294 241634 204914 241718
rect 204294 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 204914 241634
rect 204294 222000 204914 241398
rect 222294 259954 222914 278000
rect 222294 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 222914 259954
rect 222294 259634 222914 259718
rect 222294 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 222914 259634
rect 222294 223954 222914 259398
rect 222294 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 222914 223954
rect 222294 223634 222914 223718
rect 222294 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 222914 223634
rect 222294 222000 222914 223398
rect 226794 264454 227414 278000
rect 226794 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 227414 264454
rect 226794 264134 227414 264218
rect 226794 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 227414 264134
rect 226794 228454 227414 263898
rect 226794 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 227414 228454
rect 226794 228134 227414 228218
rect 226794 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 227414 228134
rect 226794 192454 227414 227898
rect 226794 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 227414 192454
rect 226794 192134 227414 192218
rect 226794 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 227414 192134
rect 79568 187954 79888 187986
rect 79568 187718 79610 187954
rect 79846 187718 79888 187954
rect 79568 187634 79888 187718
rect 79568 187398 79610 187634
rect 79846 187398 79888 187634
rect 79568 187366 79888 187398
rect 110288 187954 110608 187986
rect 110288 187718 110330 187954
rect 110566 187718 110608 187954
rect 110288 187634 110608 187718
rect 110288 187398 110330 187634
rect 110566 187398 110608 187634
rect 110288 187366 110608 187398
rect 141008 187954 141328 187986
rect 141008 187718 141050 187954
rect 141286 187718 141328 187954
rect 141008 187634 141328 187718
rect 141008 187398 141050 187634
rect 141286 187398 141328 187634
rect 141008 187366 141328 187398
rect 171728 187954 172048 187986
rect 171728 187718 171770 187954
rect 172006 187718 172048 187954
rect 171728 187634 172048 187718
rect 171728 187398 171770 187634
rect 172006 187398 172048 187634
rect 171728 187366 172048 187398
rect 202448 187954 202768 187986
rect 202448 187718 202490 187954
rect 202726 187718 202768 187954
rect 202448 187634 202768 187718
rect 202448 187398 202490 187634
rect 202726 187398 202768 187634
rect 202448 187366 202768 187398
rect 64208 183454 64528 183486
rect 64208 183218 64250 183454
rect 64486 183218 64528 183454
rect 64208 183134 64528 183218
rect 64208 182898 64250 183134
rect 64486 182898 64528 183134
rect 64208 182866 64528 182898
rect 94928 183454 95248 183486
rect 94928 183218 94970 183454
rect 95206 183218 95248 183454
rect 94928 183134 95248 183218
rect 94928 182898 94970 183134
rect 95206 182898 95248 183134
rect 94928 182866 95248 182898
rect 125648 183454 125968 183486
rect 125648 183218 125690 183454
rect 125926 183218 125968 183454
rect 125648 183134 125968 183218
rect 125648 182898 125690 183134
rect 125926 182898 125968 183134
rect 125648 182866 125968 182898
rect 156368 183454 156688 183486
rect 156368 183218 156410 183454
rect 156646 183218 156688 183454
rect 156368 183134 156688 183218
rect 156368 182898 156410 183134
rect 156646 182898 156688 183134
rect 156368 182866 156688 182898
rect 187088 183454 187408 183486
rect 187088 183218 187130 183454
rect 187366 183218 187408 183454
rect 187088 183134 187408 183218
rect 187088 182898 187130 183134
rect 187366 182898 187408 183134
rect 187088 182866 187408 182898
rect 217808 183454 218128 183486
rect 217808 183218 217850 183454
rect 218086 183218 218128 183454
rect 217808 183134 218128 183218
rect 217808 182898 217850 183134
rect 218086 182898 218128 183134
rect 217808 182866 218128 182898
rect 226794 156454 227414 191898
rect 226794 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 227414 156454
rect 226794 156134 227414 156218
rect 226794 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 227414 156134
rect 79568 151954 79888 151986
rect 79568 151718 79610 151954
rect 79846 151718 79888 151954
rect 79568 151634 79888 151718
rect 79568 151398 79610 151634
rect 79846 151398 79888 151634
rect 79568 151366 79888 151398
rect 110288 151954 110608 151986
rect 110288 151718 110330 151954
rect 110566 151718 110608 151954
rect 110288 151634 110608 151718
rect 110288 151398 110330 151634
rect 110566 151398 110608 151634
rect 110288 151366 110608 151398
rect 141008 151954 141328 151986
rect 141008 151718 141050 151954
rect 141286 151718 141328 151954
rect 141008 151634 141328 151718
rect 141008 151398 141050 151634
rect 141286 151398 141328 151634
rect 141008 151366 141328 151398
rect 171728 151954 172048 151986
rect 171728 151718 171770 151954
rect 172006 151718 172048 151954
rect 171728 151634 172048 151718
rect 171728 151398 171770 151634
rect 172006 151398 172048 151634
rect 171728 151366 172048 151398
rect 202448 151954 202768 151986
rect 202448 151718 202490 151954
rect 202726 151718 202768 151954
rect 202448 151634 202768 151718
rect 202448 151398 202490 151634
rect 202726 151398 202768 151634
rect 202448 151366 202768 151398
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 57835 131748 57901 131749
rect 57835 131684 57836 131748
rect 57900 131684 57901 131748
rect 57835 131683 57901 131684
rect 51294 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 51914 124954
rect 51294 124634 51914 124718
rect 51294 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 51914 124634
rect 51294 88954 51914 124398
rect 226794 120454 227414 155898
rect 226794 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 227414 120454
rect 226794 120134 227414 120218
rect 226794 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 227414 120134
rect 79568 115954 79888 115986
rect 79568 115718 79610 115954
rect 79846 115718 79888 115954
rect 79568 115634 79888 115718
rect 79568 115398 79610 115634
rect 79846 115398 79888 115634
rect 79568 115366 79888 115398
rect 110288 115954 110608 115986
rect 110288 115718 110330 115954
rect 110566 115718 110608 115954
rect 110288 115634 110608 115718
rect 110288 115398 110330 115634
rect 110566 115398 110608 115634
rect 110288 115366 110608 115398
rect 141008 115954 141328 115986
rect 141008 115718 141050 115954
rect 141286 115718 141328 115954
rect 141008 115634 141328 115718
rect 141008 115398 141050 115634
rect 141286 115398 141328 115634
rect 141008 115366 141328 115398
rect 171728 115954 172048 115986
rect 171728 115718 171770 115954
rect 172006 115718 172048 115954
rect 171728 115634 172048 115718
rect 171728 115398 171770 115634
rect 172006 115398 172048 115634
rect 171728 115366 172048 115398
rect 202448 115954 202768 115986
rect 202448 115718 202490 115954
rect 202726 115718 202768 115954
rect 202448 115634 202768 115718
rect 202448 115398 202490 115634
rect 202726 115398 202768 115634
rect 202448 115366 202768 115398
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 51294 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 51914 88954
rect 51294 88634 51914 88718
rect 51294 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 51914 88634
rect 51294 52954 51914 88398
rect 226794 84454 227414 119898
rect 226794 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 227414 84454
rect 226794 84134 227414 84218
rect 226794 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 227414 84134
rect 79568 79954 79888 79986
rect 79568 79718 79610 79954
rect 79846 79718 79888 79954
rect 79568 79634 79888 79718
rect 79568 79398 79610 79634
rect 79846 79398 79888 79634
rect 79568 79366 79888 79398
rect 110288 79954 110608 79986
rect 110288 79718 110330 79954
rect 110566 79718 110608 79954
rect 110288 79634 110608 79718
rect 110288 79398 110330 79634
rect 110566 79398 110608 79634
rect 110288 79366 110608 79398
rect 141008 79954 141328 79986
rect 141008 79718 141050 79954
rect 141286 79718 141328 79954
rect 141008 79634 141328 79718
rect 141008 79398 141050 79634
rect 141286 79398 141328 79634
rect 141008 79366 141328 79398
rect 171728 79954 172048 79986
rect 171728 79718 171770 79954
rect 172006 79718 172048 79954
rect 171728 79634 172048 79718
rect 171728 79398 171770 79634
rect 172006 79398 172048 79634
rect 171728 79366 172048 79398
rect 202448 79954 202768 79986
rect 202448 79718 202490 79954
rect 202726 79718 202768 79954
rect 202448 79634 202768 79718
rect 202448 79398 202490 79634
rect 202726 79398 202768 79634
rect 202448 79366 202768 79398
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 51294 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 51914 52954
rect 51294 52634 51914 52718
rect 51294 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 51914 52634
rect 51294 16954 51914 52398
rect 51294 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 51914 16954
rect 51294 16634 51914 16718
rect 51294 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 51914 16634
rect 51294 -3226 51914 16398
rect 51294 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 51914 -3226
rect 51294 -3546 51914 -3462
rect 51294 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 51914 -3546
rect 51294 -7654 51914 -3782
rect 55794 57454 56414 58000
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -4186 56414 20898
rect 55794 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 56414 -4186
rect 55794 -4506 56414 -4422
rect 55794 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 56414 -4506
rect 55794 -7654 56414 -4742
rect 60294 25954 60914 58000
rect 60294 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 60914 25954
rect 60294 25634 60914 25718
rect 60294 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 60914 25634
rect 60294 -5146 60914 25398
rect 60294 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 60914 -5146
rect 60294 -5466 60914 -5382
rect 60294 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 60914 -5466
rect 60294 -7654 60914 -5702
rect 64794 30454 65414 58000
rect 64794 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 65414 30454
rect 64794 30134 65414 30218
rect 64794 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 65414 30134
rect 64794 -6106 65414 29898
rect 64794 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 65414 -6106
rect 64794 -6426 65414 -6342
rect 64794 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 65414 -6426
rect 64794 -7654 65414 -6662
rect 69294 34954 69914 58000
rect 69294 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 69914 34954
rect 69294 34634 69914 34718
rect 69294 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 69914 34634
rect 69294 -7066 69914 34398
rect 69294 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 69914 -7066
rect 69294 -7386 69914 -7302
rect 69294 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 69914 -7386
rect 69294 -7654 69914 -7622
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 78294 43954 78914 58000
rect 78294 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 78914 43954
rect 78294 43634 78914 43718
rect 78294 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 78914 43634
rect 78294 7954 78914 43398
rect 78294 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 78914 7954
rect 78294 7634 78914 7718
rect 78294 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 78914 7634
rect 78294 -1306 78914 7398
rect 78294 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 78914 -1306
rect 78294 -1626 78914 -1542
rect 78294 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 78914 -1626
rect 78294 -7654 78914 -1862
rect 82794 48454 83414 58000
rect 82794 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 83414 48454
rect 82794 48134 83414 48218
rect 82794 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 83414 48134
rect 82794 12454 83414 47898
rect 82794 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 83414 12454
rect 82794 12134 83414 12218
rect 82794 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 83414 12134
rect 82794 -2266 83414 11898
rect 82794 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 83414 -2266
rect 82794 -2586 83414 -2502
rect 82794 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 83414 -2586
rect 82794 -7654 83414 -2822
rect 87294 52954 87914 58000
rect 87294 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 87914 52954
rect 87294 52634 87914 52718
rect 87294 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 87914 52634
rect 87294 16954 87914 52398
rect 87294 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 87914 16954
rect 87294 16634 87914 16718
rect 87294 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 87914 16634
rect 87294 -3226 87914 16398
rect 87294 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 87914 -3226
rect 87294 -3546 87914 -3462
rect 87294 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 87914 -3546
rect 87294 -7654 87914 -3782
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -4186 92414 20898
rect 91794 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 92414 -4186
rect 91794 -4506 92414 -4422
rect 91794 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 92414 -4506
rect 91794 -7654 92414 -4742
rect 96294 25954 96914 58000
rect 96294 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 96914 25954
rect 96294 25634 96914 25718
rect 96294 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 96914 25634
rect 96294 -5146 96914 25398
rect 96294 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 96914 -5146
rect 96294 -5466 96914 -5382
rect 96294 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 96914 -5466
rect 96294 -7654 96914 -5702
rect 100794 30454 101414 58000
rect 100794 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 101414 30454
rect 100794 30134 101414 30218
rect 100794 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 101414 30134
rect 100794 -6106 101414 29898
rect 100794 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 101414 -6106
rect 100794 -6426 101414 -6342
rect 100794 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 101414 -6426
rect 100794 -7654 101414 -6662
rect 105294 34954 105914 58000
rect 105294 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 105914 34954
rect 105294 34634 105914 34718
rect 105294 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 105914 34634
rect 105294 -7066 105914 34398
rect 105294 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 105914 -7066
rect 105294 -7386 105914 -7302
rect 105294 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 105914 -7386
rect 105294 -7654 105914 -7622
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 114294 43954 114914 58000
rect 114294 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 114914 43954
rect 114294 43634 114914 43718
rect 114294 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 114914 43634
rect 114294 7954 114914 43398
rect 114294 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 114914 7954
rect 114294 7634 114914 7718
rect 114294 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 114914 7634
rect 114294 -1306 114914 7398
rect 114294 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 114914 -1306
rect 114294 -1626 114914 -1542
rect 114294 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 114914 -1626
rect 114294 -7654 114914 -1862
rect 118794 48454 119414 58000
rect 118794 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 119414 48454
rect 118794 48134 119414 48218
rect 118794 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 119414 48134
rect 118794 12454 119414 47898
rect 118794 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 119414 12454
rect 118794 12134 119414 12218
rect 118794 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 119414 12134
rect 118794 -2266 119414 11898
rect 118794 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 119414 -2266
rect 118794 -2586 119414 -2502
rect 118794 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 119414 -2586
rect 118794 -7654 119414 -2822
rect 123294 52954 123914 58000
rect 123294 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 123914 52954
rect 123294 52634 123914 52718
rect 123294 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 123914 52634
rect 123294 16954 123914 52398
rect 123294 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 123914 16954
rect 123294 16634 123914 16718
rect 123294 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 123914 16634
rect 123294 -3226 123914 16398
rect 123294 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 123914 -3226
rect 123294 -3546 123914 -3462
rect 123294 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 123914 -3546
rect 123294 -7654 123914 -3782
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -4186 128414 20898
rect 127794 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 128414 -4186
rect 127794 -4506 128414 -4422
rect 127794 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 128414 -4506
rect 127794 -7654 128414 -4742
rect 132294 25954 132914 58000
rect 132294 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 132914 25954
rect 132294 25634 132914 25718
rect 132294 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 132914 25634
rect 132294 -5146 132914 25398
rect 132294 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 132914 -5146
rect 132294 -5466 132914 -5382
rect 132294 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 132914 -5466
rect 132294 -7654 132914 -5702
rect 136794 30454 137414 58000
rect 136794 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 137414 30454
rect 136794 30134 137414 30218
rect 136794 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 137414 30134
rect 136794 -6106 137414 29898
rect 136794 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 137414 -6106
rect 136794 -6426 137414 -6342
rect 136794 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 137414 -6426
rect 136794 -7654 137414 -6662
rect 141294 34954 141914 58000
rect 141294 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 141914 34954
rect 141294 34634 141914 34718
rect 141294 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 141914 34634
rect 141294 -7066 141914 34398
rect 141294 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 141914 -7066
rect 141294 -7386 141914 -7302
rect 141294 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 141914 -7386
rect 141294 -7654 141914 -7622
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 150294 43954 150914 58000
rect 150294 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 150914 43954
rect 150294 43634 150914 43718
rect 150294 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 150914 43634
rect 150294 7954 150914 43398
rect 150294 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 150914 7954
rect 150294 7634 150914 7718
rect 150294 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 150914 7634
rect 150294 -1306 150914 7398
rect 150294 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 150914 -1306
rect 150294 -1626 150914 -1542
rect 150294 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 150914 -1626
rect 150294 -7654 150914 -1862
rect 154794 48454 155414 58000
rect 154794 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 155414 48454
rect 154794 48134 155414 48218
rect 154794 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 155414 48134
rect 154794 12454 155414 47898
rect 154794 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 155414 12454
rect 154794 12134 155414 12218
rect 154794 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 155414 12134
rect 154794 -2266 155414 11898
rect 154794 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 155414 -2266
rect 154794 -2586 155414 -2502
rect 154794 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 155414 -2586
rect 154794 -7654 155414 -2822
rect 159294 52954 159914 58000
rect 159294 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 159914 52954
rect 159294 52634 159914 52718
rect 159294 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 159914 52634
rect 159294 16954 159914 52398
rect 159294 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 159914 16954
rect 159294 16634 159914 16718
rect 159294 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 159914 16634
rect 159294 -3226 159914 16398
rect 159294 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 159914 -3226
rect 159294 -3546 159914 -3462
rect 159294 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 159914 -3546
rect 159294 -7654 159914 -3782
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -4186 164414 20898
rect 163794 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 164414 -4186
rect 163794 -4506 164414 -4422
rect 163794 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 164414 -4506
rect 163794 -7654 164414 -4742
rect 168294 25954 168914 58000
rect 168294 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 168914 25954
rect 168294 25634 168914 25718
rect 168294 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 168914 25634
rect 168294 -5146 168914 25398
rect 168294 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 168914 -5146
rect 168294 -5466 168914 -5382
rect 168294 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 168914 -5466
rect 168294 -7654 168914 -5702
rect 172794 30454 173414 58000
rect 172794 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 173414 30454
rect 172794 30134 173414 30218
rect 172794 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 173414 30134
rect 172794 -6106 173414 29898
rect 172794 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 173414 -6106
rect 172794 -6426 173414 -6342
rect 172794 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 173414 -6426
rect 172794 -7654 173414 -6662
rect 177294 34954 177914 58000
rect 177294 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 177914 34954
rect 177294 34634 177914 34718
rect 177294 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 177914 34634
rect 177294 -7066 177914 34398
rect 177294 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 177914 -7066
rect 177294 -7386 177914 -7302
rect 177294 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 177914 -7386
rect 177294 -7654 177914 -7622
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 186294 43954 186914 58000
rect 186294 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 186914 43954
rect 186294 43634 186914 43718
rect 186294 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 186914 43634
rect 186294 7954 186914 43398
rect 186294 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 186914 7954
rect 186294 7634 186914 7718
rect 186294 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 186914 7634
rect 186294 -1306 186914 7398
rect 186294 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 186914 -1306
rect 186294 -1626 186914 -1542
rect 186294 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 186914 -1626
rect 186294 -7654 186914 -1862
rect 190794 48454 191414 58000
rect 190794 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 191414 48454
rect 190794 48134 191414 48218
rect 190794 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 191414 48134
rect 190794 12454 191414 47898
rect 190794 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 191414 12454
rect 190794 12134 191414 12218
rect 190794 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 191414 12134
rect 190794 -2266 191414 11898
rect 190794 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 191414 -2266
rect 190794 -2586 191414 -2502
rect 190794 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 191414 -2586
rect 190794 -7654 191414 -2822
rect 195294 52954 195914 58000
rect 195294 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 195914 52954
rect 195294 52634 195914 52718
rect 195294 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 195914 52634
rect 195294 16954 195914 52398
rect 195294 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 195914 16954
rect 195294 16634 195914 16718
rect 195294 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 195914 16634
rect 195294 -3226 195914 16398
rect 195294 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 195914 -3226
rect 195294 -3546 195914 -3462
rect 195294 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 195914 -3546
rect 195294 -7654 195914 -3782
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -4186 200414 20898
rect 199794 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 200414 -4186
rect 199794 -4506 200414 -4422
rect 199794 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 200414 -4506
rect 199794 -7654 200414 -4742
rect 204294 25954 204914 58000
rect 204294 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 204914 25954
rect 204294 25634 204914 25718
rect 204294 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 204914 25634
rect 204294 -5146 204914 25398
rect 204294 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 204914 -5146
rect 204294 -5466 204914 -5382
rect 204294 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 204914 -5466
rect 204294 -7654 204914 -5702
rect 208794 30454 209414 58000
rect 208794 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 209414 30454
rect 208794 30134 209414 30218
rect 208794 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 209414 30134
rect 208794 -6106 209414 29898
rect 208794 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 209414 -6106
rect 208794 -6426 209414 -6342
rect 208794 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 209414 -6426
rect 208794 -7654 209414 -6662
rect 213294 34954 213914 58000
rect 213294 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 213914 34954
rect 213294 34634 213914 34718
rect 213294 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 213914 34634
rect 213294 -7066 213914 34398
rect 213294 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 213914 -7066
rect 213294 -7386 213914 -7302
rect 213294 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 213914 -7386
rect 213294 -7654 213914 -7622
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 222294 43954 222914 58000
rect 222294 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 222914 43954
rect 222294 43634 222914 43718
rect 222294 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 222914 43634
rect 222294 7954 222914 43398
rect 222294 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 222914 7954
rect 222294 7634 222914 7718
rect 222294 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 222914 7634
rect 222294 -1306 222914 7398
rect 222294 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 222914 -1306
rect 222294 -1626 222914 -1542
rect 222294 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 222914 -1626
rect 222294 -7654 222914 -1862
rect 226794 48454 227414 83898
rect 226794 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 227414 48454
rect 226794 48134 227414 48218
rect 226794 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 227414 48134
rect 226794 12454 227414 47898
rect 226794 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 227414 12454
rect 226794 12134 227414 12218
rect 226794 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 227414 12134
rect 226794 -2266 227414 11898
rect 226794 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 227414 -2266
rect 226794 -2586 227414 -2502
rect 226794 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 227414 -2586
rect 226794 -7654 227414 -2822
rect 231294 268954 231914 278000
rect 231294 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 231914 268954
rect 231294 268634 231914 268718
rect 231294 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 231914 268634
rect 231294 232954 231914 268398
rect 231294 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 231914 232954
rect 231294 232634 231914 232718
rect 231294 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 231914 232634
rect 231294 196954 231914 232398
rect 231294 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 231914 196954
rect 231294 196634 231914 196718
rect 231294 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 231914 196634
rect 231294 160954 231914 196398
rect 231294 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 231914 160954
rect 231294 160634 231914 160718
rect 231294 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 231914 160634
rect 231294 124954 231914 160398
rect 231294 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 231914 124954
rect 231294 124634 231914 124718
rect 231294 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 231914 124634
rect 231294 88954 231914 124398
rect 231294 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 231914 88954
rect 231294 88634 231914 88718
rect 231294 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 231914 88634
rect 231294 52954 231914 88398
rect 231294 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 231914 52954
rect 231294 52634 231914 52718
rect 231294 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 231914 52634
rect 231294 16954 231914 52398
rect 231294 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 231914 16954
rect 231294 16634 231914 16718
rect 231294 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 231914 16634
rect 231294 -3226 231914 16398
rect 231294 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 231914 -3226
rect 231294 -3546 231914 -3462
rect 231294 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 231914 -3546
rect 231294 -7654 231914 -3782
rect 235794 273454 236414 278000
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -4186 236414 20898
rect 235794 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 236414 -4186
rect 235794 -4506 236414 -4422
rect 235794 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 236414 -4506
rect 235794 -7654 236414 -4742
rect 240294 277954 240914 278000
rect 240294 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 240914 277954
rect 240294 277634 240914 277718
rect 240294 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 240914 277634
rect 240294 241954 240914 277398
rect 240294 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 240914 241954
rect 240294 241634 240914 241718
rect 240294 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 240914 241634
rect 240294 205954 240914 241398
rect 240294 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 240914 205954
rect 240294 205634 240914 205718
rect 240294 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 240914 205634
rect 240294 169954 240914 205398
rect 240294 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 240914 169954
rect 240294 169634 240914 169718
rect 240294 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 240914 169634
rect 240294 133954 240914 169398
rect 240294 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 240914 133954
rect 240294 133634 240914 133718
rect 240294 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 240914 133634
rect 240294 97954 240914 133398
rect 240294 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 240914 97954
rect 240294 97634 240914 97718
rect 240294 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 240914 97634
rect 240294 61954 240914 97398
rect 240294 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 240914 61954
rect 240294 61634 240914 61718
rect 240294 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 240914 61634
rect 240294 25954 240914 61398
rect 240294 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 240914 25954
rect 240294 25634 240914 25718
rect 240294 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 240914 25634
rect 240294 -5146 240914 25398
rect 240294 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 240914 -5146
rect 240294 -5466 240914 -5382
rect 240294 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 240914 -5466
rect 240294 -7654 240914 -5702
rect 244794 246454 245414 278000
rect 244794 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 245414 246454
rect 244794 246134 245414 246218
rect 244794 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 245414 246134
rect 244794 210454 245414 245898
rect 244794 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 245414 210454
rect 244794 210134 245414 210218
rect 244794 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 245414 210134
rect 244794 174454 245414 209898
rect 244794 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 245414 174454
rect 244794 174134 245414 174218
rect 244794 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 245414 174134
rect 244794 138454 245414 173898
rect 244794 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 245414 138454
rect 244794 138134 245414 138218
rect 244794 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 245414 138134
rect 244794 102454 245414 137898
rect 244794 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 245414 102454
rect 244794 102134 245414 102218
rect 244794 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 245414 102134
rect 244794 66454 245414 101898
rect 244794 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 245414 66454
rect 244794 66134 245414 66218
rect 244794 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 245414 66134
rect 244794 30454 245414 65898
rect 244794 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 245414 30454
rect 244794 30134 245414 30218
rect 244794 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 245414 30134
rect 244794 -6106 245414 29898
rect 244794 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 245414 -6106
rect 244794 -6426 245414 -6342
rect 244794 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 245414 -6426
rect 244794 -7654 245414 -6662
rect 249294 250954 249914 278000
rect 249294 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 249914 250954
rect 249294 250634 249914 250718
rect 249294 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 249914 250634
rect 249294 214954 249914 250398
rect 249294 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 249914 214954
rect 249294 214634 249914 214718
rect 249294 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 249914 214634
rect 249294 178954 249914 214398
rect 249294 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 249914 178954
rect 249294 178634 249914 178718
rect 249294 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 249914 178634
rect 249294 142954 249914 178398
rect 249294 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 249914 142954
rect 249294 142634 249914 142718
rect 249294 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 249914 142634
rect 249294 106954 249914 142398
rect 249294 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 249914 106954
rect 249294 106634 249914 106718
rect 249294 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 249914 106634
rect 249294 70954 249914 106398
rect 249294 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 249914 70954
rect 249294 70634 249914 70718
rect 249294 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 249914 70634
rect 249294 34954 249914 70398
rect 249294 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 249914 34954
rect 249294 34634 249914 34718
rect 249294 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 249914 34634
rect 249294 -7066 249914 34398
rect 249294 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 249914 -7066
rect 249294 -7386 249914 -7302
rect 249294 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 249914 -7386
rect 249294 -7654 249914 -7622
rect 253794 255454 254414 278000
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 258294 259954 258914 295398
rect 258294 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 258914 259954
rect 258294 259634 258914 259718
rect 258294 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 258914 259634
rect 258294 223954 258914 259398
rect 258294 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 258914 223954
rect 258294 223634 258914 223718
rect 258294 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 258914 223634
rect 258294 187954 258914 223398
rect 258294 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 258914 187954
rect 258294 187634 258914 187718
rect 258294 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 258914 187634
rect 258294 151954 258914 187398
rect 258294 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 258914 151954
rect 258294 151634 258914 151718
rect 258294 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 258914 151634
rect 258294 115954 258914 151398
rect 258294 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 258914 115954
rect 258294 115634 258914 115718
rect 258294 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 258914 115634
rect 258294 79954 258914 115398
rect 258294 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 258914 79954
rect 258294 79634 258914 79718
rect 258294 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 258914 79634
rect 258294 43954 258914 79398
rect 258294 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 258914 43954
rect 258294 43634 258914 43718
rect 258294 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 258914 43634
rect 258294 7954 258914 43398
rect 258294 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 258914 7954
rect 258294 7634 258914 7718
rect 258294 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 258914 7634
rect 258294 -1306 258914 7398
rect 258294 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 258914 -1306
rect 258294 -1626 258914 -1542
rect 258294 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 258914 -1626
rect 258294 -7654 258914 -1862
rect 262794 706758 263414 711590
rect 262794 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 263414 706758
rect 262794 706438 263414 706522
rect 262794 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 263414 706438
rect 262794 696454 263414 706202
rect 262794 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 263414 696454
rect 262794 696134 263414 696218
rect 262794 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 263414 696134
rect 262794 660454 263414 695898
rect 262794 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 263414 660454
rect 262794 660134 263414 660218
rect 262794 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 263414 660134
rect 262794 624454 263414 659898
rect 262794 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 263414 624454
rect 262794 624134 263414 624218
rect 262794 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 263414 624134
rect 262794 588454 263414 623898
rect 262794 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 263414 588454
rect 262794 588134 263414 588218
rect 262794 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 263414 588134
rect 262794 552454 263414 587898
rect 262794 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 263414 552454
rect 262794 552134 263414 552218
rect 262794 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 263414 552134
rect 262794 516454 263414 551898
rect 262794 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 263414 516454
rect 262794 516134 263414 516218
rect 262794 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 263414 516134
rect 262794 480454 263414 515898
rect 262794 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 263414 480454
rect 262794 480134 263414 480218
rect 262794 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 263414 480134
rect 262794 444454 263414 479898
rect 262794 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 263414 444454
rect 262794 444134 263414 444218
rect 262794 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 263414 444134
rect 262794 408454 263414 443898
rect 262794 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 263414 408454
rect 262794 408134 263414 408218
rect 262794 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 263414 408134
rect 262794 372454 263414 407898
rect 262794 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 263414 372454
rect 262794 372134 263414 372218
rect 262794 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 263414 372134
rect 262794 336454 263414 371898
rect 262794 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 263414 336454
rect 262794 336134 263414 336218
rect 262794 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 263414 336134
rect 262794 300454 263414 335898
rect 262794 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 263414 300454
rect 262794 300134 263414 300218
rect 262794 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 263414 300134
rect 262794 264454 263414 299898
rect 262794 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 263414 264454
rect 262794 264134 263414 264218
rect 262794 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 263414 264134
rect 262794 228454 263414 263898
rect 262794 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 263414 228454
rect 262794 228134 263414 228218
rect 262794 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 263414 228134
rect 262794 192454 263414 227898
rect 262794 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 263414 192454
rect 262794 192134 263414 192218
rect 262794 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 263414 192134
rect 262794 156454 263414 191898
rect 262794 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 263414 156454
rect 262794 156134 263414 156218
rect 262794 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 263414 156134
rect 262794 120454 263414 155898
rect 262794 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 263414 120454
rect 262794 120134 263414 120218
rect 262794 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 263414 120134
rect 262794 84454 263414 119898
rect 262794 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 263414 84454
rect 262794 84134 263414 84218
rect 262794 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 263414 84134
rect 262794 48454 263414 83898
rect 262794 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 263414 48454
rect 262794 48134 263414 48218
rect 262794 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 263414 48134
rect 262794 12454 263414 47898
rect 262794 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 263414 12454
rect 262794 12134 263414 12218
rect 262794 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 263414 12134
rect 262794 -2266 263414 11898
rect 262794 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 263414 -2266
rect 262794 -2586 263414 -2502
rect 262794 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 263414 -2586
rect 262794 -7654 263414 -2822
rect 267294 707718 267914 711590
rect 267294 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 267914 707718
rect 267294 707398 267914 707482
rect 267294 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 267914 707398
rect 267294 700954 267914 707162
rect 267294 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 267914 700954
rect 267294 700634 267914 700718
rect 267294 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 267914 700634
rect 267294 664954 267914 700398
rect 267294 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 267914 664954
rect 267294 664634 267914 664718
rect 267294 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 267914 664634
rect 267294 628954 267914 664398
rect 267294 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 267914 628954
rect 267294 628634 267914 628718
rect 267294 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 267914 628634
rect 267294 592954 267914 628398
rect 267294 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 267914 592954
rect 267294 592634 267914 592718
rect 267294 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 267914 592634
rect 267294 556954 267914 592398
rect 267294 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 267914 556954
rect 267294 556634 267914 556718
rect 267294 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 267914 556634
rect 267294 520954 267914 556398
rect 267294 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 267914 520954
rect 267294 520634 267914 520718
rect 267294 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 267914 520634
rect 267294 484954 267914 520398
rect 267294 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 267914 484954
rect 267294 484634 267914 484718
rect 267294 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 267914 484634
rect 267294 448954 267914 484398
rect 267294 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 267914 448954
rect 267294 448634 267914 448718
rect 267294 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 267914 448634
rect 267294 412954 267914 448398
rect 267294 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 267914 412954
rect 267294 412634 267914 412718
rect 267294 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 267914 412634
rect 267294 376954 267914 412398
rect 267294 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 267914 376954
rect 267294 376634 267914 376718
rect 267294 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 267914 376634
rect 267294 340954 267914 376398
rect 267294 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 267914 340954
rect 267294 340634 267914 340718
rect 267294 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 267914 340634
rect 267294 304954 267914 340398
rect 267294 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 267914 304954
rect 267294 304634 267914 304718
rect 267294 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 267914 304634
rect 267294 268954 267914 304398
rect 267294 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 267914 268954
rect 267294 268634 267914 268718
rect 267294 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 267914 268634
rect 267294 232954 267914 268398
rect 267294 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 267914 232954
rect 267294 232634 267914 232718
rect 267294 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 267914 232634
rect 267294 196954 267914 232398
rect 267294 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 267914 196954
rect 267294 196634 267914 196718
rect 267294 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 267914 196634
rect 267294 160954 267914 196398
rect 267294 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 267914 160954
rect 267294 160634 267914 160718
rect 267294 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 267914 160634
rect 267294 124954 267914 160398
rect 267294 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 267914 124954
rect 267294 124634 267914 124718
rect 267294 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 267914 124634
rect 267294 88954 267914 124398
rect 267294 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 267914 88954
rect 267294 88634 267914 88718
rect 267294 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 267914 88634
rect 267294 52954 267914 88398
rect 267294 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 267914 52954
rect 267294 52634 267914 52718
rect 267294 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 267914 52634
rect 267294 16954 267914 52398
rect 267294 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 267914 16954
rect 267294 16634 267914 16718
rect 267294 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 267914 16634
rect 267294 -3226 267914 16398
rect 267294 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 267914 -3226
rect 267294 -3546 267914 -3462
rect 267294 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 267914 -3546
rect 267294 -7654 267914 -3782
rect 271794 708678 272414 711590
rect 271794 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 272414 708678
rect 271794 708358 272414 708442
rect 271794 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 272414 708358
rect 271794 669454 272414 708122
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 276294 709638 276914 711590
rect 276294 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 276914 709638
rect 276294 709318 276914 709402
rect 276294 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 276914 709318
rect 276294 673954 276914 709082
rect 276294 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 276914 673954
rect 276294 673634 276914 673718
rect 276294 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 276914 673634
rect 276294 642000 276914 673398
rect 280794 710598 281414 711590
rect 280794 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 281414 710598
rect 280794 710278 281414 710362
rect 280794 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 281414 710278
rect 280794 678454 281414 710042
rect 280794 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 281414 678454
rect 280794 678134 281414 678218
rect 280794 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 281414 678134
rect 279371 660652 279437 660653
rect 279371 660588 279372 660652
rect 279436 660588 279437 660652
rect 279371 660587 279437 660588
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 279374 543149 279434 660587
rect 280794 642361 281414 677898
rect 285294 711558 285914 711590
rect 285294 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 285914 711558
rect 285294 711238 285914 711322
rect 285294 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 285914 711238
rect 285294 682954 285914 711002
rect 285294 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 285914 682954
rect 285294 682634 285914 682718
rect 285294 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 285914 682634
rect 283419 663236 283485 663237
rect 283419 663172 283420 663236
rect 283484 663172 283485 663236
rect 283419 663171 283485 663172
rect 282315 661876 282381 661877
rect 282315 661812 282316 661876
rect 282380 661812 282381 661876
rect 282315 661811 282381 661812
rect 280794 642125 280826 642361
rect 281062 642125 281146 642361
rect 281382 642125 281414 642361
rect 280794 642000 281414 642125
rect 279371 543148 279437 543149
rect 279371 543084 279372 543148
rect 279436 543084 279437 543148
rect 279371 543083 279437 543084
rect 282318 543013 282378 661811
rect 283422 543285 283482 663171
rect 285294 646954 285914 682398
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 286179 662964 286245 662965
rect 286179 662900 286180 662964
rect 286244 662900 286245 662964
rect 286179 662899 286245 662900
rect 285294 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 285914 646954
rect 285294 646634 285914 646718
rect 285294 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 285914 646634
rect 285294 642000 285914 646398
rect 285443 639300 285509 639301
rect 285443 639236 285444 639300
rect 285508 639236 285509 639300
rect 285443 639235 285509 639236
rect 284208 615454 284528 615486
rect 284208 615218 284250 615454
rect 284486 615218 284528 615454
rect 284208 615134 284528 615218
rect 284208 614898 284250 615134
rect 284486 614898 284528 615134
rect 284208 614866 284528 614898
rect 285446 560965 285506 639235
rect 285443 560964 285509 560965
rect 285443 560900 285444 560964
rect 285508 560900 285509 560964
rect 285443 560899 285509 560900
rect 286182 543421 286242 662899
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 642000 290414 650898
rect 294294 705798 294914 711590
rect 294294 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 294914 705798
rect 294294 705478 294914 705562
rect 294294 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 294914 705478
rect 294294 691954 294914 705242
rect 294294 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 294914 691954
rect 294294 691634 294914 691718
rect 294294 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 294914 691634
rect 294294 655954 294914 691398
rect 298794 706758 299414 711590
rect 298794 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 299414 706758
rect 298794 706438 299414 706522
rect 298794 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 299414 706438
rect 298794 696454 299414 706202
rect 298794 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 299414 696454
rect 298794 696134 299414 696218
rect 298794 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 299414 696134
rect 295011 661740 295077 661741
rect 295011 661676 295012 661740
rect 295076 661676 295077 661740
rect 295011 661675 295077 661676
rect 294294 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 294914 655954
rect 294294 655634 294914 655718
rect 294294 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 294914 655634
rect 294294 642000 294914 655398
rect 288203 639300 288269 639301
rect 288203 639236 288204 639300
rect 288268 639236 288269 639300
rect 288203 639235 288269 639236
rect 289491 639300 289557 639301
rect 289491 639236 289492 639300
rect 289556 639236 289557 639300
rect 289491 639235 289557 639236
rect 290963 639300 291029 639301
rect 290963 639236 290964 639300
rect 291028 639236 291029 639300
rect 290963 639235 291029 639236
rect 292435 639300 292501 639301
rect 292435 639236 292436 639300
rect 292500 639236 292501 639300
rect 292435 639235 292501 639236
rect 293723 639300 293789 639301
rect 293723 639236 293724 639300
rect 293788 639236 293789 639300
rect 293723 639235 293789 639236
rect 288206 558245 288266 639235
rect 289494 562325 289554 639235
rect 289794 579454 290414 598000
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289491 562324 289557 562325
rect 289491 562260 289492 562324
rect 289556 562260 289557 562324
rect 289491 562259 289557 562260
rect 288203 558244 288269 558245
rect 288203 558180 288204 558244
rect 288268 558180 288269 558244
rect 288203 558179 288269 558180
rect 289794 543454 290414 578898
rect 290966 569261 291026 639235
rect 292438 581637 292498 639235
rect 292435 581636 292501 581637
rect 292435 581572 292436 581636
rect 292500 581572 292501 581636
rect 292435 581571 292501 581572
rect 290963 569260 291029 569261
rect 290963 569196 290964 569260
rect 291028 569196 291029 569260
rect 290963 569195 291029 569196
rect 293726 551309 293786 639235
rect 294294 583954 294914 598000
rect 294294 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 294914 583954
rect 294294 583634 294914 583718
rect 294294 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 294914 583634
rect 293723 551308 293789 551309
rect 293723 551244 293724 551308
rect 293788 551244 293789 551308
rect 293723 551243 293789 551244
rect 286179 543420 286245 543421
rect 286179 543356 286180 543420
rect 286244 543356 286245 543420
rect 286179 543355 286245 543356
rect 283419 543284 283485 543285
rect 283419 543220 283420 543284
rect 283484 543220 283485 543284
rect 283419 543219 283485 543220
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 282315 543012 282381 543013
rect 282315 542948 282316 543012
rect 282380 542948 282381 543012
rect 282315 542947 282381 542948
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 282131 542740 282197 542741
rect 282131 542676 282132 542740
rect 282196 542676 282197 542740
rect 282131 542675 282197 542676
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -4186 272414 20898
rect 271794 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 272414 -4186
rect 271794 -4506 272414 -4422
rect 271794 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 272414 -4506
rect 271794 -7654 272414 -4742
rect 276294 493954 276914 498000
rect 276294 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 276914 493954
rect 276294 493634 276914 493718
rect 276294 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 276914 493634
rect 276294 457954 276914 493398
rect 276294 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 276914 457954
rect 276294 457634 276914 457718
rect 276294 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 276914 457634
rect 276294 421954 276914 457398
rect 276294 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 276914 421954
rect 276294 421634 276914 421718
rect 276294 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 276914 421634
rect 276294 385954 276914 421398
rect 276294 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 276914 385954
rect 276294 385634 276914 385718
rect 276294 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 276914 385634
rect 276294 349954 276914 385398
rect 276294 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 276914 349954
rect 276294 349634 276914 349718
rect 276294 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 276914 349634
rect 276294 313954 276914 349398
rect 276294 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 276914 313954
rect 276294 313634 276914 313718
rect 276294 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 276914 313634
rect 276294 277954 276914 313398
rect 276294 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 276914 277954
rect 276294 277634 276914 277718
rect 276294 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 276914 277634
rect 276294 241954 276914 277398
rect 276294 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 276914 241954
rect 276294 241634 276914 241718
rect 276294 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 276914 241634
rect 276294 205954 276914 241398
rect 276294 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 276914 205954
rect 276294 205634 276914 205718
rect 276294 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 276914 205634
rect 276294 169954 276914 205398
rect 276294 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 276914 169954
rect 276294 169634 276914 169718
rect 276294 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 276914 169634
rect 276294 133954 276914 169398
rect 276294 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 276914 133954
rect 276294 133634 276914 133718
rect 276294 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 276914 133634
rect 276294 97954 276914 133398
rect 276294 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 276914 97954
rect 276294 97634 276914 97718
rect 276294 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 276914 97634
rect 276294 61954 276914 97398
rect 276294 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 276914 61954
rect 276294 61634 276914 61718
rect 276294 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 276914 61634
rect 276294 25954 276914 61398
rect 276294 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 276914 25954
rect 276294 25634 276914 25718
rect 276294 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 276914 25634
rect 276294 -5146 276914 25398
rect 276294 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 276914 -5146
rect 276294 -5466 276914 -5382
rect 276294 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 276914 -5466
rect 276294 -7654 276914 -5702
rect 280794 462454 281414 498000
rect 280794 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 281414 462454
rect 280794 462134 281414 462218
rect 280794 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 281414 462134
rect 280794 426454 281414 461898
rect 280794 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 281414 426454
rect 280794 426134 281414 426218
rect 280794 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 281414 426134
rect 280794 390454 281414 425898
rect 280794 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 281414 390454
rect 280794 390134 281414 390218
rect 280794 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 281414 390134
rect 280794 354454 281414 389898
rect 280794 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 281414 354454
rect 280794 354134 281414 354218
rect 280794 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 281414 354134
rect 280794 318454 281414 353898
rect 280794 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 281414 318454
rect 280794 318134 281414 318218
rect 280794 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 281414 318134
rect 280794 282454 281414 317898
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 246454 281414 281898
rect 282134 280669 282194 542675
rect 289794 542000 290414 542898
rect 294294 547954 294914 583398
rect 294294 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 294914 547954
rect 294294 547634 294914 547718
rect 294294 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 294914 547634
rect 294294 542000 294914 547398
rect 295014 543557 295074 661675
rect 295931 661604 295997 661605
rect 295931 661540 295932 661604
rect 295996 661540 295997 661604
rect 295931 661539 295997 661540
rect 295934 543693 295994 661539
rect 297219 661468 297285 661469
rect 297219 661404 297220 661468
rect 297284 661404 297285 661468
rect 297219 661403 297285 661404
rect 295931 543692 295997 543693
rect 295931 543628 295932 543692
rect 295996 543628 295997 543692
rect 295931 543627 295997 543628
rect 295011 543556 295077 543557
rect 295011 543492 295012 543556
rect 295076 543492 295077 543556
rect 295011 543491 295077 543492
rect 297222 543421 297282 661403
rect 298794 660454 299414 695898
rect 298794 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 299414 660454
rect 298794 660134 299414 660218
rect 298794 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 299414 660134
rect 298794 642000 299414 659898
rect 303294 707718 303914 711590
rect 303294 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 303914 707718
rect 303294 707398 303914 707482
rect 303294 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 303914 707398
rect 303294 700954 303914 707162
rect 303294 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 303914 700954
rect 303294 700634 303914 700718
rect 303294 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 303914 700634
rect 303294 664954 303914 700398
rect 303294 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 303914 664954
rect 303294 664634 303914 664718
rect 303294 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 303914 664634
rect 303294 642000 303914 664398
rect 307794 708678 308414 711590
rect 307794 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 308414 708678
rect 307794 708358 308414 708442
rect 307794 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 308414 708358
rect 307794 669454 308414 708122
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 642000 308414 668898
rect 312294 709638 312914 711590
rect 312294 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 312914 709638
rect 312294 709318 312914 709402
rect 312294 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 312914 709318
rect 312294 673954 312914 709082
rect 312294 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 312914 673954
rect 312294 673634 312914 673718
rect 312294 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 312914 673634
rect 311019 661468 311085 661469
rect 311019 661404 311020 661468
rect 311084 661404 311085 661468
rect 311019 661403 311085 661404
rect 308627 661332 308693 661333
rect 308627 661268 308628 661332
rect 308692 661268 308693 661332
rect 308627 661267 308693 661268
rect 304763 641068 304829 641069
rect 304763 641004 304764 641068
rect 304828 641004 304829 641068
rect 304763 641003 304829 641004
rect 301451 640388 301517 640389
rect 301451 640324 301452 640388
rect 301516 640324 301517 640388
rect 301451 640323 301517 640324
rect 298507 639300 298573 639301
rect 298507 639236 298508 639300
rect 298572 639236 298573 639300
rect 298507 639235 298573 639236
rect 298510 561101 298570 639235
rect 300715 639164 300781 639165
rect 300715 639100 300716 639164
rect 300780 639100 300781 639164
rect 300715 639099 300781 639100
rect 299568 619954 299888 619986
rect 299568 619718 299610 619954
rect 299846 619718 299888 619954
rect 299568 619634 299888 619718
rect 299568 619398 299610 619634
rect 299846 619398 299888 619634
rect 299568 619366 299888 619398
rect 300718 600133 300778 639099
rect 300715 600132 300781 600133
rect 300715 600068 300716 600132
rect 300780 600068 300781 600132
rect 300715 600067 300781 600068
rect 301454 598909 301514 640323
rect 303475 639028 303541 639029
rect 303475 638964 303476 639028
rect 303540 638964 303541 639028
rect 303475 638963 303541 638964
rect 303478 600677 303538 638963
rect 304766 600677 304826 641003
rect 306235 640932 306301 640933
rect 306235 640868 306236 640932
rect 306300 640868 306301 640932
rect 306235 640867 306301 640868
rect 306238 600677 306298 640867
rect 306971 639300 307037 639301
rect 306971 639236 306972 639300
rect 307036 639236 307037 639300
rect 306971 639235 307037 639236
rect 303475 600676 303541 600677
rect 303475 600612 303476 600676
rect 303540 600612 303541 600676
rect 303475 600611 303541 600612
rect 304763 600676 304829 600677
rect 304763 600612 304764 600676
rect 304828 600612 304829 600676
rect 304763 600611 304829 600612
rect 306235 600676 306301 600677
rect 306235 600612 306236 600676
rect 306300 600612 306301 600676
rect 306235 600611 306301 600612
rect 306974 600541 307034 639235
rect 306971 600540 307037 600541
rect 306971 600476 306972 600540
rect 307036 600476 307037 600540
rect 306971 600475 307037 600476
rect 301451 598908 301517 598909
rect 301451 598844 301452 598908
rect 301516 598844 301517 598908
rect 301451 598843 301517 598844
rect 298794 588454 299414 598000
rect 298794 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 299414 588454
rect 298794 588134 299414 588218
rect 298794 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 299414 588134
rect 298507 561100 298573 561101
rect 298507 561036 298508 561100
rect 298572 561036 298573 561100
rect 298507 561035 298573 561036
rect 298794 552454 299414 587898
rect 298794 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 299414 552454
rect 298794 552134 299414 552218
rect 298794 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 299414 552134
rect 297219 543420 297285 543421
rect 297219 543356 297220 543420
rect 297284 543356 297285 543420
rect 297219 543355 297285 543356
rect 298794 542000 299414 551898
rect 303294 592954 303914 598000
rect 306974 597685 307034 600475
rect 306971 597684 307037 597685
rect 306971 597620 306972 597684
rect 307036 597620 307037 597684
rect 306971 597619 307037 597620
rect 303294 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 303914 592954
rect 303294 592634 303914 592718
rect 303294 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 303914 592634
rect 303294 556954 303914 592398
rect 303294 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 303914 556954
rect 303294 556634 303914 556718
rect 303294 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 303914 556634
rect 303294 542000 303914 556398
rect 307794 597454 308414 598000
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 542000 308414 560898
rect 308630 542469 308690 661267
rect 309363 661196 309429 661197
rect 309363 661132 309364 661196
rect 309428 661132 309429 661196
rect 309363 661131 309429 661132
rect 309179 661060 309245 661061
rect 309179 660996 309180 661060
rect 309244 660996 309245 661060
rect 309179 660995 309245 660996
rect 308811 660380 308877 660381
rect 308811 660316 308812 660380
rect 308876 660316 308877 660380
rect 308811 660315 308877 660316
rect 308814 542605 308874 660315
rect 308811 542604 308877 542605
rect 308811 542540 308812 542604
rect 308876 542540 308877 542604
rect 308811 542539 308877 542540
rect 309182 542469 309242 660995
rect 309366 542605 309426 661131
rect 310467 660244 310533 660245
rect 310467 660180 310468 660244
rect 310532 660180 310533 660244
rect 310467 660179 310533 660180
rect 310470 542605 310530 660179
rect 309363 542604 309429 542605
rect 309363 542540 309364 542604
rect 309428 542540 309429 542604
rect 309363 542539 309429 542540
rect 310467 542604 310533 542605
rect 310467 542540 310468 542604
rect 310532 542540 310533 542604
rect 310467 542539 310533 542540
rect 311022 542469 311082 661403
rect 311939 660108 312005 660109
rect 311939 660044 311940 660108
rect 312004 660044 312005 660108
rect 311939 660043 312005 660044
rect 311942 543149 312002 660043
rect 312294 642000 312914 673398
rect 316794 710598 317414 711590
rect 316794 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 317414 710598
rect 316794 710278 317414 710362
rect 316794 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 317414 710278
rect 316794 678454 317414 710042
rect 316794 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 317414 678454
rect 316794 678134 317414 678218
rect 316794 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 317414 678134
rect 316794 642361 317414 677898
rect 321294 711558 321914 711590
rect 321294 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 321914 711558
rect 321294 711238 321914 711322
rect 321294 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 321914 711238
rect 321294 682954 321914 711002
rect 321294 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 321914 682954
rect 321294 682634 321914 682718
rect 321294 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 321914 682634
rect 317643 662828 317709 662829
rect 317643 662764 317644 662828
rect 317708 662764 317709 662828
rect 317643 662763 317709 662764
rect 316794 642125 316826 642361
rect 317062 642125 317146 642361
rect 317382 642125 317414 642361
rect 316794 642000 317414 642125
rect 314928 615454 315248 615486
rect 314928 615218 314970 615454
rect 315206 615218 315248 615454
rect 314928 615134 315248 615218
rect 314928 614898 314970 615134
rect 315206 614898 315248 615134
rect 314928 614866 315248 614898
rect 317646 543693 317706 662763
rect 321294 646954 321914 682398
rect 321294 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 321914 646954
rect 321294 646634 321914 646718
rect 321294 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 321914 646634
rect 321294 642000 321914 646398
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 317643 543692 317709 543693
rect 317643 543628 317644 543692
rect 317708 543628 317709 543692
rect 317643 543627 317709 543628
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 311939 543148 312005 543149
rect 311939 543084 311940 543148
rect 312004 543084 312005 543148
rect 311939 543083 312005 543084
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 308627 542468 308693 542469
rect 308627 542404 308628 542468
rect 308692 542404 308693 542468
rect 308627 542403 308693 542404
rect 309179 542468 309245 542469
rect 309179 542404 309180 542468
rect 309244 542404 309245 542468
rect 309179 542403 309245 542404
rect 311019 542468 311085 542469
rect 311019 542404 311020 542468
rect 311084 542404 311085 542468
rect 311019 542403 311085 542404
rect 287283 539748 287349 539749
rect 287283 539684 287284 539748
rect 287348 539684 287349 539748
rect 287283 539683 287349 539684
rect 288571 539748 288637 539749
rect 288571 539684 288572 539748
rect 288636 539684 288637 539748
rect 288571 539683 288637 539684
rect 290595 539748 290661 539749
rect 290595 539684 290596 539748
rect 290660 539684 290661 539748
rect 290595 539683 290661 539684
rect 284891 539612 284957 539613
rect 284891 539548 284892 539612
rect 284956 539548 284957 539612
rect 284891 539547 284957 539548
rect 285995 539612 286061 539613
rect 285995 539548 285996 539612
rect 286060 539548 286061 539612
rect 285995 539547 286061 539548
rect 284208 507454 284528 507486
rect 284208 507218 284250 507454
rect 284486 507218 284528 507454
rect 284208 507134 284528 507218
rect 284208 506898 284250 507134
rect 284486 506898 284528 507134
rect 284208 506866 284528 506898
rect 284894 292637 284954 539547
rect 285294 466954 285914 498000
rect 285294 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 285914 466954
rect 285294 466634 285914 466718
rect 285294 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 285914 466634
rect 285294 430954 285914 466398
rect 285294 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 285914 430954
rect 285294 430634 285914 430718
rect 285294 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 285914 430634
rect 285294 394954 285914 430398
rect 285294 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 285914 394954
rect 285294 394634 285914 394718
rect 285294 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 285914 394634
rect 285294 358954 285914 394398
rect 285294 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 285914 358954
rect 285294 358634 285914 358718
rect 285294 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 285914 358634
rect 285294 322954 285914 358398
rect 285294 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 285914 322954
rect 285294 322634 285914 322718
rect 285294 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 285914 322634
rect 284891 292636 284957 292637
rect 284891 292572 284892 292636
rect 284956 292572 284957 292636
rect 284891 292571 284957 292572
rect 285294 286954 285914 322398
rect 285294 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 285914 286954
rect 285294 286634 285914 286718
rect 285294 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 285914 286634
rect 282131 280668 282197 280669
rect 282131 280604 282132 280668
rect 282196 280604 282197 280668
rect 282131 280603 282197 280604
rect 280794 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 281414 246454
rect 280794 246134 281414 246218
rect 280794 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 281414 246134
rect 280794 210454 281414 245898
rect 280794 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 281414 210454
rect 280794 210134 281414 210218
rect 280794 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 281414 210134
rect 280794 174454 281414 209898
rect 280794 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 281414 174454
rect 280794 174134 281414 174218
rect 280794 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 281414 174134
rect 280794 138454 281414 173898
rect 280794 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 281414 138454
rect 280794 138134 281414 138218
rect 280794 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 281414 138134
rect 280794 102454 281414 137898
rect 280794 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 281414 102454
rect 280794 102134 281414 102218
rect 280794 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 281414 102134
rect 280794 66454 281414 101898
rect 280794 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 281414 66454
rect 280794 66134 281414 66218
rect 280794 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 281414 66134
rect 280794 30454 281414 65898
rect 280794 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 281414 30454
rect 280794 30134 281414 30218
rect 280794 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 281414 30134
rect 280794 -6106 281414 29898
rect 280794 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 281414 -6106
rect 280794 -6426 281414 -6342
rect 280794 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 281414 -6426
rect 280794 -7654 281414 -6662
rect 285294 250954 285914 286398
rect 285998 281893 286058 539547
rect 285995 281892 286061 281893
rect 285995 281828 285996 281892
rect 286060 281828 286061 281892
rect 285995 281827 286061 281828
rect 287286 281077 287346 539683
rect 287651 539612 287717 539613
rect 287651 539548 287652 539612
rect 287716 539548 287717 539612
rect 287651 539547 287717 539548
rect 288387 539612 288453 539613
rect 288387 539548 288388 539612
rect 288452 539548 288453 539612
rect 288387 539547 288453 539548
rect 287283 281076 287349 281077
rect 287283 281012 287284 281076
rect 287348 281012 287349 281076
rect 287283 281011 287349 281012
rect 287654 280805 287714 539547
rect 288390 280941 288450 539547
rect 288574 281485 288634 539683
rect 289794 471454 290414 498000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 288571 281484 288637 281485
rect 288571 281420 288572 281484
rect 288636 281420 288637 281484
rect 288571 281419 288637 281420
rect 288387 280940 288453 280941
rect 288387 280876 288388 280940
rect 288452 280876 288453 280940
rect 288387 280875 288453 280876
rect 287651 280804 287717 280805
rect 287651 280740 287652 280804
rect 287716 280740 287717 280804
rect 287651 280739 287717 280740
rect 285294 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 285914 250954
rect 285294 250634 285914 250718
rect 285294 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 285914 250634
rect 285294 214954 285914 250398
rect 285294 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 285914 214954
rect 285294 214634 285914 214718
rect 285294 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 285914 214634
rect 285294 178954 285914 214398
rect 285294 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 285914 178954
rect 285294 178634 285914 178718
rect 285294 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 285914 178634
rect 285294 142954 285914 178398
rect 285294 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 285914 142954
rect 285294 142634 285914 142718
rect 285294 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 285914 142634
rect 285294 106954 285914 142398
rect 285294 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 285914 106954
rect 285294 106634 285914 106718
rect 285294 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 285914 106634
rect 285294 70954 285914 106398
rect 285294 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 285914 70954
rect 285294 70634 285914 70718
rect 285294 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 285914 70634
rect 285294 34954 285914 70398
rect 285294 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 285914 34954
rect 285294 34634 285914 34718
rect 285294 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 285914 34634
rect 285294 -7066 285914 34398
rect 285294 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 285914 -7066
rect 285294 -7386 285914 -7302
rect 285294 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 285914 -7386
rect 285294 -7654 285914 -7622
rect 289794 255454 290414 290898
rect 290598 281213 290658 539683
rect 290779 539612 290845 539613
rect 290779 539548 290780 539612
rect 290844 539548 290845 539612
rect 290779 539547 290845 539548
rect 291147 539612 291213 539613
rect 291147 539548 291148 539612
rect 291212 539548 291213 539612
rect 291147 539547 291213 539548
rect 292619 539612 292685 539613
rect 292619 539548 292620 539612
rect 292684 539548 292685 539612
rect 292619 539547 292685 539548
rect 293907 539612 293973 539613
rect 293907 539548 293908 539612
rect 293972 539548 293973 539612
rect 293907 539547 293973 539548
rect 295379 539612 295445 539613
rect 295379 539548 295380 539612
rect 295444 539548 295445 539612
rect 295379 539547 295445 539548
rect 290782 281349 290842 539547
rect 291150 282029 291210 539547
rect 291147 282028 291213 282029
rect 291147 281964 291148 282028
rect 291212 281964 291213 282028
rect 291147 281963 291213 281964
rect 290779 281348 290845 281349
rect 290779 281284 290780 281348
rect 290844 281284 290845 281348
rect 290779 281283 290845 281284
rect 290595 281212 290661 281213
rect 290595 281148 290596 281212
rect 290660 281148 290661 281212
rect 290595 281147 290661 281148
rect 292622 280533 292682 539547
rect 292619 280532 292685 280533
rect 292619 280468 292620 280532
rect 292684 280468 292685 280532
rect 292619 280467 292685 280468
rect 293910 279989 293970 539547
rect 294294 475954 294914 498000
rect 294294 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 294914 475954
rect 294294 475634 294914 475718
rect 294294 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 294914 475634
rect 294294 439954 294914 475398
rect 294294 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 294914 439954
rect 294294 439634 294914 439718
rect 294294 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 294914 439634
rect 294294 403954 294914 439398
rect 294294 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 294914 403954
rect 294294 403634 294914 403718
rect 294294 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 294914 403634
rect 294294 367954 294914 403398
rect 294294 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 294914 367954
rect 294294 367634 294914 367718
rect 294294 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 294914 367634
rect 294294 331954 294914 367398
rect 294294 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 294914 331954
rect 294294 331634 294914 331718
rect 294294 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 294914 331634
rect 294294 295954 294914 331398
rect 294294 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 294914 295954
rect 294294 295634 294914 295718
rect 294294 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 294914 295634
rect 293907 279988 293973 279989
rect 293907 279924 293908 279988
rect 293972 279924 293973 279988
rect 293907 279923 293973 279924
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 294294 259954 294914 295398
rect 295382 280125 295442 539547
rect 299568 511954 299888 511986
rect 299568 511718 299610 511954
rect 299846 511718 299888 511954
rect 299568 511634 299888 511718
rect 299568 511398 299610 511634
rect 299846 511398 299888 511634
rect 299568 511366 299888 511398
rect 314928 507454 315248 507486
rect 314928 507218 314970 507454
rect 315206 507218 315248 507454
rect 314928 507134 315248 507218
rect 314928 506898 314970 507134
rect 315206 506898 315248 507134
rect 314928 506866 315248 506898
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 298323 498812 298389 498813
rect 298323 498748 298324 498812
rect 298388 498748 298389 498812
rect 298323 498747 298389 498748
rect 297219 310044 297285 310045
rect 297219 309980 297220 310044
rect 297284 309980 297285 310044
rect 297219 309979 297285 309980
rect 295379 280124 295445 280125
rect 295379 280060 295380 280124
rect 295444 280060 295445 280124
rect 295379 280059 295445 280060
rect 297222 279445 297282 309979
rect 298326 282437 298386 498747
rect 298794 480454 299414 498000
rect 298794 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 299414 480454
rect 298794 480134 299414 480218
rect 298794 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 299414 480134
rect 298794 444454 299414 479898
rect 298794 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 299414 444454
rect 298794 444134 299414 444218
rect 298794 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 299414 444134
rect 298794 408454 299414 443898
rect 298794 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 299414 408454
rect 298794 408134 299414 408218
rect 298794 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 299414 408134
rect 298794 372454 299414 407898
rect 298794 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 299414 372454
rect 298794 372134 299414 372218
rect 298794 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 299414 372134
rect 298507 349756 298573 349757
rect 298507 349692 298508 349756
rect 298572 349692 298573 349756
rect 298507 349691 298573 349692
rect 298323 282436 298389 282437
rect 298323 282372 298324 282436
rect 298388 282372 298389 282436
rect 298323 282371 298389 282372
rect 297219 279444 297285 279445
rect 297219 279380 297220 279444
rect 297284 279380 297285 279444
rect 297219 279379 297285 279380
rect 294294 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 294914 259954
rect 294294 259634 294914 259718
rect 294294 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 294914 259634
rect 294294 223954 294914 259398
rect 294294 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 294914 223954
rect 294294 223634 294914 223718
rect 294294 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 294914 223634
rect 294294 187954 294914 223398
rect 294294 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 294914 187954
rect 294294 187634 294914 187718
rect 294294 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 294914 187634
rect 294294 151954 294914 187398
rect 294294 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 294914 151954
rect 294294 151634 294914 151718
rect 294294 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 294914 151634
rect 294294 115954 294914 151398
rect 294294 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 294914 115954
rect 294294 115634 294914 115718
rect 294294 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 294914 115634
rect 294294 79954 294914 115398
rect 294294 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 294914 79954
rect 294294 79634 294914 79718
rect 294294 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 294914 79634
rect 294294 43954 294914 79398
rect 294294 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 294914 43954
rect 294294 43634 294914 43718
rect 294294 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 294914 43634
rect 294294 7954 294914 43398
rect 294294 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 294914 7954
rect 294294 7634 294914 7718
rect 294294 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 294914 7634
rect 294294 -1306 294914 7398
rect 298510 3637 298570 349691
rect 298794 336454 299414 371898
rect 298794 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 299414 336454
rect 298794 336134 299414 336218
rect 298794 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 299414 336134
rect 303294 484954 303914 498000
rect 303294 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 303914 484954
rect 303294 484634 303914 484718
rect 303294 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 303914 484634
rect 303294 448954 303914 484398
rect 303294 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 303914 448954
rect 303294 448634 303914 448718
rect 303294 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 303914 448634
rect 303294 412954 303914 448398
rect 303294 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 303914 412954
rect 303294 412634 303914 412718
rect 303294 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 303914 412634
rect 303294 376954 303914 412398
rect 303294 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 303914 376954
rect 303294 376634 303914 376718
rect 303294 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 303914 376634
rect 303294 340954 303914 376398
rect 303294 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 303914 340954
rect 303294 340634 303914 340718
rect 303294 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 303914 340634
rect 299795 336020 299861 336021
rect 299795 335956 299796 336020
rect 299860 335956 299861 336020
rect 299795 335955 299861 335956
rect 298794 332000 299414 335898
rect 299611 331260 299677 331261
rect 299611 331196 299612 331260
rect 299676 331196 299677 331260
rect 299611 331195 299677 331196
rect 298794 264454 299414 278000
rect 298794 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 299414 264454
rect 298794 264134 299414 264218
rect 298794 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 299414 264134
rect 298794 228454 299414 263898
rect 298794 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 299414 228454
rect 298794 228134 299414 228218
rect 298794 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 299414 228134
rect 298794 222000 299414 227898
rect 299614 216749 299674 331195
rect 299611 216748 299677 216749
rect 299611 216684 299612 216748
rect 299676 216684 299677 216748
rect 299611 216683 299677 216684
rect 298794 48454 299414 58000
rect 298794 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 299414 48454
rect 298794 48134 299414 48218
rect 298794 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 299414 48134
rect 298794 12454 299414 47898
rect 298794 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 299414 12454
rect 298794 12134 299414 12218
rect 298794 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 299414 12134
rect 298507 3636 298573 3637
rect 298507 3572 298508 3636
rect 298572 3572 298573 3636
rect 298507 3571 298573 3572
rect 294294 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 294914 -1306
rect 294294 -1626 294914 -1542
rect 294294 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 294914 -1626
rect 294294 -7654 294914 -1862
rect 298794 -2266 299414 11898
rect 299798 3637 299858 335955
rect 303294 332000 303914 340398
rect 307794 489454 308414 498000
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 332000 308414 344898
rect 312294 493954 312914 498000
rect 312294 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 312914 493954
rect 312294 493634 312914 493718
rect 312294 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 312914 493634
rect 312294 457954 312914 493398
rect 312294 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 312914 457954
rect 312294 457634 312914 457718
rect 312294 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 312914 457634
rect 312294 421954 312914 457398
rect 312294 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 312914 421954
rect 312294 421634 312914 421718
rect 312294 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 312914 421634
rect 312294 385954 312914 421398
rect 312294 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 312914 385954
rect 312294 385634 312914 385718
rect 312294 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 312914 385634
rect 312294 349954 312914 385398
rect 312294 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 312914 349954
rect 312294 349634 312914 349718
rect 312294 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 312914 349634
rect 312294 332000 312914 349398
rect 316794 462454 317414 498000
rect 316794 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 317414 462454
rect 316794 462134 317414 462218
rect 316794 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 317414 462134
rect 316794 426454 317414 461898
rect 316794 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 317414 426454
rect 316794 426134 317414 426218
rect 316794 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 317414 426134
rect 316794 390454 317414 425898
rect 316794 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 317414 390454
rect 316794 390134 317414 390218
rect 316794 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 317414 390134
rect 316794 354454 317414 389898
rect 316794 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 317414 354454
rect 316794 354134 317414 354218
rect 316794 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 317414 354134
rect 316794 332000 317414 353898
rect 321294 466954 321914 498000
rect 321294 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 321914 466954
rect 321294 466634 321914 466718
rect 321294 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 321914 466634
rect 321294 430954 321914 466398
rect 321294 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 321914 430954
rect 321294 430634 321914 430718
rect 321294 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 321914 430634
rect 321294 394954 321914 430398
rect 321294 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 321914 394954
rect 321294 394634 321914 394718
rect 321294 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 321914 394634
rect 321294 358954 321914 394398
rect 321294 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 321914 358954
rect 321294 358634 321914 358718
rect 321294 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 321914 358634
rect 321294 332000 321914 358398
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 332000 326414 362898
rect 330294 705798 330914 711590
rect 330294 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 330914 705798
rect 330294 705478 330914 705562
rect 330294 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 330914 705478
rect 330294 691954 330914 705242
rect 330294 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 330914 691954
rect 330294 691634 330914 691718
rect 330294 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 330914 691634
rect 330294 655954 330914 691398
rect 330294 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 330914 655954
rect 330294 655634 330914 655718
rect 330294 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 330914 655634
rect 330294 619954 330914 655398
rect 330294 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 330914 619954
rect 330294 619634 330914 619718
rect 330294 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 330914 619634
rect 330294 583954 330914 619398
rect 330294 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 330914 583954
rect 330294 583634 330914 583718
rect 330294 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 330914 583634
rect 330294 547954 330914 583398
rect 330294 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 330914 547954
rect 330294 547634 330914 547718
rect 330294 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 330914 547634
rect 330294 511954 330914 547398
rect 330294 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 330914 511954
rect 330294 511634 330914 511718
rect 330294 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 330914 511634
rect 330294 475954 330914 511398
rect 330294 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 330914 475954
rect 330294 475634 330914 475718
rect 330294 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 330914 475634
rect 330294 439954 330914 475398
rect 330294 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 330914 439954
rect 330294 439634 330914 439718
rect 330294 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 330914 439634
rect 330294 403954 330914 439398
rect 330294 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 330914 403954
rect 330294 403634 330914 403718
rect 330294 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 330914 403634
rect 330294 367954 330914 403398
rect 330294 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 330914 367954
rect 330294 367634 330914 367718
rect 330294 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 330914 367634
rect 330294 332000 330914 367398
rect 334794 706758 335414 711590
rect 334794 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 335414 706758
rect 334794 706438 335414 706522
rect 334794 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 335414 706438
rect 334794 696454 335414 706202
rect 334794 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 335414 696454
rect 334794 696134 335414 696218
rect 334794 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 335414 696134
rect 334794 660454 335414 695898
rect 334794 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 335414 660454
rect 334794 660134 335414 660218
rect 334794 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 335414 660134
rect 334794 624454 335414 659898
rect 334794 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 335414 624454
rect 334794 624134 335414 624218
rect 334794 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 335414 624134
rect 334794 588454 335414 623898
rect 334794 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 335414 588454
rect 334794 588134 335414 588218
rect 334794 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 335414 588134
rect 334794 552454 335414 587898
rect 334794 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552218 335414 552454
rect 334794 552134 335414 552218
rect 334794 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 551898 335414 552134
rect 334794 516454 335414 551898
rect 334794 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 335414 516454
rect 334794 516134 335414 516218
rect 334794 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 335414 516134
rect 334794 480454 335414 515898
rect 334794 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 335414 480454
rect 334794 480134 335414 480218
rect 334794 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 335414 480134
rect 334794 444454 335414 479898
rect 334794 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 335414 444454
rect 334794 444134 335414 444218
rect 334794 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 335414 444134
rect 334794 408454 335414 443898
rect 334794 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 335414 408454
rect 334794 408134 335414 408218
rect 334794 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 335414 408134
rect 334794 372454 335414 407898
rect 334794 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 335414 372454
rect 334794 372134 335414 372218
rect 334794 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 335414 372134
rect 334794 336454 335414 371898
rect 334794 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 335414 336454
rect 334794 336134 335414 336218
rect 334794 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 335414 336134
rect 334794 332000 335414 335898
rect 339294 707718 339914 711590
rect 339294 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 339914 707718
rect 339294 707398 339914 707482
rect 339294 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 339914 707398
rect 339294 700954 339914 707162
rect 339294 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 339914 700954
rect 339294 700634 339914 700718
rect 339294 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 339914 700634
rect 339294 664954 339914 700398
rect 339294 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 339914 664954
rect 339294 664634 339914 664718
rect 339294 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 339914 664634
rect 339294 628954 339914 664398
rect 339294 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 339914 628954
rect 339294 628634 339914 628718
rect 339294 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 339914 628634
rect 339294 592954 339914 628398
rect 339294 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 339914 592954
rect 339294 592634 339914 592718
rect 339294 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 339914 592634
rect 339294 556954 339914 592398
rect 339294 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 339914 556954
rect 339294 556634 339914 556718
rect 339294 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 339914 556634
rect 339294 520954 339914 556398
rect 339294 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 339914 520954
rect 339294 520634 339914 520718
rect 339294 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 339914 520634
rect 339294 484954 339914 520398
rect 339294 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 339914 484954
rect 339294 484634 339914 484718
rect 339294 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 339914 484634
rect 339294 448954 339914 484398
rect 339294 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 339914 448954
rect 339294 448634 339914 448718
rect 339294 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 339914 448634
rect 339294 412954 339914 448398
rect 339294 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 339914 412954
rect 339294 412634 339914 412718
rect 339294 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 339914 412634
rect 339294 376954 339914 412398
rect 339294 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 339914 376954
rect 339294 376634 339914 376718
rect 339294 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 339914 376634
rect 339294 340954 339914 376398
rect 339294 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 339914 340954
rect 339294 340634 339914 340718
rect 339294 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 339914 340634
rect 339294 332000 339914 340398
rect 343794 708678 344414 711590
rect 343794 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 344414 708678
rect 343794 708358 344414 708442
rect 343794 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 344414 708358
rect 343794 669454 344414 708122
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 332000 344414 344898
rect 348294 709638 348914 711590
rect 348294 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 348914 709638
rect 348294 709318 348914 709402
rect 348294 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 348914 709318
rect 348294 673954 348914 709082
rect 348294 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 348914 673954
rect 348294 673634 348914 673718
rect 348294 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 348914 673634
rect 348294 637954 348914 673398
rect 352794 710598 353414 711590
rect 352794 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 353414 710598
rect 352794 710278 353414 710362
rect 352794 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 353414 710278
rect 352794 678454 353414 710042
rect 352794 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 353414 678454
rect 352794 678134 353414 678218
rect 352794 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 353414 678134
rect 352794 642454 353414 677898
rect 352794 642218 352826 642454
rect 353062 642218 353146 642454
rect 353382 642218 353414 642454
rect 352794 642134 353414 642218
rect 352794 641898 352826 642134
rect 353062 641898 353146 642134
rect 353382 641898 353414 642134
rect 357294 711558 357914 711590
rect 357294 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 357914 711558
rect 357294 711238 357914 711322
rect 357294 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 357914 711238
rect 357294 682954 357914 711002
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 360699 700364 360765 700365
rect 360699 700300 360700 700364
rect 360764 700300 360765 700364
rect 360699 700299 360765 700300
rect 357294 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 357914 682954
rect 357294 682634 357914 682718
rect 357294 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 357914 682634
rect 357294 646954 357914 682398
rect 359963 661332 360029 661333
rect 359963 661268 359964 661332
rect 360028 661268 360029 661332
rect 359963 661267 360029 661268
rect 357294 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 357914 646954
rect 357294 646634 357914 646718
rect 357294 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 357914 646634
rect 357294 642000 357914 646398
rect 358859 642020 358925 642021
rect 358859 641956 358860 642020
rect 358924 641956 358925 642020
rect 358859 641955 358925 641956
rect 351131 640660 351197 640661
rect 351131 640596 351132 640660
rect 351196 640596 351197 640660
rect 351131 640595 351197 640596
rect 348294 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 348914 637954
rect 348294 637634 348914 637718
rect 348294 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 348914 637634
rect 348294 601954 348914 637398
rect 348294 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 348914 601954
rect 348294 601634 348914 601718
rect 348294 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 348914 601634
rect 348294 565954 348914 601398
rect 348294 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 348914 565954
rect 348294 565634 348914 565718
rect 348294 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 348914 565634
rect 348294 529954 348914 565398
rect 348294 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 348914 529954
rect 348294 529634 348914 529718
rect 348294 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 348914 529634
rect 348294 493954 348914 529398
rect 349107 518940 349173 518941
rect 349107 518876 349108 518940
rect 349172 518876 349173 518940
rect 349107 518875 349173 518876
rect 348294 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 348914 493954
rect 348294 493634 348914 493718
rect 348294 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 348914 493634
rect 348294 457954 348914 493398
rect 348294 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 348914 457954
rect 348294 457634 348914 457718
rect 348294 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 348914 457634
rect 348294 421954 348914 457398
rect 348294 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 348914 421954
rect 348294 421634 348914 421718
rect 348294 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 348914 421634
rect 348294 385954 348914 421398
rect 348294 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 348914 385954
rect 348294 385634 348914 385718
rect 348294 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 348914 385634
rect 348294 349954 348914 385398
rect 348294 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 348914 349954
rect 348294 349634 348914 349718
rect 348294 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 348914 349634
rect 348294 332000 348914 349398
rect 304208 327239 304528 327376
rect 304208 327003 304250 327239
rect 304486 327003 304528 327239
rect 304208 326866 304528 327003
rect 334928 327239 335248 327376
rect 334928 327003 334970 327239
rect 335206 327003 335248 327239
rect 334928 326866 335248 327003
rect 319568 295954 319888 295986
rect 319568 295718 319610 295954
rect 319846 295718 319888 295954
rect 319568 295634 319888 295718
rect 319568 295398 319610 295634
rect 319846 295398 319888 295634
rect 319568 295366 319888 295398
rect 304208 291454 304528 291486
rect 304208 291218 304250 291454
rect 304486 291218 304528 291454
rect 304208 291134 304528 291218
rect 304208 290898 304250 291134
rect 304486 290898 304528 291134
rect 304208 290866 304528 290898
rect 334928 291454 335248 291486
rect 334928 291218 334970 291454
rect 335206 291218 335248 291454
rect 334928 291134 335248 291218
rect 334928 290898 334970 291134
rect 335206 290898 335248 291134
rect 334928 290866 335248 290898
rect 303294 268954 303914 278000
rect 303294 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 303914 268954
rect 303294 268634 303914 268718
rect 303294 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 303914 268634
rect 303294 232954 303914 268398
rect 303294 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 303914 232954
rect 303294 232634 303914 232718
rect 303294 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 303914 232634
rect 303294 222000 303914 232398
rect 307794 273454 308414 278000
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 222000 308414 236898
rect 312294 277954 312914 278000
rect 312294 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 312914 277954
rect 312294 277634 312914 277718
rect 312294 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 312914 277634
rect 312294 241954 312914 277398
rect 312294 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 312914 241954
rect 312294 241634 312914 241718
rect 312294 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 312914 241634
rect 312294 222000 312914 241398
rect 330294 259954 330914 278000
rect 330294 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 330914 259954
rect 330294 259634 330914 259718
rect 330294 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 330914 259634
rect 330294 223954 330914 259398
rect 330294 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 330914 223954
rect 330294 223634 330914 223718
rect 330294 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 330914 223634
rect 330294 222000 330914 223398
rect 334794 264454 335414 278000
rect 334794 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 335414 264454
rect 334794 264134 335414 264218
rect 334794 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 335414 264134
rect 334794 228454 335414 263898
rect 334794 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 335414 228454
rect 334794 228134 335414 228218
rect 334794 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 335414 228134
rect 334794 222000 335414 227898
rect 339294 268954 339914 278000
rect 339294 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 339914 268954
rect 339294 268634 339914 268718
rect 339294 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 339914 268634
rect 339294 232954 339914 268398
rect 339294 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 339914 232954
rect 339294 232634 339914 232718
rect 339294 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 339914 232634
rect 339294 222000 339914 232398
rect 343794 273454 344414 278000
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 222000 344414 236898
rect 348294 277954 348914 278000
rect 348294 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 348914 277954
rect 348294 277634 348914 277718
rect 348294 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 348914 277634
rect 348294 241954 348914 277398
rect 348294 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 348914 241954
rect 348294 241634 348914 241718
rect 348294 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 348914 241634
rect 348294 205954 348914 241398
rect 348294 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 348914 205954
rect 348294 205634 348914 205718
rect 348294 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 348914 205634
rect 319568 187954 319888 187986
rect 319568 187718 319610 187954
rect 319846 187718 319888 187954
rect 319568 187634 319888 187718
rect 319568 187398 319610 187634
rect 319846 187398 319888 187634
rect 319568 187366 319888 187398
rect 304208 183454 304528 183486
rect 304208 183218 304250 183454
rect 304486 183218 304528 183454
rect 304208 183134 304528 183218
rect 304208 182898 304250 183134
rect 304486 182898 304528 183134
rect 304208 182866 304528 182898
rect 334928 183454 335248 183486
rect 334928 183218 334970 183454
rect 335206 183218 335248 183454
rect 334928 183134 335248 183218
rect 334928 182898 334970 183134
rect 335206 182898 335248 183134
rect 334928 182866 335248 182898
rect 348294 169954 348914 205398
rect 348294 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 348914 169954
rect 348294 169634 348914 169718
rect 348294 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 348914 169634
rect 319568 151954 319888 151986
rect 319568 151718 319610 151954
rect 319846 151718 319888 151954
rect 319568 151634 319888 151718
rect 319568 151398 319610 151634
rect 319846 151398 319888 151634
rect 319568 151366 319888 151398
rect 304208 147454 304528 147486
rect 304208 147218 304250 147454
rect 304486 147218 304528 147454
rect 304208 147134 304528 147218
rect 304208 146898 304250 147134
rect 304486 146898 304528 147134
rect 304208 146866 304528 146898
rect 334928 147454 335248 147486
rect 334928 147218 334970 147454
rect 335206 147218 335248 147454
rect 334928 147134 335248 147218
rect 334928 146898 334970 147134
rect 335206 146898 335248 147134
rect 334928 146866 335248 146898
rect 348294 133954 348914 169398
rect 348294 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 348914 133954
rect 348294 133634 348914 133718
rect 348294 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 348914 133634
rect 319568 115954 319888 115986
rect 319568 115718 319610 115954
rect 319846 115718 319888 115954
rect 319568 115634 319888 115718
rect 319568 115398 319610 115634
rect 319846 115398 319888 115634
rect 319568 115366 319888 115398
rect 304208 111454 304528 111486
rect 304208 111218 304250 111454
rect 304486 111218 304528 111454
rect 304208 111134 304528 111218
rect 304208 110898 304250 111134
rect 304486 110898 304528 111134
rect 304208 110866 304528 110898
rect 334928 111454 335248 111486
rect 334928 111218 334970 111454
rect 335206 111218 335248 111454
rect 334928 111134 335248 111218
rect 334928 110898 334970 111134
rect 335206 110898 335248 111134
rect 334928 110866 335248 110898
rect 340827 108356 340893 108357
rect 340827 108292 340828 108356
rect 340892 108292 340893 108356
rect 340827 108291 340893 108292
rect 340091 85508 340157 85509
rect 340091 85444 340092 85508
rect 340156 85444 340157 85508
rect 340091 85443 340157 85444
rect 319568 79954 319888 79986
rect 319568 79718 319610 79954
rect 319846 79718 319888 79954
rect 319568 79634 319888 79718
rect 319568 79398 319610 79634
rect 319846 79398 319888 79634
rect 319568 79366 319888 79398
rect 304208 75454 304528 75486
rect 304208 75218 304250 75454
rect 304486 75218 304528 75454
rect 304208 75134 304528 75218
rect 304208 74898 304250 75134
rect 304486 74898 304528 75134
rect 304208 74866 304528 74898
rect 334928 75454 335248 75486
rect 334928 75218 334970 75454
rect 335206 75218 335248 75454
rect 334928 75134 335248 75218
rect 334928 74898 334970 75134
rect 335206 74898 335248 75134
rect 334928 74866 335248 74898
rect 303294 52954 303914 58000
rect 303294 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 303914 52954
rect 303294 52634 303914 52718
rect 303294 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 303914 52634
rect 303294 16954 303914 52398
rect 303294 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 303914 16954
rect 303294 16634 303914 16718
rect 303294 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 303914 16634
rect 299795 3636 299861 3637
rect 299795 3572 299796 3636
rect 299860 3572 299861 3636
rect 299795 3571 299861 3572
rect 298794 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 299414 -2266
rect 298794 -2586 299414 -2502
rect 298794 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 299414 -2586
rect 298794 -7654 299414 -2822
rect 303294 -3226 303914 16398
rect 303294 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 303914 -3226
rect 303294 -3546 303914 -3462
rect 303294 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 303914 -3546
rect 303294 -7654 303914 -3782
rect 307794 57454 308414 58000
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -4186 308414 20898
rect 307794 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 308414 -4186
rect 307794 -4506 308414 -4422
rect 307794 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 308414 -4506
rect 307794 -7654 308414 -4742
rect 312294 25954 312914 58000
rect 312294 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 312914 25954
rect 312294 25634 312914 25718
rect 312294 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 312914 25634
rect 312294 -5146 312914 25398
rect 312294 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 312914 -5146
rect 312294 -5466 312914 -5382
rect 312294 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 312914 -5466
rect 312294 -7654 312914 -5702
rect 316794 30454 317414 58000
rect 316794 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 317414 30454
rect 316794 30134 317414 30218
rect 316794 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 317414 30134
rect 316794 -6106 317414 29898
rect 316794 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 317414 -6106
rect 316794 -6426 317414 -6342
rect 316794 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 317414 -6426
rect 316794 -7654 317414 -6662
rect 321294 34954 321914 58000
rect 321294 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 321914 34954
rect 321294 34634 321914 34718
rect 321294 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 321914 34634
rect 321294 -7066 321914 34398
rect 321294 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 321914 -7066
rect 321294 -7386 321914 -7302
rect 321294 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 321914 -7386
rect 321294 -7654 321914 -7622
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 330294 43954 330914 58000
rect 330294 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 330914 43954
rect 330294 43634 330914 43718
rect 330294 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 330914 43634
rect 330294 7954 330914 43398
rect 330294 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 330914 7954
rect 330294 7634 330914 7718
rect 330294 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 330914 7634
rect 330294 -1306 330914 7398
rect 330294 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 330914 -1306
rect 330294 -1626 330914 -1542
rect 330294 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 330914 -1626
rect 330294 -7654 330914 -1862
rect 334794 48454 335414 58000
rect 334794 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 335414 48454
rect 334794 48134 335414 48218
rect 334794 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 335414 48134
rect 334794 12454 335414 47898
rect 334794 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 335414 12454
rect 334794 12134 335414 12218
rect 334794 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 335414 12134
rect 334794 -2266 335414 11898
rect 334794 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 335414 -2266
rect 334794 -2586 335414 -2502
rect 334794 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 335414 -2586
rect 334794 -7654 335414 -2822
rect 339294 52954 339914 58000
rect 339294 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 339914 52954
rect 339294 52634 339914 52718
rect 339294 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 339914 52634
rect 339294 16954 339914 52398
rect 339294 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 339914 16954
rect 339294 16634 339914 16718
rect 339294 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 339914 16634
rect 339294 -3226 339914 16398
rect 340094 3501 340154 85443
rect 340275 73540 340341 73541
rect 340275 73476 340276 73540
rect 340340 73476 340341 73540
rect 340275 73475 340341 73476
rect 340278 55861 340338 73475
rect 340275 55860 340341 55861
rect 340275 55796 340276 55860
rect 340340 55796 340341 55860
rect 340275 55795 340341 55796
rect 340830 39269 340890 108291
rect 342299 106180 342365 106181
rect 342299 106116 342300 106180
rect 342364 106116 342365 106180
rect 342299 106115 342365 106116
rect 341011 95300 341077 95301
rect 341011 95236 341012 95300
rect 341076 95236 341077 95300
rect 341011 95235 341077 95236
rect 341014 61573 341074 95235
rect 342302 85509 342362 106115
rect 348294 97954 348914 133398
rect 348294 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 348914 97954
rect 348294 97634 348914 97718
rect 348294 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 348914 97634
rect 342299 85508 342365 85509
rect 342299 85444 342300 85508
rect 342364 85444 342365 85508
rect 342299 85443 342365 85444
rect 342483 84420 342549 84421
rect 342483 84356 342484 84420
rect 342548 84356 342549 84420
rect 342483 84355 342549 84356
rect 342299 82244 342365 82245
rect 342299 82180 342300 82244
rect 342364 82180 342365 82244
rect 342299 82179 342365 82180
rect 341379 79388 341445 79389
rect 341379 79324 341380 79388
rect 341444 79324 341445 79388
rect 341379 79323 341445 79324
rect 341195 71364 341261 71365
rect 341195 71300 341196 71364
rect 341260 71300 341261 71364
rect 341195 71299 341261 71300
rect 341011 61572 341077 61573
rect 341011 61508 341012 61572
rect 341076 61508 341077 61572
rect 341011 61507 341077 61508
rect 341198 61437 341258 71299
rect 341195 61436 341261 61437
rect 341195 61372 341196 61436
rect 341260 61372 341261 61436
rect 341195 61371 341261 61372
rect 340827 39268 340893 39269
rect 340827 39204 340828 39268
rect 340892 39204 340893 39268
rect 340827 39203 340893 39204
rect 340091 3500 340157 3501
rect 340091 3436 340092 3500
rect 340156 3436 340157 3500
rect 340091 3435 340157 3436
rect 341382 3365 341442 79323
rect 342302 5133 342362 82179
rect 342486 57221 342546 84355
rect 342667 77892 342733 77893
rect 342667 77828 342668 77892
rect 342732 77828 342733 77892
rect 342667 77827 342733 77828
rect 342670 59941 342730 77827
rect 348294 61954 348914 97398
rect 348294 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 348914 61954
rect 348294 61634 348914 61718
rect 348294 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 348914 61634
rect 342667 59940 342733 59941
rect 342667 59876 342668 59940
rect 342732 59876 342733 59940
rect 342667 59875 342733 59876
rect 343794 57454 344414 58000
rect 342483 57220 342549 57221
rect 342483 57156 342484 57220
rect 342548 57156 342549 57220
rect 342483 57155 342549 57156
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 342299 5132 342365 5133
rect 342299 5068 342300 5132
rect 342364 5068 342365 5132
rect 342299 5067 342365 5068
rect 341379 3364 341445 3365
rect 341379 3300 341380 3364
rect 341444 3300 341445 3364
rect 341379 3299 341445 3300
rect 339294 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 339914 -3226
rect 339294 -3546 339914 -3462
rect 339294 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 339914 -3546
rect 339294 -7654 339914 -3782
rect 343794 -4186 344414 20898
rect 343794 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 344414 -4186
rect 343794 -4506 344414 -4422
rect 343794 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 344414 -4506
rect 343794 -7654 344414 -4742
rect 348294 25954 348914 61398
rect 348294 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 348914 25954
rect 348294 25634 348914 25718
rect 348294 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 348914 25634
rect 348294 -5146 348914 25398
rect 349110 3637 349170 518875
rect 349291 496908 349357 496909
rect 349291 496844 349292 496908
rect 349356 496844 349357 496908
rect 349291 496843 349357 496844
rect 349294 60077 349354 496843
rect 351134 218109 351194 640595
rect 352794 606454 353414 641898
rect 355179 640524 355245 640525
rect 355179 640460 355180 640524
rect 355244 640460 355245 640524
rect 355179 640459 355245 640460
rect 352794 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 353414 606454
rect 352794 606134 353414 606218
rect 352794 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 353414 606134
rect 352794 570454 353414 605898
rect 352794 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 353414 570454
rect 352794 570134 353414 570218
rect 352794 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 353414 570134
rect 352794 534454 353414 569898
rect 352794 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 353414 534454
rect 352794 534134 353414 534218
rect 352794 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 353414 534134
rect 352794 498454 353414 533898
rect 352794 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 353414 498454
rect 352794 498134 353414 498218
rect 352794 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 353414 498134
rect 352794 462454 353414 497898
rect 352794 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 353414 462454
rect 352794 462134 353414 462218
rect 352794 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 353414 462134
rect 352794 426454 353414 461898
rect 352794 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 353414 426454
rect 352794 426134 353414 426218
rect 352794 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 353414 426134
rect 352794 390454 353414 425898
rect 352794 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 353414 390454
rect 352794 390134 353414 390218
rect 352794 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 353414 390134
rect 352794 354454 353414 389898
rect 352794 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 353414 354454
rect 352794 354134 353414 354218
rect 352794 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 353414 354134
rect 352794 332000 353414 353898
rect 351867 320244 351933 320245
rect 351867 320180 351868 320244
rect 351932 320180 351933 320244
rect 351867 320179 351933 320180
rect 351870 225589 351930 320179
rect 352794 246454 353414 278000
rect 352794 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 353414 246454
rect 352794 246134 353414 246218
rect 352794 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 353414 246134
rect 351867 225588 351933 225589
rect 351867 225524 351868 225588
rect 351932 225524 351933 225588
rect 351867 225523 351933 225524
rect 351131 218108 351197 218109
rect 351131 218044 351132 218108
rect 351196 218044 351197 218108
rect 351131 218043 351197 218044
rect 352794 210454 353414 245898
rect 352794 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 353414 210454
rect 352794 210134 353414 210218
rect 352794 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 353414 210134
rect 352794 174454 353414 209898
rect 352794 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 353414 174454
rect 352794 174134 353414 174218
rect 352794 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 353414 174134
rect 352794 138454 353414 173898
rect 352794 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 353414 138454
rect 352794 138134 353414 138218
rect 352794 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 353414 138134
rect 352794 102454 353414 137898
rect 352794 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 353414 102454
rect 352794 102134 353414 102218
rect 352794 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 353414 102134
rect 352794 66454 353414 101898
rect 355182 99517 355242 640459
rect 358675 639708 358741 639709
rect 358675 639644 358676 639708
rect 358740 639644 358741 639708
rect 358675 639643 358741 639644
rect 355363 639436 355429 639437
rect 355363 639372 355364 639436
rect 355428 639372 355429 639436
rect 355363 639371 355429 639372
rect 355366 258093 355426 639371
rect 358307 559740 358373 559741
rect 358307 559676 358308 559740
rect 358372 559676 358373 559740
rect 358307 559675 358373 559676
rect 358123 555524 358189 555525
rect 358123 555460 358124 555524
rect 358188 555460 358189 555524
rect 358123 555459 358189 555460
rect 358126 547365 358186 555459
rect 358123 547364 358189 547365
rect 358123 547300 358124 547364
rect 358188 547300 358189 547364
rect 358123 547299 358189 547300
rect 358310 540701 358370 559675
rect 358491 554164 358557 554165
rect 358491 554100 358492 554164
rect 358556 554100 358557 554164
rect 358491 554099 358557 554100
rect 358307 540700 358373 540701
rect 358307 540636 358308 540700
rect 358372 540636 358373 540700
rect 358307 540635 358373 540636
rect 358494 516901 358554 554099
rect 358678 527781 358738 639643
rect 358675 527780 358741 527781
rect 358675 527716 358676 527780
rect 358740 527716 358741 527780
rect 358675 527715 358741 527716
rect 358491 516900 358557 516901
rect 358491 516836 358492 516900
rect 358556 516836 358557 516900
rect 358491 516835 358557 516836
rect 358862 502349 358922 641955
rect 359043 554028 359109 554029
rect 359043 553964 359044 554028
rect 359108 553964 359109 554028
rect 359043 553963 359109 553964
rect 359046 505069 359106 553963
rect 359966 552669 360026 661267
rect 359963 552668 360029 552669
rect 359963 552604 359964 552668
rect 360028 552604 360029 552668
rect 359963 552603 360029 552604
rect 359227 551988 359293 551989
rect 359227 551924 359228 551988
rect 359292 551924 359293 551988
rect 359227 551923 359293 551924
rect 359230 530637 359290 551923
rect 359411 551716 359477 551717
rect 359411 551652 359412 551716
rect 359476 551652 359477 551716
rect 359411 551651 359477 551652
rect 359414 542061 359474 551651
rect 359411 542060 359477 542061
rect 359411 541996 359412 542060
rect 359476 541996 359477 542060
rect 359411 541995 359477 541996
rect 359227 530636 359293 530637
rect 359227 530572 359228 530636
rect 359292 530572 359293 530636
rect 359227 530571 359293 530572
rect 359043 505068 359109 505069
rect 359043 505004 359044 505068
rect 359108 505004 359109 505068
rect 359043 505003 359109 505004
rect 358859 502348 358925 502349
rect 358859 502284 358860 502348
rect 358924 502284 358925 502348
rect 358859 502283 358925 502284
rect 360702 499357 360762 700299
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 642000 362414 650898
rect 366294 705798 366914 711590
rect 366294 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 366914 705798
rect 366294 705478 366914 705562
rect 366294 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 366914 705478
rect 366294 691954 366914 705242
rect 366294 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 366914 691954
rect 366294 691634 366914 691718
rect 366294 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 366914 691634
rect 366294 655954 366914 691398
rect 366294 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 366914 655954
rect 366294 655634 366914 655718
rect 366294 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 366914 655634
rect 366294 642000 366914 655398
rect 370794 706758 371414 711590
rect 370794 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 371414 706758
rect 370794 706438 371414 706522
rect 370794 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 371414 706438
rect 370794 696454 371414 706202
rect 370794 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 371414 696454
rect 370794 696134 371414 696218
rect 370794 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 371414 696134
rect 370794 660454 371414 695898
rect 370794 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 371414 660454
rect 370794 660134 371414 660218
rect 370794 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 371414 660134
rect 370794 642000 371414 659898
rect 375294 707718 375914 711590
rect 375294 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 375914 707718
rect 375294 707398 375914 707482
rect 375294 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 375914 707398
rect 375294 700954 375914 707162
rect 375294 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 375914 700954
rect 375294 700634 375914 700718
rect 375294 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 375914 700634
rect 375294 664954 375914 700398
rect 375294 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 375914 664954
rect 375294 664634 375914 664718
rect 375294 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 375914 664634
rect 375294 642000 375914 664398
rect 379794 708678 380414 711590
rect 379794 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 380414 708678
rect 379794 708358 380414 708442
rect 379794 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 380414 708358
rect 379794 669454 380414 708122
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 642000 380414 668898
rect 384294 709638 384914 711590
rect 384294 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 384914 709638
rect 384294 709318 384914 709402
rect 384294 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 384914 709318
rect 384294 673954 384914 709082
rect 384294 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 384914 673954
rect 384294 673634 384914 673718
rect 384294 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 384914 673634
rect 384294 642000 384914 673398
rect 388794 710598 389414 711590
rect 388794 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 389414 710598
rect 388794 710278 389414 710362
rect 388794 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 389414 710278
rect 388794 678454 389414 710042
rect 388794 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 389414 678454
rect 388794 678134 389414 678218
rect 388794 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 389414 678134
rect 388794 642361 389414 677898
rect 388794 642125 388826 642361
rect 389062 642125 389146 642361
rect 389382 642125 389414 642361
rect 388794 642000 389414 642125
rect 393294 711558 393914 711590
rect 393294 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 393914 711558
rect 393294 711238 393914 711322
rect 393294 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 393914 711238
rect 393294 682954 393914 711002
rect 393294 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 393914 682954
rect 393294 682634 393914 682718
rect 393294 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 393914 682634
rect 393294 646954 393914 682398
rect 393294 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 393914 646954
rect 393294 646634 393914 646718
rect 393294 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 393914 646634
rect 393294 642000 393914 646398
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 402294 705798 402914 711590
rect 402294 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 402914 705798
rect 402294 705478 402914 705562
rect 402294 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 402914 705478
rect 402294 691954 402914 705242
rect 402294 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 402914 691954
rect 402294 691634 402914 691718
rect 402294 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 402914 691634
rect 401547 662692 401613 662693
rect 401547 662628 401548 662692
rect 401612 662628 401613 662692
rect 401547 662627 401613 662628
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 642000 398414 650898
rect 398603 642156 398669 642157
rect 398603 642092 398604 642156
rect 398668 642092 398669 642156
rect 398603 642091 398669 642092
rect 363459 641748 363525 641749
rect 363459 641684 363460 641748
rect 363524 641684 363525 641748
rect 363459 641683 363525 641684
rect 362723 639572 362789 639573
rect 362723 639508 362724 639572
rect 362788 639508 362789 639572
rect 362723 639507 362789 639508
rect 362355 639436 362421 639437
rect 362355 639372 362356 639436
rect 362420 639372 362421 639436
rect 362355 639371 362421 639372
rect 362539 639436 362605 639437
rect 362539 639372 362540 639436
rect 362604 639372 362605 639436
rect 362539 639371 362605 639372
rect 362358 595509 362418 639371
rect 362355 595508 362421 595509
rect 362355 595444 362356 595508
rect 362420 595444 362421 595508
rect 362355 595443 362421 595444
rect 361619 571980 361685 571981
rect 361619 571916 361620 571980
rect 361684 571916 361685 571980
rect 361619 571915 361685 571916
rect 361435 558380 361501 558381
rect 361435 558316 361436 558380
rect 361500 558316 361501 558380
rect 361435 558315 361501 558316
rect 361438 499901 361498 558315
rect 361435 499900 361501 499901
rect 361435 499836 361436 499900
rect 361500 499836 361501 499900
rect 361435 499835 361501 499836
rect 361622 499765 361682 571915
rect 362542 565045 362602 639371
rect 362539 565044 362605 565045
rect 362539 564980 362540 565044
rect 362604 564980 362605 565044
rect 362539 564979 362605 564980
rect 362726 551581 362786 639507
rect 362907 593332 362973 593333
rect 362907 593268 362908 593332
rect 362972 593268 362973 593332
rect 362907 593267 362973 593268
rect 362723 551580 362789 551581
rect 362723 551516 362724 551580
rect 362788 551516 362789 551580
rect 362723 551515 362789 551516
rect 362910 499901 362970 593267
rect 363462 593197 363522 641683
rect 377259 639708 377325 639709
rect 377259 639644 377260 639708
rect 377324 639644 377325 639708
rect 377259 639643 377325 639644
rect 364011 639436 364077 639437
rect 364011 639372 364012 639436
rect 364076 639372 364077 639436
rect 364011 639371 364077 639372
rect 363459 593196 363525 593197
rect 363459 593132 363460 593196
rect 363524 593132 363525 593196
rect 363459 593131 363525 593132
rect 364014 581773 364074 639371
rect 377262 639165 377322 639643
rect 381123 639572 381189 639573
rect 381123 639508 381124 639572
rect 381188 639508 381189 639572
rect 381123 639507 381189 639508
rect 377259 639164 377325 639165
rect 377259 639100 377260 639164
rect 377324 639100 377325 639164
rect 377259 639099 377325 639100
rect 381126 639029 381186 639507
rect 381123 639028 381189 639029
rect 381123 638964 381124 639028
rect 381188 638964 381189 639028
rect 381123 638963 381189 638964
rect 379568 619954 379888 619986
rect 379568 619718 379610 619954
rect 379846 619718 379888 619954
rect 379568 619634 379888 619718
rect 379568 619398 379610 619634
rect 379846 619398 379888 619634
rect 379568 619366 379888 619398
rect 364208 615454 364528 615486
rect 364208 615218 364250 615454
rect 364486 615218 364528 615454
rect 364208 615134 364528 615218
rect 364208 614898 364250 615134
rect 364486 614898 364528 615134
rect 364208 614866 364528 614898
rect 394928 615454 395248 615486
rect 394928 615218 394970 615454
rect 395206 615218 395248 615454
rect 394928 615134 395248 615218
rect 394928 614898 394970 615134
rect 395206 614898 395248 615134
rect 394928 614866 395248 614898
rect 369899 599588 369965 599589
rect 369899 599524 369900 599588
rect 369964 599524 369965 599588
rect 369899 599523 369965 599524
rect 368979 597684 369045 597685
rect 368979 597620 368980 597684
rect 369044 597620 369045 597684
rect 368979 597619 369045 597620
rect 364011 581772 364077 581773
rect 364011 581708 364012 581772
rect 364076 581708 364077 581772
rect 364011 581707 364077 581708
rect 366219 568580 366285 568581
rect 366219 568516 366220 568580
rect 366284 568516 366285 568580
rect 366219 568515 366285 568516
rect 364747 563684 364813 563685
rect 364747 563620 364748 563684
rect 364812 563620 364813 563684
rect 364747 563619 364813 563620
rect 364208 543454 364528 543486
rect 364208 543218 364250 543454
rect 364486 543218 364528 543454
rect 364208 543134 364528 543218
rect 364208 542898 364250 543134
rect 364486 542898 364528 543134
rect 364208 542866 364528 542898
rect 364208 507454 364528 507486
rect 364208 507218 364250 507454
rect 364486 507218 364528 507454
rect 364208 507134 364528 507218
rect 364208 506898 364250 507134
rect 364486 506898 364528 507134
rect 364208 506866 364528 506898
rect 364750 499901 364810 563619
rect 362907 499900 362973 499901
rect 362907 499836 362908 499900
rect 362972 499836 362973 499900
rect 362907 499835 362973 499836
rect 364747 499900 364813 499901
rect 364747 499836 364748 499900
rect 364812 499836 364813 499900
rect 364747 499835 364813 499836
rect 361619 499764 361685 499765
rect 361619 499700 361620 499764
rect 361684 499700 361685 499764
rect 361619 499699 361685 499700
rect 366222 499493 366282 568515
rect 368243 563684 368309 563685
rect 368243 563620 368244 563684
rect 368308 563620 368309 563684
rect 368243 563619 368309 563620
rect 368246 499901 368306 563619
rect 368243 499900 368309 499901
rect 368243 499836 368244 499900
rect 368308 499836 368309 499900
rect 368243 499835 368309 499836
rect 368982 499493 369042 597619
rect 369902 499901 369962 599523
rect 382227 598228 382293 598229
rect 382227 598164 382228 598228
rect 382292 598164 382293 598228
rect 382227 598163 382293 598164
rect 370794 588454 371414 598000
rect 370794 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 371414 588454
rect 370794 588134 371414 588218
rect 370794 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 371414 588134
rect 370794 552361 371414 587898
rect 375294 592954 375914 598000
rect 375294 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 375914 592954
rect 375294 592634 375914 592718
rect 375294 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 375914 592634
rect 373211 581636 373277 581637
rect 373211 581572 373212 581636
rect 373276 581572 373277 581636
rect 373211 581571 373277 581572
rect 371555 563140 371621 563141
rect 371555 563076 371556 563140
rect 371620 563076 371621 563140
rect 371555 563075 371621 563076
rect 370794 552125 370826 552361
rect 371062 552125 371146 552361
rect 371382 552125 371414 552361
rect 370794 552000 371414 552125
rect 371558 499901 371618 563075
rect 369899 499900 369965 499901
rect 369899 499836 369900 499900
rect 369964 499836 369965 499900
rect 369899 499835 369965 499836
rect 371555 499900 371621 499901
rect 371555 499836 371556 499900
rect 371620 499836 371621 499900
rect 371555 499835 371621 499836
rect 366219 499492 366285 499493
rect 366219 499428 366220 499492
rect 366284 499428 366285 499492
rect 366219 499427 366285 499428
rect 368979 499492 369045 499493
rect 368979 499428 368980 499492
rect 369044 499428 369045 499492
rect 368979 499427 369045 499428
rect 360699 499356 360765 499357
rect 360699 499292 360700 499356
rect 360764 499292 360765 499356
rect 360699 499291 360765 499292
rect 373214 498133 373274 581571
rect 375294 556954 375914 592398
rect 379794 597454 380414 598000
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 376155 587212 376221 587213
rect 376155 587148 376156 587212
rect 376220 587148 376221 587212
rect 376155 587147 376221 587148
rect 375294 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 375914 556954
rect 375294 556634 375914 556718
rect 375294 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 375914 556634
rect 375294 552000 375914 556398
rect 376158 499901 376218 587147
rect 376891 578916 376957 578917
rect 376891 578852 376892 578916
rect 376956 578852 376957 578916
rect 376891 578851 376957 578852
rect 376339 561236 376405 561237
rect 376339 561172 376340 561236
rect 376404 561172 376405 561236
rect 376339 561171 376405 561172
rect 376155 499900 376221 499901
rect 376155 499836 376156 499900
rect 376220 499836 376221 499900
rect 376155 499835 376221 499836
rect 376342 499493 376402 561171
rect 376894 499901 376954 578851
rect 377259 569396 377325 569397
rect 377259 569332 377260 569396
rect 377324 569332 377325 569396
rect 377259 569331 377325 569332
rect 376891 499900 376957 499901
rect 376891 499836 376892 499900
rect 376956 499836 376957 499900
rect 376891 499835 376957 499836
rect 376339 499492 376405 499493
rect 376339 499428 376340 499492
rect 376404 499428 376405 499492
rect 376339 499427 376405 499428
rect 377262 498133 377322 569331
rect 378731 565860 378797 565861
rect 378731 565796 378732 565860
rect 378796 565796 378797 565860
rect 378731 565795 378797 565796
rect 373211 498132 373277 498133
rect 373211 498068 373212 498132
rect 373276 498068 373277 498132
rect 373211 498067 373277 498068
rect 377259 498132 377325 498133
rect 377259 498068 377260 498132
rect 377324 498068 377325 498132
rect 377259 498067 377325 498068
rect 357294 466954 357914 498000
rect 357294 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 357914 466954
rect 357294 466634 357914 466718
rect 357294 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 357914 466634
rect 357294 430954 357914 466398
rect 357294 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 357914 430954
rect 357294 430634 357914 430718
rect 357294 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 357914 430634
rect 357294 394954 357914 430398
rect 357294 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 357914 394954
rect 357294 394634 357914 394718
rect 357294 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 357914 394634
rect 357294 358954 357914 394398
rect 357294 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 357914 358954
rect 357294 358634 357914 358718
rect 357294 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 357914 358634
rect 357294 322954 357914 358398
rect 357294 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 357914 322954
rect 357294 322634 357914 322718
rect 357294 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 357914 322634
rect 357294 286954 357914 322398
rect 357294 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 357914 286954
rect 357294 286634 357914 286718
rect 357294 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 357914 286634
rect 355363 258092 355429 258093
rect 355363 258028 355364 258092
rect 355428 258028 355429 258092
rect 355363 258027 355429 258028
rect 357294 250954 357914 286398
rect 357294 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 357914 250954
rect 357294 250634 357914 250718
rect 357294 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 357914 250634
rect 357294 214954 357914 250398
rect 357294 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 357914 214954
rect 357294 214634 357914 214718
rect 357294 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 357914 214634
rect 357294 178954 357914 214398
rect 357294 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 357914 178954
rect 357294 178634 357914 178718
rect 357294 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 357914 178634
rect 357294 142954 357914 178398
rect 357294 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 357914 142954
rect 357294 142634 357914 142718
rect 357294 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 357914 142634
rect 357294 106954 357914 142398
rect 357294 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 357914 106954
rect 357294 106634 357914 106718
rect 357294 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 357914 106634
rect 355179 99516 355245 99517
rect 355179 99452 355180 99516
rect 355244 99452 355245 99516
rect 355179 99451 355245 99452
rect 352794 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 353414 66454
rect 352794 66134 353414 66218
rect 352794 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 353414 66134
rect 349291 60076 349357 60077
rect 349291 60012 349292 60076
rect 349356 60012 349357 60076
rect 349291 60011 349357 60012
rect 352794 30454 353414 65898
rect 352794 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 353414 30454
rect 352794 30134 353414 30218
rect 352794 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 353414 30134
rect 349107 3636 349173 3637
rect 349107 3572 349108 3636
rect 349172 3572 349173 3636
rect 349107 3571 349173 3572
rect 348294 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 348914 -5146
rect 348294 -5466 348914 -5382
rect 348294 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 348914 -5466
rect 348294 -7654 348914 -5702
rect 352794 -6106 353414 29898
rect 352794 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 353414 -6106
rect 352794 -6426 353414 -6342
rect 352794 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 353414 -6426
rect 352794 -7654 353414 -6662
rect 357294 70954 357914 106398
rect 357294 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 357914 70954
rect 357294 70634 357914 70718
rect 357294 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 357914 70634
rect 357294 34954 357914 70398
rect 357294 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 357914 34954
rect 357294 34634 357914 34718
rect 357294 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 357914 34634
rect 357294 -7066 357914 34398
rect 357294 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 357914 -7066
rect 357294 -7386 357914 -7302
rect 357294 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 357914 -7386
rect 357294 -7654 357914 -7622
rect 361794 471454 362414 498000
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 366294 475954 366914 498000
rect 366294 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 366914 475954
rect 366294 475634 366914 475718
rect 366294 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 366914 475634
rect 366294 439954 366914 475398
rect 366294 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 366914 439954
rect 366294 439634 366914 439718
rect 366294 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 366914 439634
rect 366294 403954 366914 439398
rect 366294 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 366914 403954
rect 366294 403634 366914 403718
rect 366294 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 366914 403634
rect 366294 367954 366914 403398
rect 366294 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 366914 367954
rect 366294 367634 366914 367718
rect 366294 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 366914 367634
rect 366294 331954 366914 367398
rect 366294 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 366914 331954
rect 366294 331634 366914 331718
rect 366294 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 366914 331634
rect 366294 295954 366914 331398
rect 366294 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 366914 295954
rect 366294 295634 366914 295718
rect 366294 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 366914 295634
rect 366294 259954 366914 295398
rect 366294 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 366914 259954
rect 366294 259634 366914 259718
rect 366294 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 366914 259634
rect 366294 223954 366914 259398
rect 366294 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 366914 223954
rect 366294 223634 366914 223718
rect 366294 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 366914 223634
rect 366294 187954 366914 223398
rect 366294 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 366914 187954
rect 366294 187634 366914 187718
rect 366294 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 366914 187634
rect 366294 151954 366914 187398
rect 366294 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 366914 151954
rect 366294 151634 366914 151718
rect 366294 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 366914 151634
rect 366294 115954 366914 151398
rect 366294 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 366914 115954
rect 366294 115634 366914 115718
rect 366294 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 366914 115634
rect 366294 79954 366914 115398
rect 366294 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 366914 79954
rect 366294 79634 366914 79718
rect 366294 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 366914 79634
rect 366294 43954 366914 79398
rect 366294 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 366914 43954
rect 366294 43634 366914 43718
rect 366294 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 366914 43634
rect 366294 7954 366914 43398
rect 366294 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 366914 7954
rect 366294 7634 366914 7718
rect 366294 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 366914 7634
rect 366294 -1306 366914 7398
rect 366294 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 366914 -1306
rect 366294 -1626 366914 -1542
rect 366294 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 366914 -1626
rect 366294 -7654 366914 -1862
rect 370794 480454 371414 498000
rect 370794 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 371414 480454
rect 370794 480134 371414 480218
rect 370794 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 371414 480134
rect 370794 444454 371414 479898
rect 370794 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 371414 444454
rect 370794 444134 371414 444218
rect 370794 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 371414 444134
rect 370794 408454 371414 443898
rect 370794 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 371414 408454
rect 370794 408134 371414 408218
rect 370794 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 371414 408134
rect 370794 372454 371414 407898
rect 370794 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 371414 372454
rect 370794 372134 371414 372218
rect 370794 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 371414 372134
rect 370794 336454 371414 371898
rect 370794 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 371414 336454
rect 370794 336134 371414 336218
rect 370794 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 371414 336134
rect 370794 300454 371414 335898
rect 370794 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 371414 300454
rect 370794 300134 371414 300218
rect 370794 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 371414 300134
rect 370794 264454 371414 299898
rect 370794 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 371414 264454
rect 370794 264134 371414 264218
rect 370794 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 371414 264134
rect 370794 228454 371414 263898
rect 370794 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 371414 228454
rect 370794 228134 371414 228218
rect 370794 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 371414 228134
rect 370794 192454 371414 227898
rect 370794 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 371414 192454
rect 370794 192134 371414 192218
rect 370794 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 371414 192134
rect 370794 156454 371414 191898
rect 370794 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 371414 156454
rect 370794 156134 371414 156218
rect 370794 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 371414 156134
rect 370794 120454 371414 155898
rect 370794 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 371414 120454
rect 370794 120134 371414 120218
rect 370794 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 371414 120134
rect 370794 84454 371414 119898
rect 370794 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 371414 84454
rect 370794 84134 371414 84218
rect 370794 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 371414 84134
rect 370794 48454 371414 83898
rect 370794 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 371414 48454
rect 370794 48134 371414 48218
rect 370794 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 371414 48134
rect 370794 12454 371414 47898
rect 370794 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 371414 12454
rect 370794 12134 371414 12218
rect 370794 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 371414 12134
rect 370794 -2266 371414 11898
rect 370794 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 371414 -2266
rect 370794 -2586 371414 -2502
rect 370794 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 371414 -2586
rect 370794 -7654 371414 -2822
rect 375294 484954 375914 498000
rect 378734 497997 378794 565795
rect 379794 561454 380414 596898
rect 380939 589932 381005 589933
rect 380939 589868 380940 589932
rect 381004 589868 381005 589932
rect 380939 589867 381005 589868
rect 380571 569260 380637 569261
rect 380571 569196 380572 569260
rect 380636 569196 380637 569260
rect 380571 569195 380637 569196
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 552000 380414 560898
rect 379568 511954 379888 511986
rect 379568 511718 379610 511954
rect 379846 511718 379888 511954
rect 379568 511634 379888 511718
rect 379568 511398 379610 511634
rect 379846 511398 379888 511634
rect 379568 511366 379888 511398
rect 380574 499901 380634 569195
rect 380942 499901 381002 589867
rect 380571 499900 380637 499901
rect 380571 499836 380572 499900
rect 380636 499836 380637 499900
rect 380571 499835 380637 499836
rect 380939 499900 381005 499901
rect 380939 499836 380940 499900
rect 381004 499836 381005 499900
rect 380939 499835 381005 499836
rect 378731 497996 378797 497997
rect 378731 497932 378732 497996
rect 378796 497932 378797 497996
rect 378731 497931 378797 497932
rect 375294 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 375914 484954
rect 375294 484634 375914 484718
rect 375294 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 375914 484634
rect 375294 448954 375914 484398
rect 375294 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 375914 448954
rect 375294 448634 375914 448718
rect 375294 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 375914 448634
rect 375294 412954 375914 448398
rect 375294 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 375914 412954
rect 375294 412634 375914 412718
rect 375294 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 375914 412634
rect 375294 376954 375914 412398
rect 375294 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 375914 376954
rect 375294 376634 375914 376718
rect 375294 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 375914 376634
rect 375294 340954 375914 376398
rect 375294 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 375914 340954
rect 375294 340634 375914 340718
rect 375294 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 375914 340634
rect 375294 304954 375914 340398
rect 375294 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 375914 304954
rect 375294 304634 375914 304718
rect 375294 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 375914 304634
rect 375294 268954 375914 304398
rect 375294 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 375914 268954
rect 375294 268634 375914 268718
rect 375294 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 375914 268634
rect 375294 232954 375914 268398
rect 375294 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 375914 232954
rect 375294 232634 375914 232718
rect 375294 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 375914 232634
rect 375294 196954 375914 232398
rect 375294 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 375914 196954
rect 375294 196634 375914 196718
rect 375294 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 375914 196634
rect 375294 160954 375914 196398
rect 375294 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 375914 160954
rect 375294 160634 375914 160718
rect 375294 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 375914 160634
rect 375294 124954 375914 160398
rect 375294 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 375914 124954
rect 375294 124634 375914 124718
rect 375294 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 375914 124634
rect 375294 88954 375914 124398
rect 375294 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 375914 88954
rect 375294 88634 375914 88718
rect 375294 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 375914 88634
rect 375294 52954 375914 88398
rect 375294 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 375914 52954
rect 375294 52634 375914 52718
rect 375294 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 375914 52634
rect 375294 16954 375914 52398
rect 375294 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 375914 16954
rect 375294 16634 375914 16718
rect 375294 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 375914 16634
rect 375294 -3226 375914 16398
rect 375294 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 375914 -3226
rect 375294 -3546 375914 -3462
rect 375294 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 375914 -3546
rect 375294 -7654 375914 -3782
rect 379794 489454 380414 498000
rect 382230 497453 382290 598163
rect 384067 582996 384133 582997
rect 384067 582932 384068 582996
rect 384132 582932 384133 582996
rect 384067 582931 384133 582932
rect 382779 563684 382845 563685
rect 382779 563620 382780 563684
rect 382844 563620 382845 563684
rect 382779 563619 382845 563620
rect 382782 499901 382842 563619
rect 382779 499900 382845 499901
rect 382779 499836 382780 499900
rect 382844 499836 382845 499900
rect 382779 499835 382845 499836
rect 384070 498133 384130 582931
rect 394739 580412 394805 580413
rect 394739 580348 394740 580412
rect 394804 580348 394805 580412
rect 394739 580347 394805 580348
rect 389587 580276 389653 580277
rect 389587 580212 389588 580276
rect 389652 580212 389653 580276
rect 389587 580211 389653 580212
rect 385539 579596 385605 579597
rect 385539 579532 385540 579596
rect 385604 579532 385605 579596
rect 385539 579531 385605 579532
rect 385542 499901 385602 579531
rect 385723 564500 385789 564501
rect 385723 564436 385724 564500
rect 385788 564436 385789 564500
rect 385723 564435 385789 564436
rect 385539 499900 385605 499901
rect 385539 499836 385540 499900
rect 385604 499836 385605 499900
rect 385539 499835 385605 499836
rect 385726 499765 385786 564435
rect 386459 562460 386525 562461
rect 386459 562396 386460 562460
rect 386524 562396 386525 562460
rect 386459 562395 386525 562396
rect 386462 499901 386522 562395
rect 389590 499901 389650 580211
rect 391979 577556 392045 577557
rect 391979 577492 391980 577556
rect 392044 577492 392045 577556
rect 391979 577491 392045 577492
rect 391059 573340 391125 573341
rect 391059 573276 391060 573340
rect 391124 573276 391125 573340
rect 391059 573275 391125 573276
rect 386459 499900 386525 499901
rect 386459 499836 386460 499900
rect 386524 499836 386525 499900
rect 386459 499835 386525 499836
rect 389587 499900 389653 499901
rect 389587 499836 389588 499900
rect 389652 499836 389653 499900
rect 389587 499835 389653 499836
rect 385723 499764 385789 499765
rect 385723 499700 385724 499764
rect 385788 499700 385789 499764
rect 385723 499699 385789 499700
rect 384067 498132 384133 498133
rect 384067 498068 384068 498132
rect 384132 498068 384133 498132
rect 384067 498067 384133 498068
rect 382227 497452 382293 497453
rect 382227 497388 382228 497452
rect 382292 497388 382293 497452
rect 382227 497387 382293 497388
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -4186 380414 20898
rect 379794 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 380414 -4186
rect 379794 -4506 380414 -4422
rect 379794 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 380414 -4506
rect 379794 -7654 380414 -4742
rect 384294 493954 384914 498000
rect 384294 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 384914 493954
rect 384294 493634 384914 493718
rect 384294 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 384914 493634
rect 384294 457954 384914 493398
rect 384294 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 384914 457954
rect 384294 457634 384914 457718
rect 384294 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 384914 457634
rect 384294 421954 384914 457398
rect 384294 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 384914 421954
rect 384294 421634 384914 421718
rect 384294 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 384914 421634
rect 384294 385954 384914 421398
rect 384294 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 384914 385954
rect 384294 385634 384914 385718
rect 384294 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 384914 385634
rect 384294 349954 384914 385398
rect 384294 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 384914 349954
rect 384294 349634 384914 349718
rect 384294 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 384914 349634
rect 384294 313954 384914 349398
rect 384294 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 384914 313954
rect 384294 313634 384914 313718
rect 384294 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 384914 313634
rect 384294 277954 384914 313398
rect 384294 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 384914 277954
rect 384294 277634 384914 277718
rect 384294 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 384914 277634
rect 384294 241954 384914 277398
rect 384294 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 384914 241954
rect 384294 241634 384914 241718
rect 384294 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 384914 241634
rect 384294 205954 384914 241398
rect 384294 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 384914 205954
rect 384294 205634 384914 205718
rect 384294 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 384914 205634
rect 384294 169954 384914 205398
rect 384294 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 384914 169954
rect 384294 169634 384914 169718
rect 384294 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 384914 169634
rect 384294 133954 384914 169398
rect 384294 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 384914 133954
rect 384294 133634 384914 133718
rect 384294 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 384914 133634
rect 384294 97954 384914 133398
rect 384294 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 384914 97954
rect 384294 97634 384914 97718
rect 384294 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 384914 97634
rect 384294 61954 384914 97398
rect 384294 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 384914 61954
rect 384294 61634 384914 61718
rect 384294 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 384914 61634
rect 384294 25954 384914 61398
rect 384294 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 384914 25954
rect 384294 25634 384914 25718
rect 384294 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 384914 25634
rect 384294 -5146 384914 25398
rect 384294 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 384914 -5146
rect 384294 -5466 384914 -5382
rect 384294 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 384914 -5466
rect 384294 -7654 384914 -5702
rect 388794 462454 389414 498000
rect 391062 497997 391122 573275
rect 391982 499901 392042 577491
rect 394003 575516 394069 575517
rect 394003 575452 394004 575516
rect 394068 575452 394069 575516
rect 394003 575451 394069 575452
rect 391979 499900 392045 499901
rect 391979 499836 391980 499900
rect 392044 499836 392045 499900
rect 391979 499835 392045 499836
rect 391059 497996 391125 497997
rect 391059 497932 391060 497996
rect 391124 497932 391125 497996
rect 391059 497931 391125 497932
rect 388794 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 389414 462454
rect 388794 462134 389414 462218
rect 388794 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 389414 462134
rect 388794 426454 389414 461898
rect 388794 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 389414 426454
rect 388794 426134 389414 426218
rect 388794 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 389414 426134
rect 388794 390454 389414 425898
rect 388794 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 389414 390454
rect 388794 390134 389414 390218
rect 388794 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 389414 390134
rect 388794 354454 389414 389898
rect 388794 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 389414 354454
rect 388794 354134 389414 354218
rect 388794 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 389414 354134
rect 388794 318454 389414 353898
rect 388794 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 389414 318454
rect 388794 318134 389414 318218
rect 388794 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 389414 318134
rect 388794 282454 389414 317898
rect 388794 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 389414 282454
rect 388794 282134 389414 282218
rect 388794 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 389414 282134
rect 388794 246454 389414 281898
rect 388794 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 389414 246454
rect 388794 246134 389414 246218
rect 388794 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 389414 246134
rect 388794 210454 389414 245898
rect 388794 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 389414 210454
rect 388794 210134 389414 210218
rect 388794 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 389414 210134
rect 388794 174454 389414 209898
rect 388794 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 389414 174454
rect 388794 174134 389414 174218
rect 388794 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 389414 174134
rect 388794 138454 389414 173898
rect 388794 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 389414 138454
rect 388794 138134 389414 138218
rect 388794 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 389414 138134
rect 388794 102454 389414 137898
rect 388794 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 389414 102454
rect 388794 102134 389414 102218
rect 388794 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 389414 102134
rect 388794 66454 389414 101898
rect 388794 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 389414 66454
rect 388794 66134 389414 66218
rect 388794 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 389414 66134
rect 388794 30454 389414 65898
rect 388794 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 389414 30454
rect 388794 30134 389414 30218
rect 388794 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 389414 30134
rect 388794 -6106 389414 29898
rect 388794 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 389414 -6106
rect 388794 -6426 389414 -6342
rect 388794 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 389414 -6426
rect 388794 -7654 389414 -6662
rect 393294 466954 393914 498000
rect 394006 497589 394066 575451
rect 394742 499901 394802 580347
rect 394928 543454 395248 543486
rect 394928 543218 394970 543454
rect 395206 543218 395248 543454
rect 394928 543134 395248 543218
rect 394928 542898 394970 543134
rect 395206 542898 395248 543134
rect 394928 542866 395248 542898
rect 394928 507454 395248 507486
rect 394928 507218 394970 507454
rect 395206 507218 395248 507454
rect 394928 507134 395248 507218
rect 394928 506898 394970 507134
rect 395206 506898 395248 507134
rect 394928 506866 395248 506898
rect 398606 499901 398666 642091
rect 400627 562324 400693 562325
rect 400627 562260 400628 562324
rect 400692 562260 400693 562324
rect 400627 562259 400693 562260
rect 400443 561100 400509 561101
rect 400443 561036 400444 561100
rect 400508 561036 400509 561100
rect 400443 561035 400509 561036
rect 399155 560964 399221 560965
rect 399155 560900 399156 560964
rect 399220 560900 399221 560964
rect 399155 560899 399221 560900
rect 398787 559604 398853 559605
rect 398787 559540 398788 559604
rect 398852 559540 398853 559604
rect 398787 559539 398853 559540
rect 398790 514450 398850 559539
rect 398971 551308 399037 551309
rect 398971 551244 398972 551308
rect 399036 551244 399037 551308
rect 398971 551243 399037 551244
rect 398974 514770 399034 551243
rect 399158 523970 399218 560899
rect 400259 556748 400325 556749
rect 400259 556684 400260 556748
rect 400324 556684 400325 556748
rect 400259 556683 400325 556684
rect 399339 555388 399405 555389
rect 399339 555324 399340 555388
rect 399404 555324 399405 555388
rect 399339 555323 399405 555324
rect 399342 527781 399402 555323
rect 399339 527780 399405 527781
rect 399339 527716 399340 527780
rect 399404 527716 399405 527780
rect 399339 527715 399405 527716
rect 399158 523910 399402 523970
rect 399342 518669 399402 523910
rect 399339 518668 399405 518669
rect 399339 518604 399340 518668
rect 399404 518604 399405 518668
rect 399339 518603 399405 518604
rect 398974 514710 399586 514770
rect 398790 514390 399402 514450
rect 399342 507789 399402 514390
rect 399339 507788 399405 507789
rect 399339 507724 399340 507788
rect 399404 507724 399405 507788
rect 399339 507723 399405 507724
rect 399526 506021 399586 514710
rect 399523 506020 399589 506021
rect 399523 505956 399524 506020
rect 399588 505956 399589 506020
rect 399523 505955 399589 505956
rect 400262 501465 400322 556683
rect 400446 523225 400506 561035
rect 400630 537845 400690 562259
rect 400811 551444 400877 551445
rect 400811 551380 400812 551444
rect 400876 551380 400877 551444
rect 400811 551379 400877 551380
rect 400627 537844 400693 537845
rect 400627 537780 400628 537844
rect 400692 537780 400693 537844
rect 400627 537779 400693 537780
rect 400814 531861 400874 551379
rect 401550 539613 401610 662627
rect 401731 661332 401797 661333
rect 401731 661268 401732 661332
rect 401796 661268 401797 661332
rect 401731 661267 401797 661268
rect 401734 549269 401794 661267
rect 402294 655954 402914 691398
rect 406794 706758 407414 711590
rect 406794 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 407414 706758
rect 406794 706438 407414 706522
rect 406794 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 407414 706438
rect 406794 696454 407414 706202
rect 406794 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 407414 696454
rect 406794 696134 407414 696218
rect 406794 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 407414 696134
rect 405043 663100 405109 663101
rect 405043 663036 405044 663100
rect 405108 663036 405109 663100
rect 405043 663035 405109 663036
rect 403019 662556 403085 662557
rect 403019 662492 403020 662556
rect 403084 662492 403085 662556
rect 403019 662491 403085 662492
rect 402294 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 402914 655954
rect 402294 655634 402914 655718
rect 402294 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 402914 655634
rect 402294 642000 402914 655398
rect 401915 550084 401981 550085
rect 401915 550020 401916 550084
rect 401980 550020 401981 550084
rect 401915 550019 401981 550020
rect 401731 549268 401797 549269
rect 401731 549204 401732 549268
rect 401796 549204 401797 549268
rect 401731 549203 401797 549204
rect 401918 543693 401978 550019
rect 401915 543692 401981 543693
rect 401915 543628 401916 543692
rect 401980 543628 401981 543692
rect 401915 543627 401981 543628
rect 401547 539612 401613 539613
rect 401547 539548 401548 539612
rect 401612 539548 401613 539612
rect 401547 539547 401613 539548
rect 400811 531860 400877 531861
rect 400811 531796 400812 531860
rect 400876 531796 400877 531860
rect 400811 531795 400877 531796
rect 400443 523224 400509 523225
rect 400443 523160 400444 523224
rect 400508 523160 400509 523224
rect 400443 523159 400509 523160
rect 403022 513365 403082 662491
rect 403571 552124 403637 552125
rect 403571 552060 403572 552124
rect 403636 552060 403637 552124
rect 403571 552059 403637 552060
rect 403019 513364 403085 513365
rect 403019 513300 403020 513364
rect 403084 513300 403085 513364
rect 403019 513299 403085 513300
rect 400259 501464 400325 501465
rect 400259 501400 400260 501464
rect 400324 501400 400325 501464
rect 400259 501399 400325 501400
rect 394739 499900 394805 499901
rect 394739 499836 394740 499900
rect 394804 499836 394805 499900
rect 394739 499835 394805 499836
rect 398603 499900 398669 499901
rect 398603 499836 398604 499900
rect 398668 499836 398669 499900
rect 398603 499835 398669 499836
rect 394003 497588 394069 497589
rect 394003 497524 394004 497588
rect 394068 497524 394069 497588
rect 394003 497523 394069 497524
rect 393294 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 393914 466954
rect 393294 466634 393914 466718
rect 393294 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 393914 466634
rect 393294 430954 393914 466398
rect 393294 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 393914 430954
rect 393294 430634 393914 430718
rect 393294 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 393914 430634
rect 393294 394954 393914 430398
rect 393294 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 393914 394954
rect 393294 394634 393914 394718
rect 393294 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 393914 394634
rect 393294 358954 393914 394398
rect 393294 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 393914 358954
rect 393294 358634 393914 358718
rect 393294 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 393914 358634
rect 393294 322954 393914 358398
rect 393294 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 393914 322954
rect 393294 322634 393914 322718
rect 393294 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 393914 322634
rect 393294 286954 393914 322398
rect 393294 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 393914 286954
rect 393294 286634 393914 286718
rect 393294 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 393914 286634
rect 393294 250954 393914 286398
rect 393294 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 393914 250954
rect 393294 250634 393914 250718
rect 393294 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 393914 250634
rect 393294 214954 393914 250398
rect 393294 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 393914 214954
rect 393294 214634 393914 214718
rect 393294 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 393914 214634
rect 393294 178954 393914 214398
rect 393294 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 393914 178954
rect 393294 178634 393914 178718
rect 393294 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 393914 178634
rect 393294 142954 393914 178398
rect 393294 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 393914 142954
rect 393294 142634 393914 142718
rect 393294 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 393914 142634
rect 393294 106954 393914 142398
rect 393294 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 393914 106954
rect 393294 106634 393914 106718
rect 393294 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 393914 106634
rect 393294 70954 393914 106398
rect 393294 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 393914 70954
rect 393294 70634 393914 70718
rect 393294 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 393914 70634
rect 393294 34954 393914 70398
rect 393294 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 393914 34954
rect 393294 34634 393914 34718
rect 393294 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 393914 34634
rect 393294 -7066 393914 34398
rect 393294 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 393914 -7066
rect 393294 -7386 393914 -7302
rect 393294 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 393914 -7386
rect 393294 -7654 393914 -7622
rect 397794 471454 398414 498000
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 402294 475954 402914 498000
rect 402294 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 402914 475954
rect 402294 475634 402914 475718
rect 402294 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 402914 475634
rect 402294 439954 402914 475398
rect 402294 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 402914 439954
rect 402294 439634 402914 439718
rect 402294 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 402914 439634
rect 402294 403954 402914 439398
rect 402294 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 402914 403954
rect 402294 403634 402914 403718
rect 402294 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 402914 403634
rect 402294 367954 402914 403398
rect 402294 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 402914 367954
rect 402294 367634 402914 367718
rect 402294 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 402914 367634
rect 402294 331954 402914 367398
rect 402294 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 402914 331954
rect 402294 331634 402914 331718
rect 402294 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 402914 331634
rect 402294 295954 402914 331398
rect 402294 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 402914 295954
rect 402294 295634 402914 295718
rect 402294 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 402914 295634
rect 402294 259954 402914 295398
rect 402294 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 402914 259954
rect 402294 259634 402914 259718
rect 402294 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 402914 259634
rect 402294 223954 402914 259398
rect 402294 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 402914 223954
rect 402294 223634 402914 223718
rect 402294 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 402914 223634
rect 402294 187954 402914 223398
rect 402294 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 402914 187954
rect 402294 187634 402914 187718
rect 402294 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 402914 187634
rect 402294 151954 402914 187398
rect 402294 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 402914 151954
rect 402294 151634 402914 151718
rect 402294 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 402914 151634
rect 402294 115954 402914 151398
rect 402294 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 402914 115954
rect 402294 115634 402914 115718
rect 402294 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 402914 115634
rect 402294 79954 402914 115398
rect 402294 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 402914 79954
rect 402294 79634 402914 79718
rect 402294 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 402914 79634
rect 402294 43954 402914 79398
rect 403574 44845 403634 552059
rect 404859 538252 404925 538253
rect 404859 538188 404860 538252
rect 404924 538188 404925 538252
rect 404859 538187 404925 538188
rect 403571 44844 403637 44845
rect 403571 44780 403572 44844
rect 403636 44780 403637 44844
rect 403571 44779 403637 44780
rect 402294 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 402914 43954
rect 402294 43634 402914 43718
rect 402294 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 402914 43634
rect 402294 7954 402914 43398
rect 404862 24173 404922 538187
rect 405046 531589 405106 663035
rect 406794 660454 407414 695898
rect 406794 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 407414 660454
rect 406794 660134 407414 660218
rect 406794 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 407414 660134
rect 406794 624454 407414 659898
rect 406794 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 407414 624454
rect 406794 624134 407414 624218
rect 406794 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 407414 624134
rect 406794 588454 407414 623898
rect 406794 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 407414 588454
rect 406794 588134 407414 588218
rect 406794 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 407414 588134
rect 406794 552454 407414 587898
rect 406794 552218 406826 552454
rect 407062 552218 407146 552454
rect 407382 552218 407414 552454
rect 406794 552134 407414 552218
rect 406794 551898 406826 552134
rect 407062 551898 407146 552134
rect 407382 551898 407414 552134
rect 405043 531588 405109 531589
rect 405043 531524 405044 531588
rect 405108 531524 405109 531588
rect 405043 531523 405109 531524
rect 406794 516454 407414 551898
rect 406794 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 407414 516454
rect 406794 516134 407414 516218
rect 406794 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 407414 516134
rect 406794 480454 407414 515898
rect 406794 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 407414 480454
rect 406794 480134 407414 480218
rect 406794 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 407414 480134
rect 406794 444454 407414 479898
rect 406794 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 407414 444454
rect 406794 444134 407414 444218
rect 406794 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 407414 444134
rect 406794 408454 407414 443898
rect 406794 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 407414 408454
rect 406794 408134 407414 408218
rect 406794 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 407414 408134
rect 406794 372454 407414 407898
rect 406794 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 407414 372454
rect 406794 372134 407414 372218
rect 406794 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 407414 372134
rect 406794 336454 407414 371898
rect 406794 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 407414 336454
rect 406794 336134 407414 336218
rect 406794 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 407414 336134
rect 406794 300454 407414 335898
rect 406794 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 407414 300454
rect 406794 300134 407414 300218
rect 406794 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 407414 300134
rect 406794 264454 407414 299898
rect 406794 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 407414 264454
rect 406794 264134 407414 264218
rect 406794 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 407414 264134
rect 406794 228454 407414 263898
rect 406794 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 407414 228454
rect 406794 228134 407414 228218
rect 406794 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 407414 228134
rect 406794 192454 407414 227898
rect 406794 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 407414 192454
rect 406794 192134 407414 192218
rect 406794 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 407414 192134
rect 406794 156454 407414 191898
rect 406794 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 407414 156454
rect 406794 156134 407414 156218
rect 406794 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 407414 156134
rect 406794 120454 407414 155898
rect 406794 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 407414 120454
rect 406794 120134 407414 120218
rect 406794 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 407414 120134
rect 406794 84454 407414 119898
rect 406794 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 407414 84454
rect 406794 84134 407414 84218
rect 406794 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 407414 84134
rect 406794 48454 407414 83898
rect 406794 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 407414 48454
rect 406794 48134 407414 48218
rect 406794 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 407414 48134
rect 404859 24172 404925 24173
rect 404859 24108 404860 24172
rect 404924 24108 404925 24172
rect 404859 24107 404925 24108
rect 402294 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 402914 7954
rect 402294 7634 402914 7718
rect 402294 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 402914 7634
rect 402294 -1306 402914 7398
rect 402294 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 402914 -1306
rect 402294 -1626 402914 -1542
rect 402294 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 402914 -1626
rect 402294 -7654 402914 -1862
rect 406794 12454 407414 47898
rect 406794 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 407414 12454
rect 406794 12134 407414 12218
rect 406794 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 407414 12134
rect 406794 -2266 407414 11898
rect 406794 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 407414 -2266
rect 406794 -2586 407414 -2502
rect 406794 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 407414 -2586
rect 406794 -7654 407414 -2822
rect 411294 707718 411914 711590
rect 411294 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 411914 707718
rect 411294 707398 411914 707482
rect 411294 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 411914 707398
rect 411294 700954 411914 707162
rect 411294 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 411914 700954
rect 411294 700634 411914 700718
rect 411294 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 411914 700634
rect 411294 664954 411914 700398
rect 411294 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 411914 664954
rect 411294 664634 411914 664718
rect 411294 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 411914 664634
rect 411294 628954 411914 664398
rect 411294 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 411914 628954
rect 411294 628634 411914 628718
rect 411294 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 411914 628634
rect 411294 592954 411914 628398
rect 411294 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 411914 592954
rect 411294 592634 411914 592718
rect 411294 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 411914 592634
rect 411294 556954 411914 592398
rect 411294 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 411914 556954
rect 411294 556634 411914 556718
rect 411294 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 411914 556634
rect 411294 520954 411914 556398
rect 411294 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 411914 520954
rect 411294 520634 411914 520718
rect 411294 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 411914 520634
rect 411294 484954 411914 520398
rect 411294 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 411914 484954
rect 411294 484634 411914 484718
rect 411294 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 411914 484634
rect 411294 448954 411914 484398
rect 411294 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 411914 448954
rect 411294 448634 411914 448718
rect 411294 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 411914 448634
rect 411294 412954 411914 448398
rect 411294 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 411914 412954
rect 411294 412634 411914 412718
rect 411294 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 411914 412634
rect 411294 376954 411914 412398
rect 411294 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 411914 376954
rect 411294 376634 411914 376718
rect 411294 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 411914 376634
rect 411294 340954 411914 376398
rect 411294 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 411914 340954
rect 411294 340634 411914 340718
rect 411294 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 411914 340634
rect 411294 304954 411914 340398
rect 411294 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 411914 304954
rect 411294 304634 411914 304718
rect 411294 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 411914 304634
rect 411294 268954 411914 304398
rect 411294 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 411914 268954
rect 411294 268634 411914 268718
rect 411294 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 411914 268634
rect 411294 232954 411914 268398
rect 411294 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 411914 232954
rect 411294 232634 411914 232718
rect 411294 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 411914 232634
rect 411294 196954 411914 232398
rect 411294 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 411914 196954
rect 411294 196634 411914 196718
rect 411294 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 411914 196634
rect 411294 160954 411914 196398
rect 411294 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 411914 160954
rect 411294 160634 411914 160718
rect 411294 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 411914 160634
rect 411294 124954 411914 160398
rect 411294 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 411914 124954
rect 411294 124634 411914 124718
rect 411294 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 411914 124634
rect 411294 88954 411914 124398
rect 411294 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 411914 88954
rect 411294 88634 411914 88718
rect 411294 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 411914 88634
rect 411294 52954 411914 88398
rect 411294 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 411914 52954
rect 411294 52634 411914 52718
rect 411294 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 411914 52634
rect 411294 16954 411914 52398
rect 411294 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 411914 16954
rect 411294 16634 411914 16718
rect 411294 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 411914 16634
rect 411294 -3226 411914 16398
rect 411294 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 411914 -3226
rect 411294 -3546 411914 -3462
rect 411294 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 411914 -3546
rect 411294 -7654 411914 -3782
rect 415794 708678 416414 711590
rect 415794 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 416414 708678
rect 415794 708358 416414 708442
rect 415794 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 416414 708358
rect 415794 669454 416414 708122
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -4186 416414 20898
rect 415794 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 416414 -4186
rect 415794 -4506 416414 -4422
rect 415794 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 416414 -4506
rect 415794 -7654 416414 -4742
rect 420294 709638 420914 711590
rect 420294 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 420914 709638
rect 420294 709318 420914 709402
rect 420294 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 420914 709318
rect 420294 673954 420914 709082
rect 420294 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 420914 673954
rect 420294 673634 420914 673718
rect 420294 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 420914 673634
rect 420294 637954 420914 673398
rect 420294 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 420914 637954
rect 420294 637634 420914 637718
rect 420294 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 420914 637634
rect 420294 601954 420914 637398
rect 420294 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 420914 601954
rect 420294 601634 420914 601718
rect 420294 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 420914 601634
rect 420294 565954 420914 601398
rect 420294 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 420914 565954
rect 420294 565634 420914 565718
rect 420294 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 420914 565634
rect 420294 529954 420914 565398
rect 420294 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 420914 529954
rect 420294 529634 420914 529718
rect 420294 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 420914 529634
rect 420294 493954 420914 529398
rect 420294 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 420914 493954
rect 420294 493634 420914 493718
rect 420294 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 420914 493634
rect 420294 457954 420914 493398
rect 420294 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 420914 457954
rect 420294 457634 420914 457718
rect 420294 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 420914 457634
rect 420294 421954 420914 457398
rect 420294 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 420914 421954
rect 420294 421634 420914 421718
rect 420294 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 420914 421634
rect 420294 385954 420914 421398
rect 420294 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 420914 385954
rect 420294 385634 420914 385718
rect 420294 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 420914 385634
rect 420294 349954 420914 385398
rect 420294 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 420914 349954
rect 420294 349634 420914 349718
rect 420294 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 420914 349634
rect 420294 313954 420914 349398
rect 420294 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 420914 313954
rect 420294 313634 420914 313718
rect 420294 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 420914 313634
rect 420294 277954 420914 313398
rect 420294 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 420914 277954
rect 420294 277634 420914 277718
rect 420294 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 420914 277634
rect 420294 241954 420914 277398
rect 420294 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 420914 241954
rect 420294 241634 420914 241718
rect 420294 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 420914 241634
rect 420294 205954 420914 241398
rect 420294 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 420914 205954
rect 420294 205634 420914 205718
rect 420294 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 420914 205634
rect 420294 169954 420914 205398
rect 420294 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 420914 169954
rect 420294 169634 420914 169718
rect 420294 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 420914 169634
rect 420294 133954 420914 169398
rect 420294 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 420914 133954
rect 420294 133634 420914 133718
rect 420294 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 420914 133634
rect 420294 97954 420914 133398
rect 420294 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 420914 97954
rect 420294 97634 420914 97718
rect 420294 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 420914 97634
rect 420294 61954 420914 97398
rect 420294 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 420914 61954
rect 420294 61634 420914 61718
rect 420294 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 420914 61634
rect 420294 25954 420914 61398
rect 420294 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 420914 25954
rect 420294 25634 420914 25718
rect 420294 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 420914 25634
rect 420294 -5146 420914 25398
rect 420294 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 420914 -5146
rect 420294 -5466 420914 -5382
rect 420294 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 420914 -5466
rect 420294 -7654 420914 -5702
rect 424794 710598 425414 711590
rect 424794 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 425414 710598
rect 424794 710278 425414 710362
rect 424794 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 425414 710278
rect 424794 678454 425414 710042
rect 424794 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 425414 678454
rect 424794 678134 425414 678218
rect 424794 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 425414 678134
rect 424794 642454 425414 677898
rect 424794 642218 424826 642454
rect 425062 642218 425146 642454
rect 425382 642218 425414 642454
rect 424794 642134 425414 642218
rect 424794 641898 424826 642134
rect 425062 641898 425146 642134
rect 425382 641898 425414 642134
rect 424794 606454 425414 641898
rect 424794 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 425414 606454
rect 424794 606134 425414 606218
rect 424794 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 425414 606134
rect 424794 570454 425414 605898
rect 424794 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 425414 570454
rect 424794 570134 425414 570218
rect 424794 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 425414 570134
rect 424794 534454 425414 569898
rect 424794 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 425414 534454
rect 424794 534134 425414 534218
rect 424794 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 425414 534134
rect 424794 498454 425414 533898
rect 424794 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 425414 498454
rect 424794 498134 425414 498218
rect 424794 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 425414 498134
rect 424794 462454 425414 497898
rect 424794 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 425414 462454
rect 424794 462134 425414 462218
rect 424794 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 425414 462134
rect 424794 426454 425414 461898
rect 424794 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 425414 426454
rect 424794 426134 425414 426218
rect 424794 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 425414 426134
rect 424794 390454 425414 425898
rect 424794 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 425414 390454
rect 424794 390134 425414 390218
rect 424794 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 425414 390134
rect 424794 354454 425414 389898
rect 424794 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 425414 354454
rect 424794 354134 425414 354218
rect 424794 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 425414 354134
rect 424794 318454 425414 353898
rect 424794 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 425414 318454
rect 424794 318134 425414 318218
rect 424794 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 425414 318134
rect 424794 282454 425414 317898
rect 424794 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 425414 282454
rect 424794 282134 425414 282218
rect 424794 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 425414 282134
rect 424794 246454 425414 281898
rect 424794 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 425414 246454
rect 424794 246134 425414 246218
rect 424794 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 425414 246134
rect 424794 210454 425414 245898
rect 424794 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 425414 210454
rect 424794 210134 425414 210218
rect 424794 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 425414 210134
rect 424794 174454 425414 209898
rect 424794 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 425414 174454
rect 424794 174134 425414 174218
rect 424794 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 425414 174134
rect 424794 138454 425414 173898
rect 424794 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 425414 138454
rect 424794 138134 425414 138218
rect 424794 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 425414 138134
rect 424794 102454 425414 137898
rect 424794 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 425414 102454
rect 424794 102134 425414 102218
rect 424794 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 425414 102134
rect 424794 66454 425414 101898
rect 424794 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 425414 66454
rect 424794 66134 425414 66218
rect 424794 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 425414 66134
rect 424794 30454 425414 65898
rect 424794 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 425414 30454
rect 424794 30134 425414 30218
rect 424794 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 425414 30134
rect 424794 -6106 425414 29898
rect 424794 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 425414 -6106
rect 424794 -6426 425414 -6342
rect 424794 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 425414 -6426
rect 424794 -7654 425414 -6662
rect 429294 711558 429914 711590
rect 429294 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 429914 711558
rect 429294 711238 429914 711322
rect 429294 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 429914 711238
rect 429294 682954 429914 711002
rect 429294 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 429914 682954
rect 429294 682634 429914 682718
rect 429294 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 429914 682634
rect 429294 646954 429914 682398
rect 429294 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 429914 646954
rect 429294 646634 429914 646718
rect 429294 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 429914 646634
rect 429294 610954 429914 646398
rect 429294 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 429914 610954
rect 429294 610634 429914 610718
rect 429294 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 429914 610634
rect 429294 574954 429914 610398
rect 429294 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 429914 574954
rect 429294 574634 429914 574718
rect 429294 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 429914 574634
rect 429294 538954 429914 574398
rect 429294 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 429914 538954
rect 429294 538634 429914 538718
rect 429294 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 429914 538634
rect 429294 502954 429914 538398
rect 429294 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 429914 502954
rect 429294 502634 429914 502718
rect 429294 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 429914 502634
rect 429294 466954 429914 502398
rect 429294 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 429914 466954
rect 429294 466634 429914 466718
rect 429294 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 429914 466634
rect 429294 430954 429914 466398
rect 429294 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 429914 430954
rect 429294 430634 429914 430718
rect 429294 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 429914 430634
rect 429294 394954 429914 430398
rect 429294 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 429914 394954
rect 429294 394634 429914 394718
rect 429294 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 429914 394634
rect 429294 358954 429914 394398
rect 429294 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 429914 358954
rect 429294 358634 429914 358718
rect 429294 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 429914 358634
rect 429294 322954 429914 358398
rect 429294 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 429914 322954
rect 429294 322634 429914 322718
rect 429294 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 429914 322634
rect 429294 286954 429914 322398
rect 429294 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 429914 286954
rect 429294 286634 429914 286718
rect 429294 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 429914 286634
rect 429294 250954 429914 286398
rect 429294 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 429914 250954
rect 429294 250634 429914 250718
rect 429294 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 429914 250634
rect 429294 214954 429914 250398
rect 429294 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 429914 214954
rect 429294 214634 429914 214718
rect 429294 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 429914 214634
rect 429294 178954 429914 214398
rect 429294 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 429914 178954
rect 429294 178634 429914 178718
rect 429294 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 429914 178634
rect 429294 142954 429914 178398
rect 429294 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 429914 142954
rect 429294 142634 429914 142718
rect 429294 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 429914 142634
rect 429294 106954 429914 142398
rect 429294 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 429914 106954
rect 429294 106634 429914 106718
rect 429294 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 429914 106634
rect 429294 70954 429914 106398
rect 429294 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 429914 70954
rect 429294 70634 429914 70718
rect 429294 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 429914 70634
rect 429294 34954 429914 70398
rect 429294 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 429914 34954
rect 429294 34634 429914 34718
rect 429294 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 429914 34634
rect 429294 -7066 429914 34398
rect 429294 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 429914 -7066
rect 429294 -7386 429914 -7302
rect 429294 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 429914 -7386
rect 429294 -7654 429914 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 438294 705798 438914 711590
rect 438294 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 438914 705798
rect 438294 705478 438914 705562
rect 438294 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 438914 705478
rect 438294 691954 438914 705242
rect 438294 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 438914 691954
rect 438294 691634 438914 691718
rect 438294 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 438914 691634
rect 438294 655954 438914 691398
rect 438294 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 438914 655954
rect 438294 655634 438914 655718
rect 438294 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 438914 655634
rect 438294 619954 438914 655398
rect 438294 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 438914 619954
rect 438294 619634 438914 619718
rect 438294 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 438914 619634
rect 438294 583954 438914 619398
rect 438294 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 438914 583954
rect 438294 583634 438914 583718
rect 438294 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 438914 583634
rect 438294 547954 438914 583398
rect 438294 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 438914 547954
rect 438294 547634 438914 547718
rect 438294 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 438914 547634
rect 438294 511954 438914 547398
rect 438294 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 438914 511954
rect 438294 511634 438914 511718
rect 438294 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 438914 511634
rect 438294 475954 438914 511398
rect 438294 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 438914 475954
rect 438294 475634 438914 475718
rect 438294 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 438914 475634
rect 438294 439954 438914 475398
rect 438294 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 438914 439954
rect 438294 439634 438914 439718
rect 438294 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 438914 439634
rect 438294 403954 438914 439398
rect 438294 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 438914 403954
rect 438294 403634 438914 403718
rect 438294 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 438914 403634
rect 438294 367954 438914 403398
rect 438294 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 438914 367954
rect 438294 367634 438914 367718
rect 438294 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 438914 367634
rect 438294 331954 438914 367398
rect 438294 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 438914 331954
rect 438294 331634 438914 331718
rect 438294 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 438914 331634
rect 438294 295954 438914 331398
rect 438294 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 438914 295954
rect 438294 295634 438914 295718
rect 438294 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 438914 295634
rect 438294 259954 438914 295398
rect 438294 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 438914 259954
rect 438294 259634 438914 259718
rect 438294 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 438914 259634
rect 438294 223954 438914 259398
rect 438294 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 438914 223954
rect 438294 223634 438914 223718
rect 438294 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 438914 223634
rect 438294 187954 438914 223398
rect 438294 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 438914 187954
rect 438294 187634 438914 187718
rect 438294 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 438914 187634
rect 438294 151954 438914 187398
rect 438294 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 438914 151954
rect 438294 151634 438914 151718
rect 438294 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 438914 151634
rect 438294 115954 438914 151398
rect 438294 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 438914 115954
rect 438294 115634 438914 115718
rect 438294 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 438914 115634
rect 438294 79954 438914 115398
rect 438294 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 438914 79954
rect 438294 79634 438914 79718
rect 438294 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 438914 79634
rect 438294 43954 438914 79398
rect 438294 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 438914 43954
rect 438294 43634 438914 43718
rect 438294 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 438914 43634
rect 438294 7954 438914 43398
rect 438294 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 438914 7954
rect 438294 7634 438914 7718
rect 438294 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 438914 7634
rect 438294 -1306 438914 7398
rect 438294 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 438914 -1306
rect 438294 -1626 438914 -1542
rect 438294 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 438914 -1626
rect 438294 -7654 438914 -1862
rect 442794 706758 443414 711590
rect 442794 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 443414 706758
rect 442794 706438 443414 706522
rect 442794 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 443414 706438
rect 442794 696454 443414 706202
rect 442794 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 443414 696454
rect 442794 696134 443414 696218
rect 442794 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 443414 696134
rect 442794 660454 443414 695898
rect 442794 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 443414 660454
rect 442794 660134 443414 660218
rect 442794 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 443414 660134
rect 442794 624454 443414 659898
rect 442794 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 443414 624454
rect 442794 624134 443414 624218
rect 442794 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 443414 624134
rect 442794 588454 443414 623898
rect 442794 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 443414 588454
rect 442794 588134 443414 588218
rect 442794 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 443414 588134
rect 442794 552454 443414 587898
rect 442794 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 443414 552454
rect 442794 552134 443414 552218
rect 442794 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 443414 552134
rect 442794 516454 443414 551898
rect 442794 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 443414 516454
rect 442794 516134 443414 516218
rect 442794 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 443414 516134
rect 442794 480454 443414 515898
rect 442794 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 443414 480454
rect 442794 480134 443414 480218
rect 442794 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 443414 480134
rect 442794 444454 443414 479898
rect 442794 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 443414 444454
rect 442794 444134 443414 444218
rect 442794 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 443414 444134
rect 442794 408454 443414 443898
rect 442794 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 443414 408454
rect 442794 408134 443414 408218
rect 442794 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 443414 408134
rect 442794 372454 443414 407898
rect 442794 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 443414 372454
rect 442794 372134 443414 372218
rect 442794 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 443414 372134
rect 442794 336454 443414 371898
rect 442794 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 443414 336454
rect 442794 336134 443414 336218
rect 442794 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 443414 336134
rect 442794 300454 443414 335898
rect 442794 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 443414 300454
rect 442794 300134 443414 300218
rect 442794 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 443414 300134
rect 442794 264454 443414 299898
rect 442794 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 443414 264454
rect 442794 264134 443414 264218
rect 442794 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 443414 264134
rect 442794 228454 443414 263898
rect 442794 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 443414 228454
rect 442794 228134 443414 228218
rect 442794 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 443414 228134
rect 442794 192454 443414 227898
rect 442794 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 443414 192454
rect 442794 192134 443414 192218
rect 442794 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 443414 192134
rect 442794 156454 443414 191898
rect 442794 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 443414 156454
rect 442794 156134 443414 156218
rect 442794 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 443414 156134
rect 442794 120454 443414 155898
rect 442794 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 443414 120454
rect 442794 120134 443414 120218
rect 442794 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 443414 120134
rect 442794 84454 443414 119898
rect 442794 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 443414 84454
rect 442794 84134 443414 84218
rect 442794 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 443414 84134
rect 442794 48454 443414 83898
rect 442794 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 443414 48454
rect 442794 48134 443414 48218
rect 442794 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 443414 48134
rect 442794 12454 443414 47898
rect 442794 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 443414 12454
rect 442794 12134 443414 12218
rect 442794 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 443414 12134
rect 442794 -2266 443414 11898
rect 442794 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 443414 -2266
rect 442794 -2586 443414 -2502
rect 442794 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 443414 -2586
rect 442794 -7654 443414 -2822
rect 447294 707718 447914 711590
rect 447294 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 447914 707718
rect 447294 707398 447914 707482
rect 447294 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 447914 707398
rect 447294 700954 447914 707162
rect 447294 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 447914 700954
rect 447294 700634 447914 700718
rect 447294 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 447914 700634
rect 447294 664954 447914 700398
rect 447294 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 447914 664954
rect 447294 664634 447914 664718
rect 447294 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 447914 664634
rect 447294 628954 447914 664398
rect 447294 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 447914 628954
rect 447294 628634 447914 628718
rect 447294 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 447914 628634
rect 447294 592954 447914 628398
rect 447294 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 447914 592954
rect 447294 592634 447914 592718
rect 447294 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 447914 592634
rect 447294 556954 447914 592398
rect 447294 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 447914 556954
rect 447294 556634 447914 556718
rect 447294 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 447914 556634
rect 447294 520954 447914 556398
rect 447294 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 447914 520954
rect 447294 520634 447914 520718
rect 447294 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 447914 520634
rect 447294 484954 447914 520398
rect 447294 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 447914 484954
rect 447294 484634 447914 484718
rect 447294 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 447914 484634
rect 447294 448954 447914 484398
rect 447294 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 447914 448954
rect 447294 448634 447914 448718
rect 447294 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 447914 448634
rect 447294 412954 447914 448398
rect 447294 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 447914 412954
rect 447294 412634 447914 412718
rect 447294 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 447914 412634
rect 447294 376954 447914 412398
rect 447294 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 447914 376954
rect 447294 376634 447914 376718
rect 447294 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 447914 376634
rect 447294 340954 447914 376398
rect 447294 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 447914 340954
rect 447294 340634 447914 340718
rect 447294 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 447914 340634
rect 447294 304954 447914 340398
rect 447294 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 447914 304954
rect 447294 304634 447914 304718
rect 447294 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 447914 304634
rect 447294 268954 447914 304398
rect 447294 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 447914 268954
rect 447294 268634 447914 268718
rect 447294 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 447914 268634
rect 447294 232954 447914 268398
rect 447294 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 447914 232954
rect 447294 232634 447914 232718
rect 447294 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 447914 232634
rect 447294 196954 447914 232398
rect 447294 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 447914 196954
rect 447294 196634 447914 196718
rect 447294 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 447914 196634
rect 447294 160954 447914 196398
rect 447294 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 447914 160954
rect 447294 160634 447914 160718
rect 447294 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 447914 160634
rect 447294 124954 447914 160398
rect 447294 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 447914 124954
rect 447294 124634 447914 124718
rect 447294 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 447914 124634
rect 447294 88954 447914 124398
rect 447294 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 447914 88954
rect 447294 88634 447914 88718
rect 447294 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 447914 88634
rect 447294 52954 447914 88398
rect 447294 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 447914 52954
rect 447294 52634 447914 52718
rect 447294 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 447914 52634
rect 447294 16954 447914 52398
rect 447294 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 447914 16954
rect 447294 16634 447914 16718
rect 447294 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 447914 16634
rect 447294 -3226 447914 16398
rect 447294 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 447914 -3226
rect 447294 -3546 447914 -3462
rect 447294 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 447914 -3546
rect 447294 -7654 447914 -3782
rect 451794 708678 452414 711590
rect 451794 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 452414 708678
rect 451794 708358 452414 708442
rect 451794 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 452414 708358
rect 451794 669454 452414 708122
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -4186 452414 20898
rect 451794 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 452414 -4186
rect 451794 -4506 452414 -4422
rect 451794 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 452414 -4506
rect 451794 -7654 452414 -4742
rect 456294 709638 456914 711590
rect 456294 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 456914 709638
rect 456294 709318 456914 709402
rect 456294 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 456914 709318
rect 456294 673954 456914 709082
rect 456294 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 456914 673954
rect 456294 673634 456914 673718
rect 456294 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 456914 673634
rect 456294 637954 456914 673398
rect 456294 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 456914 637954
rect 456294 637634 456914 637718
rect 456294 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 456914 637634
rect 456294 601954 456914 637398
rect 456294 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 456914 601954
rect 456294 601634 456914 601718
rect 456294 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 456914 601634
rect 456294 565954 456914 601398
rect 456294 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 456914 565954
rect 456294 565634 456914 565718
rect 456294 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 456914 565634
rect 456294 529954 456914 565398
rect 456294 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 456914 529954
rect 456294 529634 456914 529718
rect 456294 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 456914 529634
rect 456294 493954 456914 529398
rect 456294 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 456914 493954
rect 456294 493634 456914 493718
rect 456294 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 456914 493634
rect 456294 457954 456914 493398
rect 456294 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 456914 457954
rect 456294 457634 456914 457718
rect 456294 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 456914 457634
rect 456294 421954 456914 457398
rect 456294 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 456914 421954
rect 456294 421634 456914 421718
rect 456294 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 456914 421634
rect 456294 385954 456914 421398
rect 456294 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 456914 385954
rect 456294 385634 456914 385718
rect 456294 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 456914 385634
rect 456294 349954 456914 385398
rect 456294 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 456914 349954
rect 456294 349634 456914 349718
rect 456294 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 456914 349634
rect 456294 313954 456914 349398
rect 456294 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 456914 313954
rect 456294 313634 456914 313718
rect 456294 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 456914 313634
rect 456294 277954 456914 313398
rect 456294 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 456914 277954
rect 456294 277634 456914 277718
rect 456294 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 456914 277634
rect 456294 241954 456914 277398
rect 456294 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 456914 241954
rect 456294 241634 456914 241718
rect 456294 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 456914 241634
rect 456294 205954 456914 241398
rect 456294 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 456914 205954
rect 456294 205634 456914 205718
rect 456294 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 456914 205634
rect 456294 169954 456914 205398
rect 456294 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 456914 169954
rect 456294 169634 456914 169718
rect 456294 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 456914 169634
rect 456294 133954 456914 169398
rect 456294 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 456914 133954
rect 456294 133634 456914 133718
rect 456294 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 456914 133634
rect 456294 97954 456914 133398
rect 456294 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 456914 97954
rect 456294 97634 456914 97718
rect 456294 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 456914 97634
rect 456294 61954 456914 97398
rect 456294 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 456914 61954
rect 456294 61634 456914 61718
rect 456294 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 456914 61634
rect 456294 25954 456914 61398
rect 456294 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 456914 25954
rect 456294 25634 456914 25718
rect 456294 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 456914 25634
rect 456294 -5146 456914 25398
rect 456294 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 456914 -5146
rect 456294 -5466 456914 -5382
rect 456294 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 456914 -5466
rect 456294 -7654 456914 -5702
rect 460794 710598 461414 711590
rect 460794 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 461414 710598
rect 460794 710278 461414 710362
rect 460794 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 461414 710278
rect 460794 678454 461414 710042
rect 460794 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 461414 678454
rect 460794 678134 461414 678218
rect 460794 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 461414 678134
rect 460794 642454 461414 677898
rect 460794 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642218 461414 642454
rect 460794 642134 461414 642218
rect 460794 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 641898 461414 642134
rect 460794 606454 461414 641898
rect 460794 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 461414 606454
rect 460794 606134 461414 606218
rect 460794 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 461414 606134
rect 460794 570454 461414 605898
rect 460794 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 461414 570454
rect 460794 570134 461414 570218
rect 460794 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 461414 570134
rect 460794 534454 461414 569898
rect 460794 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 461414 534454
rect 460794 534134 461414 534218
rect 460794 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 461414 534134
rect 460794 498454 461414 533898
rect 460794 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 461414 498454
rect 460794 498134 461414 498218
rect 460794 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 461414 498134
rect 460794 462454 461414 497898
rect 460794 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 461414 462454
rect 460794 462134 461414 462218
rect 460794 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 461414 462134
rect 460794 426454 461414 461898
rect 460794 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 461414 426454
rect 460794 426134 461414 426218
rect 460794 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 461414 426134
rect 460794 390454 461414 425898
rect 460794 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 461414 390454
rect 460794 390134 461414 390218
rect 460794 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 461414 390134
rect 460794 354454 461414 389898
rect 460794 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 461414 354454
rect 460794 354134 461414 354218
rect 460794 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 461414 354134
rect 460794 318454 461414 353898
rect 460794 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 461414 318454
rect 460794 318134 461414 318218
rect 460794 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 461414 318134
rect 460794 282454 461414 317898
rect 460794 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 461414 282454
rect 460794 282134 461414 282218
rect 460794 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 461414 282134
rect 460794 246454 461414 281898
rect 460794 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 461414 246454
rect 460794 246134 461414 246218
rect 460794 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 461414 246134
rect 460794 210454 461414 245898
rect 460794 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 461414 210454
rect 460794 210134 461414 210218
rect 460794 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 461414 210134
rect 460794 174454 461414 209898
rect 460794 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 461414 174454
rect 460794 174134 461414 174218
rect 460794 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 461414 174134
rect 460794 138454 461414 173898
rect 460794 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 461414 138454
rect 460794 138134 461414 138218
rect 460794 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 461414 138134
rect 460794 102454 461414 137898
rect 460794 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 461414 102454
rect 460794 102134 461414 102218
rect 460794 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 461414 102134
rect 460794 66454 461414 101898
rect 460794 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 461414 66454
rect 460794 66134 461414 66218
rect 460794 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 461414 66134
rect 460794 30454 461414 65898
rect 460794 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 461414 30454
rect 460794 30134 461414 30218
rect 460794 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 461414 30134
rect 460794 -6106 461414 29898
rect 460794 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 461414 -6106
rect 460794 -6426 461414 -6342
rect 460794 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 461414 -6426
rect 460794 -7654 461414 -6662
rect 465294 711558 465914 711590
rect 465294 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 465914 711558
rect 465294 711238 465914 711322
rect 465294 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 465914 711238
rect 465294 682954 465914 711002
rect 465294 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 465914 682954
rect 465294 682634 465914 682718
rect 465294 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 465914 682634
rect 465294 646954 465914 682398
rect 465294 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 465914 646954
rect 465294 646634 465914 646718
rect 465294 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 465914 646634
rect 465294 610954 465914 646398
rect 465294 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 465914 610954
rect 465294 610634 465914 610718
rect 465294 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 465914 610634
rect 465294 574954 465914 610398
rect 465294 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 465914 574954
rect 465294 574634 465914 574718
rect 465294 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 465914 574634
rect 465294 538954 465914 574398
rect 465294 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 465914 538954
rect 465294 538634 465914 538718
rect 465294 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 465914 538634
rect 465294 502954 465914 538398
rect 465294 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 465914 502954
rect 465294 502634 465914 502718
rect 465294 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 465914 502634
rect 465294 466954 465914 502398
rect 465294 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 465914 466954
rect 465294 466634 465914 466718
rect 465294 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 465914 466634
rect 465294 430954 465914 466398
rect 465294 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 465914 430954
rect 465294 430634 465914 430718
rect 465294 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 465914 430634
rect 465294 394954 465914 430398
rect 465294 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 465914 394954
rect 465294 394634 465914 394718
rect 465294 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 465914 394634
rect 465294 358954 465914 394398
rect 465294 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 465914 358954
rect 465294 358634 465914 358718
rect 465294 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 465914 358634
rect 465294 322954 465914 358398
rect 465294 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 465914 322954
rect 465294 322634 465914 322718
rect 465294 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 465914 322634
rect 465294 286954 465914 322398
rect 465294 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 465914 286954
rect 465294 286634 465914 286718
rect 465294 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 465914 286634
rect 465294 250954 465914 286398
rect 465294 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 465914 250954
rect 465294 250634 465914 250718
rect 465294 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 465914 250634
rect 465294 214954 465914 250398
rect 465294 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 465914 214954
rect 465294 214634 465914 214718
rect 465294 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 465914 214634
rect 465294 178954 465914 214398
rect 465294 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 465914 178954
rect 465294 178634 465914 178718
rect 465294 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 465914 178634
rect 465294 142954 465914 178398
rect 465294 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 465914 142954
rect 465294 142634 465914 142718
rect 465294 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 465914 142634
rect 465294 106954 465914 142398
rect 465294 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 465914 106954
rect 465294 106634 465914 106718
rect 465294 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 465914 106634
rect 465294 70954 465914 106398
rect 465294 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 465914 70954
rect 465294 70634 465914 70718
rect 465294 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 465914 70634
rect 465294 34954 465914 70398
rect 465294 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 465914 34954
rect 465294 34634 465914 34718
rect 465294 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 465914 34634
rect 465294 -7066 465914 34398
rect 465294 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 465914 -7066
rect 465294 -7386 465914 -7302
rect 465294 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 465914 -7386
rect 465294 -7654 465914 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 474294 705798 474914 711590
rect 474294 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 474914 705798
rect 474294 705478 474914 705562
rect 474294 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 474914 705478
rect 474294 691954 474914 705242
rect 474294 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 474914 691954
rect 474294 691634 474914 691718
rect 474294 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 474914 691634
rect 474294 655954 474914 691398
rect 474294 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 474914 655954
rect 474294 655634 474914 655718
rect 474294 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 474914 655634
rect 474294 619954 474914 655398
rect 478794 706758 479414 711590
rect 478794 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 479414 706758
rect 478794 706438 479414 706522
rect 478794 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 479414 706438
rect 478794 696454 479414 706202
rect 478794 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 479414 696454
rect 478794 696134 479414 696218
rect 478794 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 479414 696134
rect 478794 660454 479414 695898
rect 478794 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 479414 660454
rect 478794 660134 479414 660218
rect 478794 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 479414 660134
rect 478794 642000 479414 659898
rect 483294 707718 483914 711590
rect 483294 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 483914 707718
rect 483294 707398 483914 707482
rect 483294 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 483914 707398
rect 483294 700954 483914 707162
rect 483294 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 483914 700954
rect 483294 700634 483914 700718
rect 483294 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 483914 700634
rect 483294 664954 483914 700398
rect 483294 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 483914 664954
rect 483294 664634 483914 664718
rect 483294 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 483914 664634
rect 483294 642000 483914 664398
rect 487794 708678 488414 711590
rect 487794 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 488414 708678
rect 487794 708358 488414 708442
rect 487794 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 488414 708358
rect 487794 669454 488414 708122
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 642000 488414 668898
rect 492294 709638 492914 711590
rect 492294 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 492914 709638
rect 492294 709318 492914 709402
rect 492294 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 492914 709318
rect 492294 673954 492914 709082
rect 492294 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 492914 673954
rect 492294 673634 492914 673718
rect 492294 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 492914 673634
rect 489683 659972 489749 659973
rect 489683 659908 489684 659972
rect 489748 659908 489749 659972
rect 489683 659907 489749 659908
rect 474294 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 474914 619954
rect 474294 619634 474914 619718
rect 474294 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 474914 619634
rect 474294 583954 474914 619398
rect 484208 615454 484528 615486
rect 484208 615218 484250 615454
rect 484486 615218 484528 615454
rect 484208 615134 484528 615218
rect 484208 614898 484250 615134
rect 484486 614898 484528 615134
rect 484208 614866 484528 614898
rect 474294 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 474914 583954
rect 474294 583634 474914 583718
rect 474294 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 474914 583634
rect 474294 547954 474914 583398
rect 474294 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 474914 547954
rect 474294 547634 474914 547718
rect 474294 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 474914 547634
rect 474294 511954 474914 547398
rect 478794 588454 479414 598000
rect 478794 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 479414 588454
rect 478794 588134 479414 588218
rect 478794 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 479414 588134
rect 478794 552454 479414 587898
rect 478794 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 479414 552454
rect 478794 552134 479414 552218
rect 478794 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 479414 552134
rect 478794 542000 479414 551898
rect 483294 592954 483914 598000
rect 483294 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 483914 592954
rect 483294 592634 483914 592718
rect 483294 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 483914 592634
rect 483294 556954 483914 592398
rect 483294 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 483914 556954
rect 483294 556634 483914 556718
rect 483294 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 483914 556634
rect 483294 542000 483914 556398
rect 487794 597454 488414 598000
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 542000 488414 560898
rect 489686 543690 489746 659907
rect 492294 642000 492914 673398
rect 496794 710598 497414 711590
rect 496794 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 497414 710598
rect 496794 710278 497414 710362
rect 496794 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 497414 710278
rect 496794 678454 497414 710042
rect 496794 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 497414 678454
rect 496794 678134 497414 678218
rect 496794 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 497414 678134
rect 496794 642361 497414 677898
rect 496794 642125 496826 642361
rect 497062 642125 497146 642361
rect 497382 642125 497414 642361
rect 496794 642000 497414 642125
rect 501294 711558 501914 711590
rect 501294 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 501914 711558
rect 501294 711238 501914 711322
rect 501294 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 501914 711238
rect 501294 682954 501914 711002
rect 501294 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 501914 682954
rect 501294 682634 501914 682718
rect 501294 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 501914 682634
rect 501294 646954 501914 682398
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 502931 660244 502997 660245
rect 502931 660180 502932 660244
rect 502996 660180 502997 660244
rect 502931 660179 502997 660180
rect 501294 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 501914 646954
rect 501294 646634 501914 646718
rect 501294 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 501914 646634
rect 501294 642000 501914 646398
rect 499568 619954 499888 619986
rect 499568 619718 499610 619954
rect 499846 619718 499888 619954
rect 499568 619634 499888 619718
rect 499568 619398 499610 619634
rect 499846 619398 499888 619634
rect 499568 619366 499888 619398
rect 489867 543692 489933 543693
rect 489867 543690 489868 543692
rect 489686 543630 489868 543690
rect 489867 543628 489868 543630
rect 489932 543628 489933 543692
rect 489867 543627 489933 543628
rect 495939 541108 496005 541109
rect 495939 541044 495940 541108
rect 496004 541044 496005 541108
rect 495939 541043 496005 541044
rect 485635 539884 485701 539885
rect 485635 539820 485636 539884
rect 485700 539820 485701 539884
rect 485635 539819 485701 539820
rect 474294 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 474914 511954
rect 474294 511634 474914 511718
rect 474294 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 474914 511634
rect 474294 475954 474914 511398
rect 484208 507454 484528 507486
rect 484208 507218 484250 507454
rect 484486 507218 484528 507454
rect 484208 507134 484528 507218
rect 484208 506898 484250 507134
rect 484486 506898 484528 507134
rect 484208 506866 484528 506898
rect 474294 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 474914 475954
rect 474294 475634 474914 475718
rect 474294 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 474914 475634
rect 474294 439954 474914 475398
rect 474294 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 474914 439954
rect 474294 439634 474914 439718
rect 474294 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 474914 439634
rect 474294 403954 474914 439398
rect 474294 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 474914 403954
rect 474294 403634 474914 403718
rect 474294 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 474914 403634
rect 474294 367954 474914 403398
rect 474294 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 474914 367954
rect 474294 367634 474914 367718
rect 474294 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 474914 367634
rect 474294 331954 474914 367398
rect 474294 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 474914 331954
rect 474294 331634 474914 331718
rect 474294 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 474914 331634
rect 474294 295954 474914 331398
rect 474294 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 474914 295954
rect 474294 295634 474914 295718
rect 474294 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 474914 295634
rect 474294 259954 474914 295398
rect 474294 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 474914 259954
rect 474294 259634 474914 259718
rect 474294 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 474914 259634
rect 474294 223954 474914 259398
rect 474294 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 474914 223954
rect 474294 223634 474914 223718
rect 474294 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 474914 223634
rect 474294 187954 474914 223398
rect 474294 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 474914 187954
rect 474294 187634 474914 187718
rect 474294 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 474914 187634
rect 474294 151954 474914 187398
rect 474294 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 474914 151954
rect 474294 151634 474914 151718
rect 474294 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 474914 151634
rect 474294 115954 474914 151398
rect 474294 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 474914 115954
rect 474294 115634 474914 115718
rect 474294 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 474914 115634
rect 474294 79954 474914 115398
rect 474294 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 474914 79954
rect 474294 79634 474914 79718
rect 474294 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 474914 79634
rect 474294 43954 474914 79398
rect 474294 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 474914 43954
rect 474294 43634 474914 43718
rect 474294 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 474914 43634
rect 474294 7954 474914 43398
rect 474294 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 474914 7954
rect 474294 7634 474914 7718
rect 474294 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 474914 7634
rect 474294 -1306 474914 7398
rect 474294 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 474914 -1306
rect 474294 -1626 474914 -1542
rect 474294 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 474914 -1626
rect 474294 -7654 474914 -1862
rect 478794 480454 479414 498000
rect 478794 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 479414 480454
rect 478794 480134 479414 480218
rect 478794 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 479414 480134
rect 478794 444454 479414 479898
rect 478794 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 479414 444454
rect 478794 444134 479414 444218
rect 478794 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 479414 444134
rect 478794 408454 479414 443898
rect 478794 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 479414 408454
rect 478794 408134 479414 408218
rect 478794 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 479414 408134
rect 478794 372454 479414 407898
rect 478794 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 479414 372454
rect 478794 372134 479414 372218
rect 478794 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 479414 372134
rect 478794 336454 479414 371898
rect 478794 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 479414 336454
rect 478794 336134 479414 336218
rect 478794 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 479414 336134
rect 478794 300454 479414 335898
rect 478794 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 479414 300454
rect 478794 300134 479414 300218
rect 478794 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 479414 300134
rect 478794 264454 479414 299898
rect 478794 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 479414 264454
rect 478794 264134 479414 264218
rect 478794 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 479414 264134
rect 478794 228454 479414 263898
rect 478794 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 479414 228454
rect 478794 228134 479414 228218
rect 478794 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 479414 228134
rect 478794 192454 479414 227898
rect 478794 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 479414 192454
rect 478794 192134 479414 192218
rect 478794 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 479414 192134
rect 478794 156454 479414 191898
rect 478794 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 479414 156454
rect 478794 156134 479414 156218
rect 478794 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 479414 156134
rect 478794 120454 479414 155898
rect 478794 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 479414 120454
rect 478794 120134 479414 120218
rect 478794 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 479414 120134
rect 478794 84454 479414 119898
rect 478794 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 479414 84454
rect 478794 84134 479414 84218
rect 478794 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 479414 84134
rect 478794 48454 479414 83898
rect 478794 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 479414 48454
rect 478794 48134 479414 48218
rect 478794 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 479414 48134
rect 478794 12454 479414 47898
rect 478794 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 479414 12454
rect 478794 12134 479414 12218
rect 478794 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 479414 12134
rect 478794 -2266 479414 11898
rect 478794 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 479414 -2266
rect 478794 -2586 479414 -2502
rect 478794 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 479414 -2586
rect 478794 -7654 479414 -2822
rect 483294 484954 483914 498000
rect 485638 496909 485698 539819
rect 486371 539748 486437 539749
rect 486371 539684 486372 539748
rect 486436 539684 486437 539748
rect 486371 539683 486437 539684
rect 494651 539748 494717 539749
rect 494651 539684 494652 539748
rect 494716 539684 494717 539748
rect 494651 539683 494717 539684
rect 484347 496908 484413 496909
rect 484347 496844 484348 496908
rect 484412 496844 484413 496908
rect 484347 496843 484413 496844
rect 485635 496908 485701 496909
rect 485635 496844 485636 496908
rect 485700 496844 485701 496908
rect 485635 496843 485701 496844
rect 483294 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 483914 484954
rect 483294 484634 483914 484718
rect 483294 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 483914 484634
rect 483294 448954 483914 484398
rect 483294 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 483914 448954
rect 483294 448634 483914 448718
rect 483294 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 483914 448634
rect 483294 412954 483914 448398
rect 483294 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 483914 412954
rect 483294 412634 483914 412718
rect 483294 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 483914 412634
rect 483294 376954 483914 412398
rect 483294 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 483914 376954
rect 483294 376634 483914 376718
rect 483294 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 483914 376634
rect 483294 340954 483914 376398
rect 483294 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 483914 340954
rect 483294 340634 483914 340718
rect 483294 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 483914 340634
rect 483294 304954 483914 340398
rect 483294 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 483914 304954
rect 483294 304634 483914 304718
rect 483294 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 483914 304634
rect 483294 268954 483914 304398
rect 483294 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 483914 268954
rect 483294 268634 483914 268718
rect 483294 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 483914 268634
rect 483294 232954 483914 268398
rect 483294 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 483914 232954
rect 483294 232634 483914 232718
rect 483294 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 483914 232634
rect 483294 196954 483914 232398
rect 483294 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 483914 196954
rect 483294 196634 483914 196718
rect 483294 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 483914 196634
rect 483294 160954 483914 196398
rect 483294 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 483914 160954
rect 483294 160634 483914 160718
rect 483294 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 483914 160634
rect 483294 124954 483914 160398
rect 483294 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 483914 124954
rect 483294 124634 483914 124718
rect 483294 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 483914 124634
rect 483294 88954 483914 124398
rect 483294 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 483914 88954
rect 483294 88634 483914 88718
rect 483294 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 483914 88634
rect 483294 52954 483914 88398
rect 483294 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 483914 52954
rect 483294 52634 483914 52718
rect 483294 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 483914 52634
rect 483294 16954 483914 52398
rect 483294 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 483914 16954
rect 483294 16634 483914 16718
rect 483294 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 483914 16634
rect 483294 -3226 483914 16398
rect 484350 4997 484410 496843
rect 486374 281485 486434 539683
rect 487794 489454 488414 498000
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 486371 281484 486437 281485
rect 486371 281420 486372 281484
rect 486436 281420 486437 281484
rect 486371 281419 486437 281420
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 484347 4996 484413 4997
rect 484347 4932 484348 4996
rect 484412 4932 484413 4996
rect 484347 4931 484413 4932
rect 483294 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 483914 -3226
rect 483294 -3546 483914 -3462
rect 483294 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 483914 -3546
rect 483294 -7654 483914 -3782
rect 487794 -4186 488414 20898
rect 487794 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 488414 -4186
rect 487794 -4506 488414 -4422
rect 487794 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 488414 -4506
rect 487794 -7654 488414 -4742
rect 492294 493954 492914 498000
rect 492294 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 492914 493954
rect 492294 493634 492914 493718
rect 492294 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 492914 493634
rect 492294 457954 492914 493398
rect 492294 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 492914 457954
rect 492294 457634 492914 457718
rect 492294 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 492914 457634
rect 492294 421954 492914 457398
rect 492294 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 492914 421954
rect 492294 421634 492914 421718
rect 492294 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 492914 421634
rect 492294 385954 492914 421398
rect 492294 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 492914 385954
rect 492294 385634 492914 385718
rect 492294 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 492914 385634
rect 492294 349954 492914 385398
rect 492294 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 492914 349954
rect 492294 349634 492914 349718
rect 492294 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 492914 349634
rect 492294 313954 492914 349398
rect 492294 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 492914 313954
rect 492294 313634 492914 313718
rect 492294 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 492914 313634
rect 492294 277954 492914 313398
rect 492294 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 492914 277954
rect 492294 277634 492914 277718
rect 492294 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 492914 277634
rect 492294 241954 492914 277398
rect 492294 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 492914 241954
rect 492294 241634 492914 241718
rect 492294 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 492914 241634
rect 492294 205954 492914 241398
rect 492294 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 492914 205954
rect 492294 205634 492914 205718
rect 492294 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 492914 205634
rect 492294 169954 492914 205398
rect 492294 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 492914 169954
rect 492294 169634 492914 169718
rect 492294 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 492914 169634
rect 492294 133954 492914 169398
rect 492294 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 492914 133954
rect 492294 133634 492914 133718
rect 492294 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 492914 133634
rect 492294 97954 492914 133398
rect 492294 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 492914 97954
rect 492294 97634 492914 97718
rect 492294 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 492914 97634
rect 492294 61954 492914 97398
rect 492294 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 492914 61954
rect 492294 61634 492914 61718
rect 492294 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 492914 61634
rect 492294 25954 492914 61398
rect 492294 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 492914 25954
rect 492294 25634 492914 25718
rect 492294 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 492914 25634
rect 492294 -5146 492914 25398
rect 494654 7581 494714 539683
rect 495942 499629 496002 541043
rect 502195 539748 502261 539749
rect 502195 539684 502196 539748
rect 502260 539684 502261 539748
rect 502195 539683 502261 539684
rect 499568 511954 499888 511986
rect 499568 511718 499610 511954
rect 499846 511718 499888 511954
rect 499568 511634 499888 511718
rect 499568 511398 499610 511634
rect 499846 511398 499888 511634
rect 499568 511366 499888 511398
rect 495939 499628 496005 499629
rect 495939 499564 495940 499628
rect 496004 499564 496005 499628
rect 495939 499563 496005 499564
rect 496794 462454 497414 498000
rect 496794 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 497414 462454
rect 496794 462134 497414 462218
rect 496794 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 497414 462134
rect 496794 426454 497414 461898
rect 496794 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 497414 426454
rect 496794 426134 497414 426218
rect 496794 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 497414 426134
rect 496794 390454 497414 425898
rect 496794 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 497414 390454
rect 496794 390134 497414 390218
rect 496794 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 497414 390134
rect 496794 354454 497414 389898
rect 496794 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 497414 354454
rect 496794 354134 497414 354218
rect 496794 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 497414 354134
rect 496794 318454 497414 353898
rect 496794 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 497414 318454
rect 496794 318134 497414 318218
rect 496794 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 497414 318134
rect 496794 282454 497414 317898
rect 496794 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 497414 282454
rect 496794 282134 497414 282218
rect 496794 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 497414 282134
rect 496794 246454 497414 281898
rect 496794 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 497414 246454
rect 496794 246134 497414 246218
rect 496794 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 497414 246134
rect 496794 210454 497414 245898
rect 496794 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 497414 210454
rect 496794 210134 497414 210218
rect 496794 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 497414 210134
rect 496794 174454 497414 209898
rect 496794 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 497414 174454
rect 496794 174134 497414 174218
rect 496794 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 497414 174134
rect 496794 138454 497414 173898
rect 496794 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 497414 138454
rect 496794 138134 497414 138218
rect 496794 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 497414 138134
rect 496794 102454 497414 137898
rect 496794 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 497414 102454
rect 496794 102134 497414 102218
rect 496794 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 497414 102134
rect 496794 66454 497414 101898
rect 496794 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 497414 66454
rect 496794 66134 497414 66218
rect 496794 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 497414 66134
rect 496794 30454 497414 65898
rect 496794 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 497414 30454
rect 496794 30134 497414 30218
rect 496794 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 497414 30134
rect 494651 7580 494717 7581
rect 494651 7516 494652 7580
rect 494716 7516 494717 7580
rect 494651 7515 494717 7516
rect 492294 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 492914 -5146
rect 492294 -5466 492914 -5382
rect 492294 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 492914 -5466
rect 492294 -7654 492914 -5702
rect 496794 -6106 497414 29898
rect 496794 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 497414 -6106
rect 496794 -6426 497414 -6342
rect 496794 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 497414 -6426
rect 496794 -7654 497414 -6662
rect 501294 466954 501914 498000
rect 501294 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 501914 466954
rect 501294 466634 501914 466718
rect 501294 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 501914 466634
rect 501294 430954 501914 466398
rect 501294 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 501914 430954
rect 501294 430634 501914 430718
rect 501294 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 501914 430634
rect 501294 394954 501914 430398
rect 501294 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 501914 394954
rect 501294 394634 501914 394718
rect 501294 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 501914 394634
rect 501294 358954 501914 394398
rect 501294 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 501914 358954
rect 501294 358634 501914 358718
rect 501294 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 501914 358634
rect 501294 322954 501914 358398
rect 501294 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 501914 322954
rect 501294 322634 501914 322718
rect 501294 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 501914 322634
rect 501294 286954 501914 322398
rect 501294 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 501914 286954
rect 501294 286634 501914 286718
rect 501294 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 501914 286634
rect 501294 250954 501914 286398
rect 501294 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 501914 250954
rect 501294 250634 501914 250718
rect 501294 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 501914 250634
rect 501294 214954 501914 250398
rect 501294 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 501914 214954
rect 501294 214634 501914 214718
rect 501294 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 501914 214634
rect 501294 178954 501914 214398
rect 501294 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 501914 178954
rect 501294 178634 501914 178718
rect 501294 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 501914 178634
rect 501294 142954 501914 178398
rect 501294 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 501914 142954
rect 501294 142634 501914 142718
rect 501294 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 501914 142634
rect 501294 106954 501914 142398
rect 501294 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 501914 106954
rect 501294 106634 501914 106718
rect 501294 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 501914 106634
rect 501294 70954 501914 106398
rect 501294 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 501914 70954
rect 501294 70634 501914 70718
rect 501294 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 501914 70634
rect 501294 34954 501914 70398
rect 501294 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 501914 34954
rect 501294 34634 501914 34718
rect 501294 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 501914 34634
rect 501294 -7066 501914 34398
rect 502198 3501 502258 539683
rect 502934 499901 502994 660179
rect 505794 651454 506414 686898
rect 510294 705798 510914 711590
rect 510294 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 510914 705798
rect 510294 705478 510914 705562
rect 510294 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 510914 705478
rect 510294 691954 510914 705242
rect 510294 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 510914 691954
rect 510294 691634 510914 691718
rect 510294 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 510914 691634
rect 508451 660244 508517 660245
rect 508451 660180 508452 660244
rect 508516 660180 508517 660244
rect 508451 660179 508517 660180
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 642000 506414 650898
rect 505794 579454 506414 598000
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 508454 543557 508514 660179
rect 510294 655954 510914 691398
rect 510294 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 510914 655954
rect 510294 655634 510914 655718
rect 510294 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 510914 655634
rect 510294 642000 510914 655398
rect 514794 706758 515414 711590
rect 514794 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 515414 706758
rect 514794 706438 515414 706522
rect 514794 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 515414 706438
rect 514794 696454 515414 706202
rect 514794 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 515414 696454
rect 514794 696134 515414 696218
rect 514794 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 515414 696134
rect 514794 660454 515414 695898
rect 514794 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 515414 660454
rect 514794 660134 515414 660218
rect 514794 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 515414 660134
rect 514794 642000 515414 659898
rect 519294 707718 519914 711590
rect 519294 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 519914 707718
rect 519294 707398 519914 707482
rect 519294 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 519914 707398
rect 519294 700954 519914 707162
rect 519294 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 519914 700954
rect 519294 700634 519914 700718
rect 519294 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 519914 700634
rect 519294 664954 519914 700398
rect 519294 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 519914 664954
rect 519294 664634 519914 664718
rect 519294 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 519914 664634
rect 519294 642000 519914 664398
rect 523794 708678 524414 711590
rect 523794 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 524414 708678
rect 523794 708358 524414 708442
rect 523794 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 524414 708358
rect 523794 669454 524414 708122
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 642000 524414 668898
rect 528294 709638 528914 711590
rect 528294 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 528914 709638
rect 528294 709318 528914 709402
rect 528294 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 528914 709318
rect 528294 673954 528914 709082
rect 528294 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 528914 673954
rect 528294 673634 528914 673718
rect 528294 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 528914 673634
rect 528294 637954 528914 673398
rect 528294 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 528914 637954
rect 528294 637634 528914 637718
rect 528294 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 528914 637634
rect 514928 615454 515248 615486
rect 514928 615218 514970 615454
rect 515206 615218 515248 615454
rect 514928 615134 515248 615218
rect 514928 614898 514970 615134
rect 515206 614898 515248 615134
rect 514928 614866 515248 614898
rect 528294 601954 528914 637398
rect 528294 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 528914 601954
rect 528294 601634 528914 601718
rect 528294 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 528914 601634
rect 510294 583954 510914 598000
rect 510294 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 510914 583954
rect 510294 583634 510914 583718
rect 510294 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 510914 583634
rect 510294 547954 510914 583398
rect 510294 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 510914 547954
rect 510294 547634 510914 547718
rect 510294 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 510914 547634
rect 508451 543556 508517 543557
rect 508451 543492 508452 543556
rect 508516 543492 508517 543556
rect 508451 543491 508517 543492
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 542000 506414 542898
rect 510294 542000 510914 547398
rect 514794 588454 515414 598000
rect 514794 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 515414 588454
rect 514794 588134 515414 588218
rect 514794 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 515414 588134
rect 514794 552454 515414 587898
rect 514794 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 515414 552454
rect 514794 552134 515414 552218
rect 514794 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 515414 552134
rect 514794 542000 515414 551898
rect 519294 592954 519914 598000
rect 519294 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 519914 592954
rect 519294 592634 519914 592718
rect 519294 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 519914 592634
rect 519294 556954 519914 592398
rect 519294 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 519914 556954
rect 519294 556634 519914 556718
rect 519294 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 519914 556634
rect 519294 542000 519914 556398
rect 523794 597454 524414 598000
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 542000 524414 560898
rect 528294 565954 528914 601398
rect 528294 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 528914 565954
rect 528294 565634 528914 565718
rect 528294 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 528914 565634
rect 511211 541108 511277 541109
rect 511211 541044 511212 541108
rect 511276 541044 511277 541108
rect 511211 541043 511277 541044
rect 505507 539748 505573 539749
rect 505507 539684 505508 539748
rect 505572 539684 505573 539748
rect 505507 539683 505573 539684
rect 502931 499900 502997 499901
rect 502931 499836 502932 499900
rect 502996 499836 502997 499900
rect 502931 499835 502997 499836
rect 505510 4045 505570 539683
rect 505794 471454 506414 498000
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505507 4044 505573 4045
rect 505507 3980 505508 4044
rect 505572 3980 505573 4044
rect 505507 3979 505573 3980
rect 502195 3500 502261 3501
rect 502195 3436 502196 3500
rect 502260 3436 502261 3500
rect 502195 3435 502261 3436
rect 505794 3454 506414 38898
rect 501294 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 501914 -7066
rect 501294 -7386 501914 -7302
rect 501294 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 501914 -7386
rect 501294 -7654 501914 -7622
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 510294 475954 510914 498000
rect 510294 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 510914 475954
rect 510294 475634 510914 475718
rect 510294 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 510914 475634
rect 510294 439954 510914 475398
rect 510294 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 510914 439954
rect 510294 439634 510914 439718
rect 510294 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 510914 439634
rect 510294 403954 510914 439398
rect 510294 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 510914 403954
rect 510294 403634 510914 403718
rect 510294 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 510914 403634
rect 510294 367954 510914 403398
rect 510294 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 510914 367954
rect 510294 367634 510914 367718
rect 510294 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 510914 367634
rect 510294 331954 510914 367398
rect 510294 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 510914 331954
rect 510294 331634 510914 331718
rect 510294 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 510914 331634
rect 510294 295954 510914 331398
rect 510294 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 510914 295954
rect 510294 295634 510914 295718
rect 510294 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 510914 295634
rect 510294 259954 510914 295398
rect 510294 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 510914 259954
rect 510294 259634 510914 259718
rect 510294 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 510914 259634
rect 510294 223954 510914 259398
rect 510294 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 510914 223954
rect 510294 223634 510914 223718
rect 510294 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 510914 223634
rect 510294 187954 510914 223398
rect 510294 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 510914 187954
rect 510294 187634 510914 187718
rect 510294 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 510914 187634
rect 510294 151954 510914 187398
rect 510294 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 510914 151954
rect 510294 151634 510914 151718
rect 510294 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 510914 151634
rect 510294 115954 510914 151398
rect 510294 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 510914 115954
rect 510294 115634 510914 115718
rect 510294 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 510914 115634
rect 510294 79954 510914 115398
rect 510294 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 510914 79954
rect 510294 79634 510914 79718
rect 510294 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 510914 79634
rect 510294 43954 510914 79398
rect 510294 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 510914 43954
rect 510294 43634 510914 43718
rect 510294 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 510914 43634
rect 510294 7954 510914 43398
rect 510294 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 510914 7954
rect 510294 7634 510914 7718
rect 510294 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 510914 7634
rect 510294 -1306 510914 7398
rect 511214 3365 511274 541043
rect 512499 539884 512565 539885
rect 512499 539820 512500 539884
rect 512564 539820 512565 539884
rect 512499 539819 512565 539820
rect 512502 6221 512562 539819
rect 516363 539748 516429 539749
rect 516363 539684 516364 539748
rect 516428 539684 516429 539748
rect 516363 539683 516429 539684
rect 514928 507454 515248 507486
rect 514928 507218 514970 507454
rect 515206 507218 515248 507454
rect 514928 507134 515248 507218
rect 514928 506898 514970 507134
rect 515206 506898 515248 507134
rect 514928 506866 515248 506898
rect 514794 480454 515414 498000
rect 514794 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 515414 480454
rect 514794 480134 515414 480218
rect 514794 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 515414 480134
rect 514794 444454 515414 479898
rect 514794 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 515414 444454
rect 514794 444134 515414 444218
rect 514794 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 515414 444134
rect 514794 408454 515414 443898
rect 514794 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 515414 408454
rect 514794 408134 515414 408218
rect 514794 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 515414 408134
rect 514794 372454 515414 407898
rect 514794 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 515414 372454
rect 514794 372134 515414 372218
rect 514794 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 515414 372134
rect 514794 336454 515414 371898
rect 514794 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 515414 336454
rect 514794 336134 515414 336218
rect 514794 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 515414 336134
rect 514794 300454 515414 335898
rect 514794 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 515414 300454
rect 514794 300134 515414 300218
rect 514794 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 515414 300134
rect 514794 264454 515414 299898
rect 514794 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 515414 264454
rect 514794 264134 515414 264218
rect 514794 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 515414 264134
rect 514794 228454 515414 263898
rect 514794 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 515414 228454
rect 514794 228134 515414 228218
rect 514794 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 515414 228134
rect 514794 192454 515414 227898
rect 514794 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 515414 192454
rect 514794 192134 515414 192218
rect 514794 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 515414 192134
rect 514794 156454 515414 191898
rect 514794 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 515414 156454
rect 514794 156134 515414 156218
rect 514794 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 515414 156134
rect 514794 120454 515414 155898
rect 514794 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 515414 120454
rect 514794 120134 515414 120218
rect 514794 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 515414 120134
rect 514794 84454 515414 119898
rect 514794 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 515414 84454
rect 514794 84134 515414 84218
rect 514794 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 515414 84134
rect 514794 48454 515414 83898
rect 514794 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 515414 48454
rect 514794 48134 515414 48218
rect 514794 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 515414 48134
rect 514794 12454 515414 47898
rect 514794 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 515414 12454
rect 514794 12134 515414 12218
rect 514794 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 515414 12134
rect 512499 6220 512565 6221
rect 512499 6156 512500 6220
rect 512564 6156 512565 6220
rect 512499 6155 512565 6156
rect 511211 3364 511277 3365
rect 511211 3300 511212 3364
rect 511276 3300 511277 3364
rect 511211 3299 511277 3300
rect 510294 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 510914 -1306
rect 510294 -1626 510914 -1542
rect 510294 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 510914 -1626
rect 510294 -7654 510914 -1862
rect 514794 -2266 515414 11898
rect 516366 3501 516426 539683
rect 521883 538524 521949 538525
rect 521883 538460 521884 538524
rect 521948 538460 521949 538524
rect 521883 538459 521949 538460
rect 519307 533900 519373 533901
rect 519307 533836 519308 533900
rect 519372 533836 519373 533900
rect 519307 533835 519373 533836
rect 519310 528570 519370 533835
rect 518942 528510 519370 528570
rect 518942 4861 519002 528510
rect 519307 523428 519373 523429
rect 519307 523364 519308 523428
rect 519372 523364 519373 523428
rect 519307 523363 519373 523364
rect 519310 509250 519370 523363
rect 519126 509190 519370 509250
rect 519126 224229 519186 509190
rect 521699 503028 521765 503029
rect 521699 502964 521700 503028
rect 521764 502964 521765 503028
rect 521699 502963 521765 502964
rect 519294 484954 519914 498000
rect 519294 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 519914 484954
rect 519294 484634 519914 484718
rect 519294 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 519914 484634
rect 519294 448954 519914 484398
rect 519294 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 519914 448954
rect 519294 448634 519914 448718
rect 519294 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 519914 448634
rect 519294 412954 519914 448398
rect 519294 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 519914 412954
rect 519294 412634 519914 412718
rect 519294 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 519914 412634
rect 519294 376954 519914 412398
rect 519294 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 519914 376954
rect 519294 376634 519914 376718
rect 519294 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 519914 376634
rect 519294 340954 519914 376398
rect 519294 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 519914 340954
rect 519294 340634 519914 340718
rect 519294 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 519914 340634
rect 519294 304954 519914 340398
rect 519294 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 519914 304954
rect 519294 304634 519914 304718
rect 519294 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 519914 304634
rect 519294 268954 519914 304398
rect 519294 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 519914 268954
rect 519294 268634 519914 268718
rect 519294 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 519914 268634
rect 519294 232954 519914 268398
rect 519294 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 519914 232954
rect 519294 232634 519914 232718
rect 519294 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 519914 232634
rect 519123 224228 519189 224229
rect 519123 224164 519124 224228
rect 519188 224164 519189 224228
rect 519123 224163 519189 224164
rect 519294 196954 519914 232398
rect 519294 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 519914 196954
rect 519294 196634 519914 196718
rect 519294 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 519914 196634
rect 519294 160954 519914 196398
rect 519294 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 519914 160954
rect 519294 160634 519914 160718
rect 519294 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 519914 160634
rect 519294 124954 519914 160398
rect 519294 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 519914 124954
rect 519294 124634 519914 124718
rect 519294 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 519914 124634
rect 519294 88954 519914 124398
rect 519294 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 519914 88954
rect 519294 88634 519914 88718
rect 519294 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 519914 88634
rect 519294 52954 519914 88398
rect 519294 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 519914 52954
rect 519294 52634 519914 52718
rect 519294 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 519914 52634
rect 519294 16954 519914 52398
rect 519294 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 519914 16954
rect 519294 16634 519914 16718
rect 519294 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 519914 16634
rect 518939 4860 519005 4861
rect 518939 4796 518940 4860
rect 519004 4796 519005 4860
rect 518939 4795 519005 4796
rect 516363 3500 516429 3501
rect 516363 3436 516364 3500
rect 516428 3436 516429 3500
rect 516363 3435 516429 3436
rect 514794 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 515414 -2266
rect 514794 -2586 515414 -2502
rect 514794 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 515414 -2586
rect 514794 -7654 515414 -2822
rect 519294 -3226 519914 16398
rect 521702 8941 521762 502963
rect 521886 224365 521946 538459
rect 522067 532812 522133 532813
rect 522067 532748 522068 532812
rect 522132 532748 522133 532812
rect 522067 532747 522133 532748
rect 522070 226949 522130 532747
rect 528294 529954 528914 565398
rect 528294 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 528914 529954
rect 528294 529634 528914 529718
rect 528294 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 528914 529634
rect 523794 489454 524414 498000
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 522067 226948 522133 226949
rect 522067 226884 522068 226948
rect 522132 226884 522133 226948
rect 522067 226883 522133 226884
rect 521883 224364 521949 224365
rect 521883 224300 521884 224364
rect 521948 224300 521949 224364
rect 521883 224299 521949 224300
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 521699 8940 521765 8941
rect 521699 8876 521700 8940
rect 521764 8876 521765 8940
rect 521699 8875 521765 8876
rect 519294 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 519914 -3226
rect 519294 -3546 519914 -3462
rect 519294 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 519914 -3546
rect 519294 -7654 519914 -3782
rect 523794 -4186 524414 20898
rect 523794 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 524414 -4186
rect 523794 -4506 524414 -4422
rect 523794 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 524414 -4506
rect 523794 -7654 524414 -4742
rect 528294 493954 528914 529398
rect 528294 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 528914 493954
rect 528294 493634 528914 493718
rect 528294 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 528914 493634
rect 528294 457954 528914 493398
rect 528294 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 528914 457954
rect 528294 457634 528914 457718
rect 528294 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 528914 457634
rect 528294 421954 528914 457398
rect 528294 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 528914 421954
rect 528294 421634 528914 421718
rect 528294 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 528914 421634
rect 528294 385954 528914 421398
rect 528294 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 528914 385954
rect 528294 385634 528914 385718
rect 528294 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 528914 385634
rect 528294 349954 528914 385398
rect 528294 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 528914 349954
rect 528294 349634 528914 349718
rect 528294 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 528914 349634
rect 528294 313954 528914 349398
rect 528294 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 528914 313954
rect 528294 313634 528914 313718
rect 528294 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 528914 313634
rect 528294 277954 528914 313398
rect 528294 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 528914 277954
rect 528294 277634 528914 277718
rect 528294 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 528914 277634
rect 528294 241954 528914 277398
rect 528294 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 528914 241954
rect 528294 241634 528914 241718
rect 528294 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 528914 241634
rect 528294 205954 528914 241398
rect 528294 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 528914 205954
rect 528294 205634 528914 205718
rect 528294 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 528914 205634
rect 528294 169954 528914 205398
rect 528294 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 528914 169954
rect 528294 169634 528914 169718
rect 528294 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 528914 169634
rect 528294 133954 528914 169398
rect 528294 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 528914 133954
rect 528294 133634 528914 133718
rect 528294 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 528914 133634
rect 528294 97954 528914 133398
rect 528294 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 528914 97954
rect 528294 97634 528914 97718
rect 528294 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 528914 97634
rect 528294 61954 528914 97398
rect 528294 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 528914 61954
rect 528294 61634 528914 61718
rect 528294 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 528914 61634
rect 528294 25954 528914 61398
rect 528294 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 528914 25954
rect 528294 25634 528914 25718
rect 528294 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 528914 25634
rect 528294 -5146 528914 25398
rect 528294 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 528914 -5146
rect 528294 -5466 528914 -5382
rect 528294 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 528914 -5466
rect 528294 -7654 528914 -5702
rect 532794 710598 533414 711590
rect 532794 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 533414 710598
rect 532794 710278 533414 710362
rect 532794 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 533414 710278
rect 532794 678454 533414 710042
rect 532794 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 533414 678454
rect 532794 678134 533414 678218
rect 532794 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 533414 678134
rect 532794 642454 533414 677898
rect 532794 642218 532826 642454
rect 533062 642218 533146 642454
rect 533382 642218 533414 642454
rect 532794 642134 533414 642218
rect 532794 641898 532826 642134
rect 533062 641898 533146 642134
rect 533382 641898 533414 642134
rect 532794 606454 533414 641898
rect 532794 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 533414 606454
rect 532794 606134 533414 606218
rect 532794 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 533414 606134
rect 532794 570454 533414 605898
rect 532794 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 533414 570454
rect 532794 570134 533414 570218
rect 532794 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 533414 570134
rect 532794 534454 533414 569898
rect 532794 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 533414 534454
rect 532794 534134 533414 534218
rect 532794 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 533414 534134
rect 532794 498454 533414 533898
rect 532794 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 533414 498454
rect 532794 498134 533414 498218
rect 532794 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 533414 498134
rect 532794 462454 533414 497898
rect 532794 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 533414 462454
rect 532794 462134 533414 462218
rect 532794 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 533414 462134
rect 532794 426454 533414 461898
rect 532794 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 533414 426454
rect 532794 426134 533414 426218
rect 532794 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 533414 426134
rect 532794 390454 533414 425898
rect 532794 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 533414 390454
rect 532794 390134 533414 390218
rect 532794 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 533414 390134
rect 532794 354454 533414 389898
rect 532794 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 533414 354454
rect 532794 354134 533414 354218
rect 532794 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 533414 354134
rect 532794 318454 533414 353898
rect 532794 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 533414 318454
rect 532794 318134 533414 318218
rect 532794 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 533414 318134
rect 532794 282454 533414 317898
rect 532794 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 533414 282454
rect 532794 282134 533414 282218
rect 532794 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 533414 282134
rect 532794 246454 533414 281898
rect 532794 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 533414 246454
rect 532794 246134 533414 246218
rect 532794 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 533414 246134
rect 532794 210454 533414 245898
rect 532794 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 533414 210454
rect 532794 210134 533414 210218
rect 532794 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 533414 210134
rect 532794 174454 533414 209898
rect 532794 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 533414 174454
rect 532794 174134 533414 174218
rect 532794 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 533414 174134
rect 532794 138454 533414 173898
rect 532794 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 533414 138454
rect 532794 138134 533414 138218
rect 532794 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 533414 138134
rect 532794 102454 533414 137898
rect 532794 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 533414 102454
rect 532794 102134 533414 102218
rect 532794 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 533414 102134
rect 532794 66454 533414 101898
rect 532794 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 533414 66454
rect 532794 66134 533414 66218
rect 532794 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 533414 66134
rect 532794 30454 533414 65898
rect 532794 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 533414 30454
rect 532794 30134 533414 30218
rect 532794 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 533414 30134
rect 532794 -6106 533414 29898
rect 532794 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 533414 -6106
rect 532794 -6426 533414 -6342
rect 532794 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 533414 -6426
rect 532794 -7654 533414 -6662
rect 537294 711558 537914 711590
rect 537294 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 537914 711558
rect 537294 711238 537914 711322
rect 537294 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 537914 711238
rect 537294 682954 537914 711002
rect 537294 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 537914 682954
rect 537294 682634 537914 682718
rect 537294 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 537914 682634
rect 537294 646954 537914 682398
rect 537294 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 537914 646954
rect 537294 646634 537914 646718
rect 537294 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 537914 646634
rect 537294 610954 537914 646398
rect 537294 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 537914 610954
rect 537294 610634 537914 610718
rect 537294 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 537914 610634
rect 537294 574954 537914 610398
rect 537294 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 537914 574954
rect 537294 574634 537914 574718
rect 537294 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 537914 574634
rect 537294 538954 537914 574398
rect 537294 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 537914 538954
rect 537294 538634 537914 538718
rect 537294 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 537914 538634
rect 537294 502954 537914 538398
rect 537294 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 537914 502954
rect 537294 502634 537914 502718
rect 537294 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 537914 502634
rect 537294 466954 537914 502398
rect 537294 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 537914 466954
rect 537294 466634 537914 466718
rect 537294 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 537914 466634
rect 537294 430954 537914 466398
rect 537294 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 537914 430954
rect 537294 430634 537914 430718
rect 537294 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 537914 430634
rect 537294 394954 537914 430398
rect 537294 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 537914 394954
rect 537294 394634 537914 394718
rect 537294 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 537914 394634
rect 537294 358954 537914 394398
rect 537294 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 537914 358954
rect 537294 358634 537914 358718
rect 537294 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 537914 358634
rect 537294 322954 537914 358398
rect 537294 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 537914 322954
rect 537294 322634 537914 322718
rect 537294 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 537914 322634
rect 537294 286954 537914 322398
rect 537294 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 537914 286954
rect 537294 286634 537914 286718
rect 537294 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 537914 286634
rect 537294 250954 537914 286398
rect 537294 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 537914 250954
rect 537294 250634 537914 250718
rect 537294 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 537914 250634
rect 537294 214954 537914 250398
rect 537294 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 537914 214954
rect 537294 214634 537914 214718
rect 537294 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 537914 214634
rect 537294 178954 537914 214398
rect 537294 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 537914 178954
rect 537294 178634 537914 178718
rect 537294 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 537914 178634
rect 537294 142954 537914 178398
rect 537294 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 537914 142954
rect 537294 142634 537914 142718
rect 537294 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 537914 142634
rect 537294 106954 537914 142398
rect 537294 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 537914 106954
rect 537294 106634 537914 106718
rect 537294 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 537914 106634
rect 537294 70954 537914 106398
rect 537294 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 537914 70954
rect 537294 70634 537914 70718
rect 537294 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 537914 70634
rect 537294 34954 537914 70398
rect 537294 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 537914 34954
rect 537294 34634 537914 34718
rect 537294 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 537914 34634
rect 537294 -7066 537914 34398
rect 537294 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 537914 -7066
rect 537294 -7386 537914 -7302
rect 537294 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 537914 -7386
rect 537294 -7654 537914 -7622
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 546294 705798 546914 711590
rect 546294 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 546914 705798
rect 546294 705478 546914 705562
rect 546294 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 546914 705478
rect 546294 691954 546914 705242
rect 546294 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 546914 691954
rect 546294 691634 546914 691718
rect 546294 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 546914 691634
rect 546294 655954 546914 691398
rect 546294 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 546914 655954
rect 546294 655634 546914 655718
rect 546294 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 546914 655634
rect 546294 619954 546914 655398
rect 546294 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 546914 619954
rect 546294 619634 546914 619718
rect 546294 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 546914 619634
rect 546294 583954 546914 619398
rect 546294 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 546914 583954
rect 546294 583634 546914 583718
rect 546294 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 546914 583634
rect 546294 547954 546914 583398
rect 546294 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 546914 547954
rect 546294 547634 546914 547718
rect 546294 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 546914 547634
rect 546294 511954 546914 547398
rect 546294 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 546914 511954
rect 546294 511634 546914 511718
rect 546294 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 546914 511634
rect 546294 475954 546914 511398
rect 546294 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 546914 475954
rect 546294 475634 546914 475718
rect 546294 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 546914 475634
rect 546294 439954 546914 475398
rect 546294 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 546914 439954
rect 546294 439634 546914 439718
rect 546294 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 546914 439634
rect 546294 403954 546914 439398
rect 546294 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 546914 403954
rect 546294 403634 546914 403718
rect 546294 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 546914 403634
rect 546294 367954 546914 403398
rect 546294 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 546914 367954
rect 546294 367634 546914 367718
rect 546294 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 546914 367634
rect 546294 331954 546914 367398
rect 546294 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 546914 331954
rect 546294 331634 546914 331718
rect 546294 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 546914 331634
rect 546294 295954 546914 331398
rect 546294 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 546914 295954
rect 546294 295634 546914 295718
rect 546294 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 546914 295634
rect 546294 259954 546914 295398
rect 546294 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 546914 259954
rect 546294 259634 546914 259718
rect 546294 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 546914 259634
rect 546294 223954 546914 259398
rect 546294 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 546914 223954
rect 546294 223634 546914 223718
rect 546294 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 546914 223634
rect 546294 187954 546914 223398
rect 546294 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 546914 187954
rect 546294 187634 546914 187718
rect 546294 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 546914 187634
rect 546294 151954 546914 187398
rect 546294 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 546914 151954
rect 546294 151634 546914 151718
rect 546294 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 546914 151634
rect 546294 115954 546914 151398
rect 546294 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 546914 115954
rect 546294 115634 546914 115718
rect 546294 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 546914 115634
rect 546294 79954 546914 115398
rect 546294 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 546914 79954
rect 546294 79634 546914 79718
rect 546294 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 546914 79634
rect 546294 43954 546914 79398
rect 546294 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 546914 43954
rect 546294 43634 546914 43718
rect 546294 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 546914 43634
rect 546294 7954 546914 43398
rect 546294 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 546914 7954
rect 546294 7634 546914 7718
rect 546294 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 546914 7634
rect 546294 -1306 546914 7398
rect 546294 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 546914 -1306
rect 546294 -1626 546914 -1542
rect 546294 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 546914 -1626
rect 546294 -7654 546914 -1862
rect 550794 706758 551414 711590
rect 550794 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 551414 706758
rect 550794 706438 551414 706522
rect 550794 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 551414 706438
rect 550794 696454 551414 706202
rect 550794 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 551414 696454
rect 550794 696134 551414 696218
rect 550794 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 551414 696134
rect 550794 660454 551414 695898
rect 550794 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 551414 660454
rect 550794 660134 551414 660218
rect 550794 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 551414 660134
rect 550794 624454 551414 659898
rect 550794 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 551414 624454
rect 550794 624134 551414 624218
rect 550794 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 551414 624134
rect 550794 588454 551414 623898
rect 550794 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 551414 588454
rect 550794 588134 551414 588218
rect 550794 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 551414 588134
rect 550794 552454 551414 587898
rect 550794 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 551414 552454
rect 550794 552134 551414 552218
rect 550794 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 551414 552134
rect 550794 516454 551414 551898
rect 550794 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 551414 516454
rect 550794 516134 551414 516218
rect 550794 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 551414 516134
rect 550794 480454 551414 515898
rect 550794 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 551414 480454
rect 550794 480134 551414 480218
rect 550794 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 551414 480134
rect 550794 444454 551414 479898
rect 550794 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 551414 444454
rect 550794 444134 551414 444218
rect 550794 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 551414 444134
rect 550794 408454 551414 443898
rect 550794 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 551414 408454
rect 550794 408134 551414 408218
rect 550794 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 551414 408134
rect 550794 372454 551414 407898
rect 550794 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 551414 372454
rect 550794 372134 551414 372218
rect 550794 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 551414 372134
rect 550794 336454 551414 371898
rect 550794 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 551414 336454
rect 550794 336134 551414 336218
rect 550794 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 551414 336134
rect 550794 300454 551414 335898
rect 550794 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 551414 300454
rect 550794 300134 551414 300218
rect 550794 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 551414 300134
rect 550794 264454 551414 299898
rect 550794 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 551414 264454
rect 550794 264134 551414 264218
rect 550794 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 551414 264134
rect 550794 228454 551414 263898
rect 550794 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 551414 228454
rect 550794 228134 551414 228218
rect 550794 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 551414 228134
rect 550794 192454 551414 227898
rect 550794 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 551414 192454
rect 550794 192134 551414 192218
rect 550794 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 551414 192134
rect 550794 156454 551414 191898
rect 550794 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 551414 156454
rect 550794 156134 551414 156218
rect 550794 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 551414 156134
rect 550794 120454 551414 155898
rect 550794 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 551414 120454
rect 550794 120134 551414 120218
rect 550794 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 551414 120134
rect 550794 84454 551414 119898
rect 550794 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 551414 84454
rect 550794 84134 551414 84218
rect 550794 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 551414 84134
rect 550794 48454 551414 83898
rect 550794 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 551414 48454
rect 550794 48134 551414 48218
rect 550794 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 551414 48134
rect 550794 12454 551414 47898
rect 550794 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 551414 12454
rect 550794 12134 551414 12218
rect 550794 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 551414 12134
rect 550794 -2266 551414 11898
rect 550794 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 551414 -2266
rect 550794 -2586 551414 -2502
rect 550794 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 551414 -2586
rect 550794 -7654 551414 -2822
rect 555294 707718 555914 711590
rect 555294 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 555914 707718
rect 555294 707398 555914 707482
rect 555294 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 555914 707398
rect 555294 700954 555914 707162
rect 555294 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 555914 700954
rect 555294 700634 555914 700718
rect 555294 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 555914 700634
rect 555294 664954 555914 700398
rect 555294 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 555914 664954
rect 555294 664634 555914 664718
rect 555294 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 555914 664634
rect 555294 628954 555914 664398
rect 555294 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 555914 628954
rect 555294 628634 555914 628718
rect 555294 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 555914 628634
rect 555294 592954 555914 628398
rect 555294 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 555914 592954
rect 555294 592634 555914 592718
rect 555294 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 555914 592634
rect 555294 556954 555914 592398
rect 555294 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 555914 556954
rect 555294 556634 555914 556718
rect 555294 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 555914 556634
rect 555294 520954 555914 556398
rect 555294 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 555914 520954
rect 555294 520634 555914 520718
rect 555294 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 555914 520634
rect 555294 484954 555914 520398
rect 555294 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 555914 484954
rect 555294 484634 555914 484718
rect 555294 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 555914 484634
rect 555294 448954 555914 484398
rect 555294 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 555914 448954
rect 555294 448634 555914 448718
rect 555294 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 555914 448634
rect 555294 412954 555914 448398
rect 555294 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 555914 412954
rect 555294 412634 555914 412718
rect 555294 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 555914 412634
rect 555294 376954 555914 412398
rect 555294 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 555914 376954
rect 555294 376634 555914 376718
rect 555294 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 555914 376634
rect 555294 340954 555914 376398
rect 555294 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 555914 340954
rect 555294 340634 555914 340718
rect 555294 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 555914 340634
rect 555294 304954 555914 340398
rect 555294 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 555914 304954
rect 555294 304634 555914 304718
rect 555294 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 555914 304634
rect 555294 268954 555914 304398
rect 555294 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 555914 268954
rect 555294 268634 555914 268718
rect 555294 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 555914 268634
rect 555294 232954 555914 268398
rect 555294 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 555914 232954
rect 555294 232634 555914 232718
rect 555294 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 555914 232634
rect 555294 196954 555914 232398
rect 555294 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 555914 196954
rect 555294 196634 555914 196718
rect 555294 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 555914 196634
rect 555294 160954 555914 196398
rect 555294 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 555914 160954
rect 555294 160634 555914 160718
rect 555294 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 555914 160634
rect 555294 124954 555914 160398
rect 555294 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 555914 124954
rect 555294 124634 555914 124718
rect 555294 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 555914 124634
rect 555294 88954 555914 124398
rect 555294 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 555914 88954
rect 555294 88634 555914 88718
rect 555294 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 555914 88634
rect 555294 52954 555914 88398
rect 555294 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 555914 52954
rect 555294 52634 555914 52718
rect 555294 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 555914 52634
rect 555294 16954 555914 52398
rect 555294 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 555914 16954
rect 555294 16634 555914 16718
rect 555294 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 555914 16634
rect 555294 -3226 555914 16398
rect 555294 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 555914 -3226
rect 555294 -3546 555914 -3462
rect 555294 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 555914 -3546
rect 555294 -7654 555914 -3782
rect 559794 708678 560414 711590
rect 559794 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 560414 708678
rect 559794 708358 560414 708442
rect 559794 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 560414 708358
rect 559794 669454 560414 708122
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -4186 560414 20898
rect 559794 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 560414 -4186
rect 559794 -4506 560414 -4422
rect 559794 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 560414 -4506
rect 559794 -7654 560414 -4742
rect 564294 709638 564914 711590
rect 564294 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 564914 709638
rect 564294 709318 564914 709402
rect 564294 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 564914 709318
rect 564294 673954 564914 709082
rect 564294 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 564914 673954
rect 564294 673634 564914 673718
rect 564294 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 564914 673634
rect 564294 637954 564914 673398
rect 564294 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 564914 637954
rect 564294 637634 564914 637718
rect 564294 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 564914 637634
rect 564294 601954 564914 637398
rect 564294 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 564914 601954
rect 564294 601634 564914 601718
rect 564294 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 564914 601634
rect 564294 565954 564914 601398
rect 564294 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 564914 565954
rect 564294 565634 564914 565718
rect 564294 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 564914 565634
rect 564294 529954 564914 565398
rect 564294 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 564914 529954
rect 564294 529634 564914 529718
rect 564294 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 564914 529634
rect 564294 493954 564914 529398
rect 564294 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 564914 493954
rect 564294 493634 564914 493718
rect 564294 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 564914 493634
rect 564294 457954 564914 493398
rect 564294 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 564914 457954
rect 564294 457634 564914 457718
rect 564294 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 564914 457634
rect 564294 421954 564914 457398
rect 564294 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 564914 421954
rect 564294 421634 564914 421718
rect 564294 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 564914 421634
rect 564294 385954 564914 421398
rect 564294 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 564914 385954
rect 564294 385634 564914 385718
rect 564294 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 564914 385634
rect 564294 349954 564914 385398
rect 564294 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 564914 349954
rect 564294 349634 564914 349718
rect 564294 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 564914 349634
rect 564294 313954 564914 349398
rect 564294 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 564914 313954
rect 564294 313634 564914 313718
rect 564294 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 564914 313634
rect 564294 277954 564914 313398
rect 564294 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 564914 277954
rect 564294 277634 564914 277718
rect 564294 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 564914 277634
rect 564294 241954 564914 277398
rect 564294 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 564914 241954
rect 564294 241634 564914 241718
rect 564294 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 564914 241634
rect 564294 205954 564914 241398
rect 564294 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 564914 205954
rect 564294 205634 564914 205718
rect 564294 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 564914 205634
rect 564294 169954 564914 205398
rect 564294 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 564914 169954
rect 564294 169634 564914 169718
rect 564294 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 564914 169634
rect 564294 133954 564914 169398
rect 564294 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 564914 133954
rect 564294 133634 564914 133718
rect 564294 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 564914 133634
rect 564294 97954 564914 133398
rect 564294 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 564914 97954
rect 564294 97634 564914 97718
rect 564294 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 564914 97634
rect 564294 61954 564914 97398
rect 564294 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 564914 61954
rect 564294 61634 564914 61718
rect 564294 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 564914 61634
rect 564294 25954 564914 61398
rect 564294 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 564914 25954
rect 564294 25634 564914 25718
rect 564294 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 564914 25634
rect 564294 -5146 564914 25398
rect 564294 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 564914 -5146
rect 564294 -5466 564914 -5382
rect 564294 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 564914 -5466
rect 564294 -7654 564914 -5702
rect 568794 710598 569414 711590
rect 568794 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 569414 710598
rect 568794 710278 569414 710362
rect 568794 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 569414 710278
rect 568794 678454 569414 710042
rect 568794 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 569414 678454
rect 568794 678134 569414 678218
rect 568794 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 569414 678134
rect 568794 642454 569414 677898
rect 568794 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 569414 642454
rect 568794 642134 569414 642218
rect 568794 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 569414 642134
rect 568794 606454 569414 641898
rect 568794 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 569414 606454
rect 568794 606134 569414 606218
rect 568794 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 569414 606134
rect 568794 570454 569414 605898
rect 568794 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 569414 570454
rect 568794 570134 569414 570218
rect 568794 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 569414 570134
rect 568794 534454 569414 569898
rect 568794 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 569414 534454
rect 568794 534134 569414 534218
rect 568794 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 569414 534134
rect 568794 498454 569414 533898
rect 568794 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 569414 498454
rect 568794 498134 569414 498218
rect 568794 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 569414 498134
rect 568794 462454 569414 497898
rect 568794 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 569414 462454
rect 568794 462134 569414 462218
rect 568794 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 569414 462134
rect 568794 426454 569414 461898
rect 568794 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 569414 426454
rect 568794 426134 569414 426218
rect 568794 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 569414 426134
rect 568794 390454 569414 425898
rect 568794 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 569414 390454
rect 568794 390134 569414 390218
rect 568794 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 569414 390134
rect 568794 354454 569414 389898
rect 568794 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 569414 354454
rect 568794 354134 569414 354218
rect 568794 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 569414 354134
rect 568794 318454 569414 353898
rect 568794 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 569414 318454
rect 568794 318134 569414 318218
rect 568794 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 569414 318134
rect 568794 282454 569414 317898
rect 568794 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 569414 282454
rect 568794 282134 569414 282218
rect 568794 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 569414 282134
rect 568794 246454 569414 281898
rect 568794 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 569414 246454
rect 568794 246134 569414 246218
rect 568794 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 569414 246134
rect 568794 210454 569414 245898
rect 568794 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 569414 210454
rect 568794 210134 569414 210218
rect 568794 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 569414 210134
rect 568794 174454 569414 209898
rect 568794 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 569414 174454
rect 568794 174134 569414 174218
rect 568794 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 569414 174134
rect 568794 138454 569414 173898
rect 568794 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 569414 138454
rect 568794 138134 569414 138218
rect 568794 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 569414 138134
rect 568794 102454 569414 137898
rect 568794 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 569414 102454
rect 568794 102134 569414 102218
rect 568794 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 569414 102134
rect 568794 66454 569414 101898
rect 568794 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 569414 66454
rect 568794 66134 569414 66218
rect 568794 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 569414 66134
rect 568794 30454 569414 65898
rect 568794 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 569414 30454
rect 568794 30134 569414 30218
rect 568794 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 569414 30134
rect 568794 -6106 569414 29898
rect 568794 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 569414 -6106
rect 568794 -6426 569414 -6342
rect 568794 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 569414 -6426
rect 568794 -7654 569414 -6662
rect 573294 711558 573914 711590
rect 573294 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 573914 711558
rect 573294 711238 573914 711322
rect 573294 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 573914 711238
rect 573294 682954 573914 711002
rect 573294 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 573914 682954
rect 573294 682634 573914 682718
rect 573294 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 573914 682634
rect 573294 646954 573914 682398
rect 573294 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 573914 646954
rect 573294 646634 573914 646718
rect 573294 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 573914 646634
rect 573294 610954 573914 646398
rect 573294 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 573914 610954
rect 573294 610634 573914 610718
rect 573294 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 573914 610634
rect 573294 574954 573914 610398
rect 573294 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 573914 574954
rect 573294 574634 573914 574718
rect 573294 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 573914 574634
rect 573294 538954 573914 574398
rect 573294 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 573914 538954
rect 573294 538634 573914 538718
rect 573294 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 573914 538634
rect 573294 502954 573914 538398
rect 573294 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 573914 502954
rect 573294 502634 573914 502718
rect 573294 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 573914 502634
rect 573294 466954 573914 502398
rect 573294 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 573914 466954
rect 573294 466634 573914 466718
rect 573294 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 573914 466634
rect 573294 430954 573914 466398
rect 573294 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 573914 430954
rect 573294 430634 573914 430718
rect 573294 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 573914 430634
rect 573294 394954 573914 430398
rect 573294 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 573914 394954
rect 573294 394634 573914 394718
rect 573294 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 573914 394634
rect 573294 358954 573914 394398
rect 573294 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 573914 358954
rect 573294 358634 573914 358718
rect 573294 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 573914 358634
rect 573294 322954 573914 358398
rect 573294 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 573914 322954
rect 573294 322634 573914 322718
rect 573294 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 573914 322634
rect 573294 286954 573914 322398
rect 573294 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 573914 286954
rect 573294 286634 573914 286718
rect 573294 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 573914 286634
rect 573294 250954 573914 286398
rect 573294 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 573914 250954
rect 573294 250634 573914 250718
rect 573294 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 573914 250634
rect 573294 214954 573914 250398
rect 573294 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 573914 214954
rect 573294 214634 573914 214718
rect 573294 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 573914 214634
rect 573294 178954 573914 214398
rect 573294 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 573914 178954
rect 573294 178634 573914 178718
rect 573294 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 573914 178634
rect 573294 142954 573914 178398
rect 573294 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 573914 142954
rect 573294 142634 573914 142718
rect 573294 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 573914 142634
rect 573294 106954 573914 142398
rect 573294 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 573914 106954
rect 573294 106634 573914 106718
rect 573294 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 573914 106634
rect 573294 70954 573914 106398
rect 573294 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 573914 70954
rect 573294 70634 573914 70718
rect 573294 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 573914 70634
rect 573294 34954 573914 70398
rect 573294 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 573914 34954
rect 573294 34634 573914 34718
rect 573294 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 573914 34634
rect 573294 -7066 573914 34398
rect 573294 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 573914 -7066
rect 573294 -7386 573914 -7302
rect 573294 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 573914 -7386
rect 573294 -7654 573914 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect 582294 691954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 582914 691954
rect 582294 691634 582914 691718
rect 582294 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 582914 691634
rect 582294 655954 582914 691398
rect 582294 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 582914 655954
rect 582294 655634 582914 655718
rect 582294 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 582914 655634
rect 582294 619954 582914 655398
rect 582294 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 582914 619954
rect 582294 619634 582914 619718
rect 582294 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 582914 619634
rect 582294 583954 582914 619398
rect 582294 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 582914 583954
rect 582294 583634 582914 583718
rect 582294 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 582914 583634
rect 582294 547954 582914 583398
rect 582294 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 582914 547954
rect 582294 547634 582914 547718
rect 582294 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 582914 547634
rect 582294 511954 582914 547398
rect 582294 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 582914 511954
rect 582294 511634 582914 511718
rect 582294 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 582914 511634
rect 582294 475954 582914 511398
rect 582294 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 582914 475954
rect 582294 475634 582914 475718
rect 582294 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 582914 475634
rect 582294 439954 582914 475398
rect 582294 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 582914 439954
rect 582294 439634 582914 439718
rect 582294 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 582914 439634
rect 582294 403954 582914 439398
rect 582294 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 582914 403954
rect 582294 403634 582914 403718
rect 582294 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 582914 403634
rect 582294 367954 582914 403398
rect 582294 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 582914 367954
rect 582294 367634 582914 367718
rect 582294 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 582914 367634
rect 582294 331954 582914 367398
rect 582294 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 582914 331954
rect 582294 331634 582914 331718
rect 582294 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 582914 331634
rect 582294 295954 582914 331398
rect 582294 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 582914 295954
rect 582294 295634 582914 295718
rect 582294 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 582914 295634
rect 582294 259954 582914 295398
rect 582294 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 582914 259954
rect 582294 259634 582914 259718
rect 582294 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 582914 259634
rect 582294 223954 582914 259398
rect 582294 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 582914 223954
rect 582294 223634 582914 223718
rect 582294 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 582914 223634
rect 582294 187954 582914 223398
rect 582294 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 582914 187954
rect 582294 187634 582914 187718
rect 582294 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 582914 187634
rect 582294 151954 582914 187398
rect 582294 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 582914 151954
rect 582294 151634 582914 151718
rect 582294 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 582914 151634
rect 582294 115954 582914 151398
rect 582294 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 582914 115954
rect 582294 115634 582914 115718
rect 582294 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 582914 115634
rect 582294 79954 582914 115398
rect 582294 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 582914 79954
rect 582294 79634 582914 79718
rect 582294 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 582914 79634
rect 582294 43954 582914 79398
rect 582294 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 582914 43954
rect 582294 43634 582914 43718
rect 582294 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 582914 43634
rect 582294 7954 582914 43398
rect 582294 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 582914 7954
rect 582294 7634 582914 7718
rect 582294 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 582914 7634
rect 582294 -1306 582914 7398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691954 586890 705242
rect 586270 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 586890 691954
rect 586270 691634 586890 691718
rect 586270 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 586890 691634
rect 586270 655954 586890 691398
rect 586270 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 586890 655954
rect 586270 655634 586890 655718
rect 586270 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 586890 655634
rect 586270 619954 586890 655398
rect 586270 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 586890 619954
rect 586270 619634 586890 619718
rect 586270 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 586890 619634
rect 586270 583954 586890 619398
rect 586270 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 586890 583954
rect 586270 583634 586890 583718
rect 586270 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 586890 583634
rect 586270 547954 586890 583398
rect 586270 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 586890 547954
rect 586270 547634 586890 547718
rect 586270 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 586890 547634
rect 586270 511954 586890 547398
rect 586270 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 586890 511954
rect 586270 511634 586890 511718
rect 586270 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 586890 511634
rect 586270 475954 586890 511398
rect 586270 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 586890 475954
rect 586270 475634 586890 475718
rect 586270 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 586890 475634
rect 586270 439954 586890 475398
rect 586270 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 586890 439954
rect 586270 439634 586890 439718
rect 586270 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 586890 439634
rect 586270 403954 586890 439398
rect 586270 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 586890 403954
rect 586270 403634 586890 403718
rect 586270 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 586890 403634
rect 586270 367954 586890 403398
rect 586270 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 586890 367954
rect 586270 367634 586890 367718
rect 586270 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 586890 367634
rect 586270 331954 586890 367398
rect 586270 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 586890 331954
rect 586270 331634 586890 331718
rect 586270 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 586890 331634
rect 586270 295954 586890 331398
rect 586270 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 586890 295954
rect 586270 295634 586890 295718
rect 586270 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 586890 295634
rect 586270 259954 586890 295398
rect 586270 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 586890 259954
rect 586270 259634 586890 259718
rect 586270 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 586890 259634
rect 586270 223954 586890 259398
rect 586270 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 586890 223954
rect 586270 223634 586890 223718
rect 586270 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 586890 223634
rect 586270 187954 586890 223398
rect 586270 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 586890 187954
rect 586270 187634 586890 187718
rect 586270 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 586890 187634
rect 586270 151954 586890 187398
rect 586270 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 586890 151954
rect 586270 151634 586890 151718
rect 586270 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 586890 151634
rect 586270 115954 586890 151398
rect 586270 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 586890 115954
rect 586270 115634 586890 115718
rect 586270 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 586890 115634
rect 586270 79954 586890 115398
rect 586270 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 586890 79954
rect 586270 79634 586890 79718
rect 586270 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 586890 79634
rect 586270 43954 586890 79398
rect 586270 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 586890 43954
rect 586270 43634 586890 43718
rect 586270 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 586890 43634
rect 586270 7954 586890 43398
rect 586270 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 586890 7954
rect 586270 7634 586890 7718
rect 586270 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 586890 7634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 7398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 696454 587850 706202
rect 587230 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 587850 696454
rect 587230 696134 587850 696218
rect 587230 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 587850 696134
rect 587230 660454 587850 695898
rect 587230 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 587850 660454
rect 587230 660134 587850 660218
rect 587230 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 587850 660134
rect 587230 624454 587850 659898
rect 587230 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 587850 624454
rect 587230 624134 587850 624218
rect 587230 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 587850 624134
rect 587230 588454 587850 623898
rect 587230 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 587850 588454
rect 587230 588134 587850 588218
rect 587230 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 587850 588134
rect 587230 552454 587850 587898
rect 587230 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 587850 552454
rect 587230 552134 587850 552218
rect 587230 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 587850 552134
rect 587230 516454 587850 551898
rect 587230 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 587850 516454
rect 587230 516134 587850 516218
rect 587230 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 587850 516134
rect 587230 480454 587850 515898
rect 587230 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 587850 480454
rect 587230 480134 587850 480218
rect 587230 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 587850 480134
rect 587230 444454 587850 479898
rect 587230 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 587850 444454
rect 587230 444134 587850 444218
rect 587230 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 587850 444134
rect 587230 408454 587850 443898
rect 587230 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 587850 408454
rect 587230 408134 587850 408218
rect 587230 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 587850 408134
rect 587230 372454 587850 407898
rect 587230 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 587850 372454
rect 587230 372134 587850 372218
rect 587230 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 587850 372134
rect 587230 336454 587850 371898
rect 587230 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 587850 336454
rect 587230 336134 587850 336218
rect 587230 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 587850 336134
rect 587230 300454 587850 335898
rect 587230 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 587850 300454
rect 587230 300134 587850 300218
rect 587230 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 587850 300134
rect 587230 264454 587850 299898
rect 587230 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 587850 264454
rect 587230 264134 587850 264218
rect 587230 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 587850 264134
rect 587230 228454 587850 263898
rect 587230 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 587850 228454
rect 587230 228134 587850 228218
rect 587230 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 587850 228134
rect 587230 192454 587850 227898
rect 587230 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 587850 192454
rect 587230 192134 587850 192218
rect 587230 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 587850 192134
rect 587230 156454 587850 191898
rect 587230 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 587850 156454
rect 587230 156134 587850 156218
rect 587230 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 587850 156134
rect 587230 120454 587850 155898
rect 587230 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 587850 120454
rect 587230 120134 587850 120218
rect 587230 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 587850 120134
rect 587230 84454 587850 119898
rect 587230 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 587850 84454
rect 587230 84134 587850 84218
rect 587230 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 587850 84134
rect 587230 48454 587850 83898
rect 587230 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 587850 48454
rect 587230 48134 587850 48218
rect 587230 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 587850 48134
rect 587230 12454 587850 47898
rect 587230 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 587850 12454
rect 587230 12134 587850 12218
rect 587230 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 587850 12134
rect 587230 -2266 587850 11898
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 700954 588810 707162
rect 588190 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 588810 700954
rect 588190 700634 588810 700718
rect 588190 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 588810 700634
rect 588190 664954 588810 700398
rect 588190 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 588810 664954
rect 588190 664634 588810 664718
rect 588190 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 588810 664634
rect 588190 628954 588810 664398
rect 588190 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 588810 628954
rect 588190 628634 588810 628718
rect 588190 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 588810 628634
rect 588190 592954 588810 628398
rect 588190 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 588810 592954
rect 588190 592634 588810 592718
rect 588190 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 588810 592634
rect 588190 556954 588810 592398
rect 588190 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 588810 556954
rect 588190 556634 588810 556718
rect 588190 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 588810 556634
rect 588190 520954 588810 556398
rect 588190 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 588810 520954
rect 588190 520634 588810 520718
rect 588190 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 588810 520634
rect 588190 484954 588810 520398
rect 588190 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 588810 484954
rect 588190 484634 588810 484718
rect 588190 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 588810 484634
rect 588190 448954 588810 484398
rect 588190 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 588810 448954
rect 588190 448634 588810 448718
rect 588190 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 588810 448634
rect 588190 412954 588810 448398
rect 588190 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 588810 412954
rect 588190 412634 588810 412718
rect 588190 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 588810 412634
rect 588190 376954 588810 412398
rect 588190 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 588810 376954
rect 588190 376634 588810 376718
rect 588190 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 588810 376634
rect 588190 340954 588810 376398
rect 588190 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 588810 340954
rect 588190 340634 588810 340718
rect 588190 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 588810 340634
rect 588190 304954 588810 340398
rect 588190 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 588810 304954
rect 588190 304634 588810 304718
rect 588190 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 588810 304634
rect 588190 268954 588810 304398
rect 588190 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 588810 268954
rect 588190 268634 588810 268718
rect 588190 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 588810 268634
rect 588190 232954 588810 268398
rect 588190 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 588810 232954
rect 588190 232634 588810 232718
rect 588190 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 588810 232634
rect 588190 196954 588810 232398
rect 588190 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 588810 196954
rect 588190 196634 588810 196718
rect 588190 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 588810 196634
rect 588190 160954 588810 196398
rect 588190 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 588810 160954
rect 588190 160634 588810 160718
rect 588190 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 588810 160634
rect 588190 124954 588810 160398
rect 588190 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 588810 124954
rect 588190 124634 588810 124718
rect 588190 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 588810 124634
rect 588190 88954 588810 124398
rect 588190 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 588810 88954
rect 588190 88634 588810 88718
rect 588190 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 588810 88634
rect 588190 52954 588810 88398
rect 588190 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 588810 52954
rect 588190 52634 588810 52718
rect 588190 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 588810 52634
rect 588190 16954 588810 52398
rect 588190 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 588810 16954
rect 588190 16634 588810 16718
rect 588190 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 588810 16634
rect 588190 -3226 588810 16398
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 669454 589770 708122
rect 589150 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 589770 669454
rect 589150 669134 589770 669218
rect 589150 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 589770 669134
rect 589150 633454 589770 668898
rect 589150 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 589770 633454
rect 589150 633134 589770 633218
rect 589150 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 589770 633134
rect 589150 597454 589770 632898
rect 589150 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 589770 597454
rect 589150 597134 589770 597218
rect 589150 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 589770 597134
rect 589150 561454 589770 596898
rect 589150 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 589770 561454
rect 589150 561134 589770 561218
rect 589150 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 589770 561134
rect 589150 525454 589770 560898
rect 589150 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 589770 525454
rect 589150 525134 589770 525218
rect 589150 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 589770 525134
rect 589150 489454 589770 524898
rect 589150 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 589770 489454
rect 589150 489134 589770 489218
rect 589150 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 589770 489134
rect 589150 453454 589770 488898
rect 589150 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 589770 453454
rect 589150 453134 589770 453218
rect 589150 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 589770 453134
rect 589150 417454 589770 452898
rect 589150 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 589770 417454
rect 589150 417134 589770 417218
rect 589150 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 589770 417134
rect 589150 381454 589770 416898
rect 589150 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 589770 381454
rect 589150 381134 589770 381218
rect 589150 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 589770 381134
rect 589150 345454 589770 380898
rect 589150 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 589770 345454
rect 589150 345134 589770 345218
rect 589150 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 589770 345134
rect 589150 309454 589770 344898
rect 589150 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 589770 309454
rect 589150 309134 589770 309218
rect 589150 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 589770 309134
rect 589150 273454 589770 308898
rect 589150 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 589770 273454
rect 589150 273134 589770 273218
rect 589150 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 589770 273134
rect 589150 237454 589770 272898
rect 589150 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 589770 237454
rect 589150 237134 589770 237218
rect 589150 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 589770 237134
rect 589150 201454 589770 236898
rect 589150 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 589770 201454
rect 589150 201134 589770 201218
rect 589150 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 589770 201134
rect 589150 165454 589770 200898
rect 589150 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 589770 165454
rect 589150 165134 589770 165218
rect 589150 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 589770 165134
rect 589150 129454 589770 164898
rect 589150 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 589770 129454
rect 589150 129134 589770 129218
rect 589150 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 589770 129134
rect 589150 93454 589770 128898
rect 589150 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 589770 93454
rect 589150 93134 589770 93218
rect 589150 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 589770 93134
rect 589150 57454 589770 92898
rect 589150 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 589770 57454
rect 589150 57134 589770 57218
rect 589150 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 589770 57134
rect 589150 21454 589770 56898
rect 589150 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 589770 21454
rect 589150 21134 589770 21218
rect 589150 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 589770 21134
rect 589150 -4186 589770 20898
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 673954 590730 709082
rect 590110 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 590730 673954
rect 590110 673634 590730 673718
rect 590110 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 590730 673634
rect 590110 637954 590730 673398
rect 590110 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 590730 637954
rect 590110 637634 590730 637718
rect 590110 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 590730 637634
rect 590110 601954 590730 637398
rect 590110 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 590730 601954
rect 590110 601634 590730 601718
rect 590110 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 590730 601634
rect 590110 565954 590730 601398
rect 590110 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 590730 565954
rect 590110 565634 590730 565718
rect 590110 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 590730 565634
rect 590110 529954 590730 565398
rect 590110 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 590730 529954
rect 590110 529634 590730 529718
rect 590110 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 590730 529634
rect 590110 493954 590730 529398
rect 590110 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 590730 493954
rect 590110 493634 590730 493718
rect 590110 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 590730 493634
rect 590110 457954 590730 493398
rect 590110 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 590730 457954
rect 590110 457634 590730 457718
rect 590110 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 590730 457634
rect 590110 421954 590730 457398
rect 590110 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 590730 421954
rect 590110 421634 590730 421718
rect 590110 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 590730 421634
rect 590110 385954 590730 421398
rect 590110 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 590730 385954
rect 590110 385634 590730 385718
rect 590110 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 590730 385634
rect 590110 349954 590730 385398
rect 590110 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 590730 349954
rect 590110 349634 590730 349718
rect 590110 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 590730 349634
rect 590110 313954 590730 349398
rect 590110 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 590730 313954
rect 590110 313634 590730 313718
rect 590110 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 590730 313634
rect 590110 277954 590730 313398
rect 590110 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 590730 277954
rect 590110 277634 590730 277718
rect 590110 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 590730 277634
rect 590110 241954 590730 277398
rect 590110 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 590730 241954
rect 590110 241634 590730 241718
rect 590110 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 590730 241634
rect 590110 205954 590730 241398
rect 590110 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 590730 205954
rect 590110 205634 590730 205718
rect 590110 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 590730 205634
rect 590110 169954 590730 205398
rect 590110 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 590730 169954
rect 590110 169634 590730 169718
rect 590110 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 590730 169634
rect 590110 133954 590730 169398
rect 590110 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 590730 133954
rect 590110 133634 590730 133718
rect 590110 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 590730 133634
rect 590110 97954 590730 133398
rect 590110 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 590730 97954
rect 590110 97634 590730 97718
rect 590110 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 590730 97634
rect 590110 61954 590730 97398
rect 590110 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 590730 61954
rect 590110 61634 590730 61718
rect 590110 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 590730 61634
rect 590110 25954 590730 61398
rect 590110 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 590730 25954
rect 590110 25634 590730 25718
rect 590110 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 590730 25634
rect 590110 -5146 590730 25398
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 678454 591690 710042
rect 591070 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 591690 678454
rect 591070 678134 591690 678218
rect 591070 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 591690 678134
rect 591070 642454 591690 677898
rect 591070 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 591690 642454
rect 591070 642134 591690 642218
rect 591070 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 591690 642134
rect 591070 606454 591690 641898
rect 591070 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 591690 606454
rect 591070 606134 591690 606218
rect 591070 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 591690 606134
rect 591070 570454 591690 605898
rect 591070 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 591690 570454
rect 591070 570134 591690 570218
rect 591070 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 591690 570134
rect 591070 534454 591690 569898
rect 591070 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 591690 534454
rect 591070 534134 591690 534218
rect 591070 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 591690 534134
rect 591070 498454 591690 533898
rect 591070 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 591690 498454
rect 591070 498134 591690 498218
rect 591070 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 591690 498134
rect 591070 462454 591690 497898
rect 591070 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 591690 462454
rect 591070 462134 591690 462218
rect 591070 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 591690 462134
rect 591070 426454 591690 461898
rect 591070 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 591690 426454
rect 591070 426134 591690 426218
rect 591070 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 591690 426134
rect 591070 390454 591690 425898
rect 591070 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 591690 390454
rect 591070 390134 591690 390218
rect 591070 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 591690 390134
rect 591070 354454 591690 389898
rect 591070 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 591690 354454
rect 591070 354134 591690 354218
rect 591070 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 591690 354134
rect 591070 318454 591690 353898
rect 591070 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 591690 318454
rect 591070 318134 591690 318218
rect 591070 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 591690 318134
rect 591070 282454 591690 317898
rect 591070 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 591690 282454
rect 591070 282134 591690 282218
rect 591070 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 591690 282134
rect 591070 246454 591690 281898
rect 591070 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 591690 246454
rect 591070 246134 591690 246218
rect 591070 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 591690 246134
rect 591070 210454 591690 245898
rect 591070 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 591690 210454
rect 591070 210134 591690 210218
rect 591070 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 591690 210134
rect 591070 174454 591690 209898
rect 591070 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 591690 174454
rect 591070 174134 591690 174218
rect 591070 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 591690 174134
rect 591070 138454 591690 173898
rect 591070 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 591690 138454
rect 591070 138134 591690 138218
rect 591070 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 591690 138134
rect 591070 102454 591690 137898
rect 591070 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 591690 102454
rect 591070 102134 591690 102218
rect 591070 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 591690 102134
rect 591070 66454 591690 101898
rect 591070 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 591690 66454
rect 591070 66134 591690 66218
rect 591070 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 591690 66134
rect 591070 30454 591690 65898
rect 591070 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 591690 30454
rect 591070 30134 591690 30218
rect 591070 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 591690 30134
rect 591070 -6106 591690 29898
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 682954 592650 711002
rect 592030 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect 592030 682634 592650 682718
rect 592030 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect 592030 646954 592650 682398
rect 592030 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect 592030 646634 592650 646718
rect 592030 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect 592030 610954 592650 646398
rect 592030 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect 592030 610634 592650 610718
rect 592030 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect 592030 574954 592650 610398
rect 592030 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect 592030 574634 592650 574718
rect 592030 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect 592030 538954 592650 574398
rect 592030 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect 592030 538634 592650 538718
rect 592030 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect 592030 502954 592650 538398
rect 592030 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect 592030 502634 592650 502718
rect 592030 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect 592030 466954 592650 502398
rect 592030 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect 592030 466634 592650 466718
rect 592030 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect 592030 430954 592650 466398
rect 592030 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect 592030 430634 592650 430718
rect 592030 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect 592030 394954 592650 430398
rect 592030 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect 592030 394634 592650 394718
rect 592030 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect 592030 358954 592650 394398
rect 592030 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect 592030 358634 592650 358718
rect 592030 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect 592030 322954 592650 358398
rect 592030 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect 592030 322634 592650 322718
rect 592030 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect 592030 286954 592650 322398
rect 592030 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect 592030 286634 592650 286718
rect 592030 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect 592030 250954 592650 286398
rect 592030 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect 592030 250634 592650 250718
rect 592030 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect 592030 214954 592650 250398
rect 592030 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect 592030 214634 592650 214718
rect 592030 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect 592030 178954 592650 214398
rect 592030 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect 592030 178634 592650 178718
rect 592030 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect 592030 142954 592650 178398
rect 592030 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect 592030 142634 592650 142718
rect 592030 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect 592030 106954 592650 142398
rect 592030 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect 592030 106634 592650 106718
rect 592030 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect 592030 70954 592650 106398
rect 592030 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect 592030 70634 592650 70718
rect 592030 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect 592030 34954 592650 70398
rect 592030 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect 592030 34634 592650 34718
rect 592030 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect 592030 -7066 592650 34398
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 682718 -8458 682954
rect -8374 682718 -8138 682954
rect -8694 682398 -8458 682634
rect -8374 682398 -8138 682634
rect -8694 646718 -8458 646954
rect -8374 646718 -8138 646954
rect -8694 646398 -8458 646634
rect -8374 646398 -8138 646634
rect -8694 610718 -8458 610954
rect -8374 610718 -8138 610954
rect -8694 610398 -8458 610634
rect -8374 610398 -8138 610634
rect -8694 574718 -8458 574954
rect -8374 574718 -8138 574954
rect -8694 574398 -8458 574634
rect -8374 574398 -8138 574634
rect -8694 538718 -8458 538954
rect -8374 538718 -8138 538954
rect -8694 538398 -8458 538634
rect -8374 538398 -8138 538634
rect -8694 502718 -8458 502954
rect -8374 502718 -8138 502954
rect -8694 502398 -8458 502634
rect -8374 502398 -8138 502634
rect -8694 466718 -8458 466954
rect -8374 466718 -8138 466954
rect -8694 466398 -8458 466634
rect -8374 466398 -8138 466634
rect -8694 430718 -8458 430954
rect -8374 430718 -8138 430954
rect -8694 430398 -8458 430634
rect -8374 430398 -8138 430634
rect -8694 394718 -8458 394954
rect -8374 394718 -8138 394954
rect -8694 394398 -8458 394634
rect -8374 394398 -8138 394634
rect -8694 358718 -8458 358954
rect -8374 358718 -8138 358954
rect -8694 358398 -8458 358634
rect -8374 358398 -8138 358634
rect -8694 322718 -8458 322954
rect -8374 322718 -8138 322954
rect -8694 322398 -8458 322634
rect -8374 322398 -8138 322634
rect -8694 286718 -8458 286954
rect -8374 286718 -8138 286954
rect -8694 286398 -8458 286634
rect -8374 286398 -8138 286634
rect -8694 250718 -8458 250954
rect -8374 250718 -8138 250954
rect -8694 250398 -8458 250634
rect -8374 250398 -8138 250634
rect -8694 214718 -8458 214954
rect -8374 214718 -8138 214954
rect -8694 214398 -8458 214634
rect -8374 214398 -8138 214634
rect -8694 178718 -8458 178954
rect -8374 178718 -8138 178954
rect -8694 178398 -8458 178634
rect -8374 178398 -8138 178634
rect -8694 142718 -8458 142954
rect -8374 142718 -8138 142954
rect -8694 142398 -8458 142634
rect -8374 142398 -8138 142634
rect -8694 106718 -8458 106954
rect -8374 106718 -8138 106954
rect -8694 106398 -8458 106634
rect -8374 106398 -8138 106634
rect -8694 70718 -8458 70954
rect -8374 70718 -8138 70954
rect -8694 70398 -8458 70634
rect -8374 70398 -8138 70634
rect -8694 34718 -8458 34954
rect -8374 34718 -8138 34954
rect -8694 34398 -8458 34634
rect -8374 34398 -8138 34634
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 678218 -7498 678454
rect -7414 678218 -7178 678454
rect -7734 677898 -7498 678134
rect -7414 677898 -7178 678134
rect -7734 642218 -7498 642454
rect -7414 642218 -7178 642454
rect -7734 641898 -7498 642134
rect -7414 641898 -7178 642134
rect -7734 606218 -7498 606454
rect -7414 606218 -7178 606454
rect -7734 605898 -7498 606134
rect -7414 605898 -7178 606134
rect -7734 570218 -7498 570454
rect -7414 570218 -7178 570454
rect -7734 569898 -7498 570134
rect -7414 569898 -7178 570134
rect -7734 534218 -7498 534454
rect -7414 534218 -7178 534454
rect -7734 533898 -7498 534134
rect -7414 533898 -7178 534134
rect -7734 498218 -7498 498454
rect -7414 498218 -7178 498454
rect -7734 497898 -7498 498134
rect -7414 497898 -7178 498134
rect -7734 462218 -7498 462454
rect -7414 462218 -7178 462454
rect -7734 461898 -7498 462134
rect -7414 461898 -7178 462134
rect -7734 426218 -7498 426454
rect -7414 426218 -7178 426454
rect -7734 425898 -7498 426134
rect -7414 425898 -7178 426134
rect -7734 390218 -7498 390454
rect -7414 390218 -7178 390454
rect -7734 389898 -7498 390134
rect -7414 389898 -7178 390134
rect -7734 354218 -7498 354454
rect -7414 354218 -7178 354454
rect -7734 353898 -7498 354134
rect -7414 353898 -7178 354134
rect -7734 318218 -7498 318454
rect -7414 318218 -7178 318454
rect -7734 317898 -7498 318134
rect -7414 317898 -7178 318134
rect -7734 282218 -7498 282454
rect -7414 282218 -7178 282454
rect -7734 281898 -7498 282134
rect -7414 281898 -7178 282134
rect -7734 246218 -7498 246454
rect -7414 246218 -7178 246454
rect -7734 245898 -7498 246134
rect -7414 245898 -7178 246134
rect -7734 210218 -7498 210454
rect -7414 210218 -7178 210454
rect -7734 209898 -7498 210134
rect -7414 209898 -7178 210134
rect -7734 174218 -7498 174454
rect -7414 174218 -7178 174454
rect -7734 173898 -7498 174134
rect -7414 173898 -7178 174134
rect -7734 138218 -7498 138454
rect -7414 138218 -7178 138454
rect -7734 137898 -7498 138134
rect -7414 137898 -7178 138134
rect -7734 102218 -7498 102454
rect -7414 102218 -7178 102454
rect -7734 101898 -7498 102134
rect -7414 101898 -7178 102134
rect -7734 66218 -7498 66454
rect -7414 66218 -7178 66454
rect -7734 65898 -7498 66134
rect -7414 65898 -7178 66134
rect -7734 30218 -7498 30454
rect -7414 30218 -7178 30454
rect -7734 29898 -7498 30134
rect -7414 29898 -7178 30134
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 673718 -6538 673954
rect -6454 673718 -6218 673954
rect -6774 673398 -6538 673634
rect -6454 673398 -6218 673634
rect -6774 637718 -6538 637954
rect -6454 637718 -6218 637954
rect -6774 637398 -6538 637634
rect -6454 637398 -6218 637634
rect -6774 601718 -6538 601954
rect -6454 601718 -6218 601954
rect -6774 601398 -6538 601634
rect -6454 601398 -6218 601634
rect -6774 565718 -6538 565954
rect -6454 565718 -6218 565954
rect -6774 565398 -6538 565634
rect -6454 565398 -6218 565634
rect -6774 529718 -6538 529954
rect -6454 529718 -6218 529954
rect -6774 529398 -6538 529634
rect -6454 529398 -6218 529634
rect -6774 493718 -6538 493954
rect -6454 493718 -6218 493954
rect -6774 493398 -6538 493634
rect -6454 493398 -6218 493634
rect -6774 457718 -6538 457954
rect -6454 457718 -6218 457954
rect -6774 457398 -6538 457634
rect -6454 457398 -6218 457634
rect -6774 421718 -6538 421954
rect -6454 421718 -6218 421954
rect -6774 421398 -6538 421634
rect -6454 421398 -6218 421634
rect -6774 385718 -6538 385954
rect -6454 385718 -6218 385954
rect -6774 385398 -6538 385634
rect -6454 385398 -6218 385634
rect -6774 349718 -6538 349954
rect -6454 349718 -6218 349954
rect -6774 349398 -6538 349634
rect -6454 349398 -6218 349634
rect -6774 313718 -6538 313954
rect -6454 313718 -6218 313954
rect -6774 313398 -6538 313634
rect -6454 313398 -6218 313634
rect -6774 277718 -6538 277954
rect -6454 277718 -6218 277954
rect -6774 277398 -6538 277634
rect -6454 277398 -6218 277634
rect -6774 241718 -6538 241954
rect -6454 241718 -6218 241954
rect -6774 241398 -6538 241634
rect -6454 241398 -6218 241634
rect -6774 205718 -6538 205954
rect -6454 205718 -6218 205954
rect -6774 205398 -6538 205634
rect -6454 205398 -6218 205634
rect -6774 169718 -6538 169954
rect -6454 169718 -6218 169954
rect -6774 169398 -6538 169634
rect -6454 169398 -6218 169634
rect -6774 133718 -6538 133954
rect -6454 133718 -6218 133954
rect -6774 133398 -6538 133634
rect -6454 133398 -6218 133634
rect -6774 97718 -6538 97954
rect -6454 97718 -6218 97954
rect -6774 97398 -6538 97634
rect -6454 97398 -6218 97634
rect -6774 61718 -6538 61954
rect -6454 61718 -6218 61954
rect -6774 61398 -6538 61634
rect -6454 61398 -6218 61634
rect -6774 25718 -6538 25954
rect -6454 25718 -6218 25954
rect -6774 25398 -6538 25634
rect -6454 25398 -6218 25634
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 669218 -5578 669454
rect -5494 669218 -5258 669454
rect -5814 668898 -5578 669134
rect -5494 668898 -5258 669134
rect -5814 633218 -5578 633454
rect -5494 633218 -5258 633454
rect -5814 632898 -5578 633134
rect -5494 632898 -5258 633134
rect -5814 597218 -5578 597454
rect -5494 597218 -5258 597454
rect -5814 596898 -5578 597134
rect -5494 596898 -5258 597134
rect -5814 561218 -5578 561454
rect -5494 561218 -5258 561454
rect -5814 560898 -5578 561134
rect -5494 560898 -5258 561134
rect -5814 525218 -5578 525454
rect -5494 525218 -5258 525454
rect -5814 524898 -5578 525134
rect -5494 524898 -5258 525134
rect -5814 489218 -5578 489454
rect -5494 489218 -5258 489454
rect -5814 488898 -5578 489134
rect -5494 488898 -5258 489134
rect -5814 453218 -5578 453454
rect -5494 453218 -5258 453454
rect -5814 452898 -5578 453134
rect -5494 452898 -5258 453134
rect -5814 417218 -5578 417454
rect -5494 417218 -5258 417454
rect -5814 416898 -5578 417134
rect -5494 416898 -5258 417134
rect -5814 381218 -5578 381454
rect -5494 381218 -5258 381454
rect -5814 380898 -5578 381134
rect -5494 380898 -5258 381134
rect -5814 345218 -5578 345454
rect -5494 345218 -5258 345454
rect -5814 344898 -5578 345134
rect -5494 344898 -5258 345134
rect -5814 309218 -5578 309454
rect -5494 309218 -5258 309454
rect -5814 308898 -5578 309134
rect -5494 308898 -5258 309134
rect -5814 273218 -5578 273454
rect -5494 273218 -5258 273454
rect -5814 272898 -5578 273134
rect -5494 272898 -5258 273134
rect -5814 237218 -5578 237454
rect -5494 237218 -5258 237454
rect -5814 236898 -5578 237134
rect -5494 236898 -5258 237134
rect -5814 201218 -5578 201454
rect -5494 201218 -5258 201454
rect -5814 200898 -5578 201134
rect -5494 200898 -5258 201134
rect -5814 165218 -5578 165454
rect -5494 165218 -5258 165454
rect -5814 164898 -5578 165134
rect -5494 164898 -5258 165134
rect -5814 129218 -5578 129454
rect -5494 129218 -5258 129454
rect -5814 128898 -5578 129134
rect -5494 128898 -5258 129134
rect -5814 93218 -5578 93454
rect -5494 93218 -5258 93454
rect -5814 92898 -5578 93134
rect -5494 92898 -5258 93134
rect -5814 57218 -5578 57454
rect -5494 57218 -5258 57454
rect -5814 56898 -5578 57134
rect -5494 56898 -5258 57134
rect -5814 21218 -5578 21454
rect -5494 21218 -5258 21454
rect -5814 20898 -5578 21134
rect -5494 20898 -5258 21134
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 700718 -4618 700954
rect -4534 700718 -4298 700954
rect -4854 700398 -4618 700634
rect -4534 700398 -4298 700634
rect -4854 664718 -4618 664954
rect -4534 664718 -4298 664954
rect -4854 664398 -4618 664634
rect -4534 664398 -4298 664634
rect -4854 628718 -4618 628954
rect -4534 628718 -4298 628954
rect -4854 628398 -4618 628634
rect -4534 628398 -4298 628634
rect -4854 592718 -4618 592954
rect -4534 592718 -4298 592954
rect -4854 592398 -4618 592634
rect -4534 592398 -4298 592634
rect -4854 556718 -4618 556954
rect -4534 556718 -4298 556954
rect -4854 556398 -4618 556634
rect -4534 556398 -4298 556634
rect -4854 520718 -4618 520954
rect -4534 520718 -4298 520954
rect -4854 520398 -4618 520634
rect -4534 520398 -4298 520634
rect -4854 484718 -4618 484954
rect -4534 484718 -4298 484954
rect -4854 484398 -4618 484634
rect -4534 484398 -4298 484634
rect -4854 448718 -4618 448954
rect -4534 448718 -4298 448954
rect -4854 448398 -4618 448634
rect -4534 448398 -4298 448634
rect -4854 412718 -4618 412954
rect -4534 412718 -4298 412954
rect -4854 412398 -4618 412634
rect -4534 412398 -4298 412634
rect -4854 376718 -4618 376954
rect -4534 376718 -4298 376954
rect -4854 376398 -4618 376634
rect -4534 376398 -4298 376634
rect -4854 340718 -4618 340954
rect -4534 340718 -4298 340954
rect -4854 340398 -4618 340634
rect -4534 340398 -4298 340634
rect -4854 304718 -4618 304954
rect -4534 304718 -4298 304954
rect -4854 304398 -4618 304634
rect -4534 304398 -4298 304634
rect -4854 268718 -4618 268954
rect -4534 268718 -4298 268954
rect -4854 268398 -4618 268634
rect -4534 268398 -4298 268634
rect -4854 232718 -4618 232954
rect -4534 232718 -4298 232954
rect -4854 232398 -4618 232634
rect -4534 232398 -4298 232634
rect -4854 196718 -4618 196954
rect -4534 196718 -4298 196954
rect -4854 196398 -4618 196634
rect -4534 196398 -4298 196634
rect -4854 160718 -4618 160954
rect -4534 160718 -4298 160954
rect -4854 160398 -4618 160634
rect -4534 160398 -4298 160634
rect -4854 124718 -4618 124954
rect -4534 124718 -4298 124954
rect -4854 124398 -4618 124634
rect -4534 124398 -4298 124634
rect -4854 88718 -4618 88954
rect -4534 88718 -4298 88954
rect -4854 88398 -4618 88634
rect -4534 88398 -4298 88634
rect -4854 52718 -4618 52954
rect -4534 52718 -4298 52954
rect -4854 52398 -4618 52634
rect -4534 52398 -4298 52634
rect -4854 16718 -4618 16954
rect -4534 16718 -4298 16954
rect -4854 16398 -4618 16634
rect -4534 16398 -4298 16634
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 696218 -3658 696454
rect -3574 696218 -3338 696454
rect -3894 695898 -3658 696134
rect -3574 695898 -3338 696134
rect -3894 660218 -3658 660454
rect -3574 660218 -3338 660454
rect -3894 659898 -3658 660134
rect -3574 659898 -3338 660134
rect -3894 624218 -3658 624454
rect -3574 624218 -3338 624454
rect -3894 623898 -3658 624134
rect -3574 623898 -3338 624134
rect -3894 588218 -3658 588454
rect -3574 588218 -3338 588454
rect -3894 587898 -3658 588134
rect -3574 587898 -3338 588134
rect -3894 552218 -3658 552454
rect -3574 552218 -3338 552454
rect -3894 551898 -3658 552134
rect -3574 551898 -3338 552134
rect -3894 516218 -3658 516454
rect -3574 516218 -3338 516454
rect -3894 515898 -3658 516134
rect -3574 515898 -3338 516134
rect -3894 480218 -3658 480454
rect -3574 480218 -3338 480454
rect -3894 479898 -3658 480134
rect -3574 479898 -3338 480134
rect -3894 444218 -3658 444454
rect -3574 444218 -3338 444454
rect -3894 443898 -3658 444134
rect -3574 443898 -3338 444134
rect -3894 408218 -3658 408454
rect -3574 408218 -3338 408454
rect -3894 407898 -3658 408134
rect -3574 407898 -3338 408134
rect -3894 372218 -3658 372454
rect -3574 372218 -3338 372454
rect -3894 371898 -3658 372134
rect -3574 371898 -3338 372134
rect -3894 336218 -3658 336454
rect -3574 336218 -3338 336454
rect -3894 335898 -3658 336134
rect -3574 335898 -3338 336134
rect -3894 300218 -3658 300454
rect -3574 300218 -3338 300454
rect -3894 299898 -3658 300134
rect -3574 299898 -3338 300134
rect -3894 264218 -3658 264454
rect -3574 264218 -3338 264454
rect -3894 263898 -3658 264134
rect -3574 263898 -3338 264134
rect -3894 228218 -3658 228454
rect -3574 228218 -3338 228454
rect -3894 227898 -3658 228134
rect -3574 227898 -3338 228134
rect -3894 192218 -3658 192454
rect -3574 192218 -3338 192454
rect -3894 191898 -3658 192134
rect -3574 191898 -3338 192134
rect -3894 156218 -3658 156454
rect -3574 156218 -3338 156454
rect -3894 155898 -3658 156134
rect -3574 155898 -3338 156134
rect -3894 120218 -3658 120454
rect -3574 120218 -3338 120454
rect -3894 119898 -3658 120134
rect -3574 119898 -3338 120134
rect -3894 84218 -3658 84454
rect -3574 84218 -3338 84454
rect -3894 83898 -3658 84134
rect -3574 83898 -3338 84134
rect -3894 48218 -3658 48454
rect -3574 48218 -3338 48454
rect -3894 47898 -3658 48134
rect -3574 47898 -3338 48134
rect -3894 12218 -3658 12454
rect -3574 12218 -3338 12454
rect -3894 11898 -3658 12134
rect -3574 11898 -3338 12134
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 691718 -2698 691954
rect -2614 691718 -2378 691954
rect -2934 691398 -2698 691634
rect -2614 691398 -2378 691634
rect -2934 655718 -2698 655954
rect -2614 655718 -2378 655954
rect -2934 655398 -2698 655634
rect -2614 655398 -2378 655634
rect -2934 619718 -2698 619954
rect -2614 619718 -2378 619954
rect -2934 619398 -2698 619634
rect -2614 619398 -2378 619634
rect -2934 583718 -2698 583954
rect -2614 583718 -2378 583954
rect -2934 583398 -2698 583634
rect -2614 583398 -2378 583634
rect -2934 547718 -2698 547954
rect -2614 547718 -2378 547954
rect -2934 547398 -2698 547634
rect -2614 547398 -2378 547634
rect -2934 511718 -2698 511954
rect -2614 511718 -2378 511954
rect -2934 511398 -2698 511634
rect -2614 511398 -2378 511634
rect -2934 475718 -2698 475954
rect -2614 475718 -2378 475954
rect -2934 475398 -2698 475634
rect -2614 475398 -2378 475634
rect -2934 439718 -2698 439954
rect -2614 439718 -2378 439954
rect -2934 439398 -2698 439634
rect -2614 439398 -2378 439634
rect -2934 403718 -2698 403954
rect -2614 403718 -2378 403954
rect -2934 403398 -2698 403634
rect -2614 403398 -2378 403634
rect -2934 367718 -2698 367954
rect -2614 367718 -2378 367954
rect -2934 367398 -2698 367634
rect -2614 367398 -2378 367634
rect -2934 331718 -2698 331954
rect -2614 331718 -2378 331954
rect -2934 331398 -2698 331634
rect -2614 331398 -2378 331634
rect -2934 295718 -2698 295954
rect -2614 295718 -2378 295954
rect -2934 295398 -2698 295634
rect -2614 295398 -2378 295634
rect -2934 259718 -2698 259954
rect -2614 259718 -2378 259954
rect -2934 259398 -2698 259634
rect -2614 259398 -2378 259634
rect -2934 223718 -2698 223954
rect -2614 223718 -2378 223954
rect -2934 223398 -2698 223634
rect -2614 223398 -2378 223634
rect -2934 187718 -2698 187954
rect -2614 187718 -2378 187954
rect -2934 187398 -2698 187634
rect -2614 187398 -2378 187634
rect -2934 151718 -2698 151954
rect -2614 151718 -2378 151954
rect -2934 151398 -2698 151634
rect -2614 151398 -2378 151634
rect -2934 115718 -2698 115954
rect -2614 115718 -2378 115954
rect -2934 115398 -2698 115634
rect -2614 115398 -2378 115634
rect -2934 79718 -2698 79954
rect -2614 79718 -2378 79954
rect -2934 79398 -2698 79634
rect -2614 79398 -2378 79634
rect -2934 43718 -2698 43954
rect -2614 43718 -2378 43954
rect -2934 43398 -2698 43634
rect -2614 43398 -2378 43634
rect -2934 7718 -2698 7954
rect -2614 7718 -2378 7954
rect -2934 7398 -2698 7634
rect -2614 7398 -2378 7634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 6326 705562 6562 705798
rect 6646 705562 6882 705798
rect 6326 705242 6562 705478
rect 6646 705242 6882 705478
rect 6326 691718 6562 691954
rect 6646 691718 6882 691954
rect 6326 691398 6562 691634
rect 6646 691398 6882 691634
rect 6326 655718 6562 655954
rect 6646 655718 6882 655954
rect 6326 655398 6562 655634
rect 6646 655398 6882 655634
rect 6326 619718 6562 619954
rect 6646 619718 6882 619954
rect 6326 619398 6562 619634
rect 6646 619398 6882 619634
rect 6326 583718 6562 583954
rect 6646 583718 6882 583954
rect 6326 583398 6562 583634
rect 6646 583398 6882 583634
rect 6326 547718 6562 547954
rect 6646 547718 6882 547954
rect 6326 547398 6562 547634
rect 6646 547398 6882 547634
rect 6326 511718 6562 511954
rect 6646 511718 6882 511954
rect 6326 511398 6562 511634
rect 6646 511398 6882 511634
rect 6326 475718 6562 475954
rect 6646 475718 6882 475954
rect 6326 475398 6562 475634
rect 6646 475398 6882 475634
rect 6326 439718 6562 439954
rect 6646 439718 6882 439954
rect 6326 439398 6562 439634
rect 6646 439398 6882 439634
rect 6326 403718 6562 403954
rect 6646 403718 6882 403954
rect 6326 403398 6562 403634
rect 6646 403398 6882 403634
rect 6326 367718 6562 367954
rect 6646 367718 6882 367954
rect 6326 367398 6562 367634
rect 6646 367398 6882 367634
rect 6326 331718 6562 331954
rect 6646 331718 6882 331954
rect 6326 331398 6562 331634
rect 6646 331398 6882 331634
rect 6326 295718 6562 295954
rect 6646 295718 6882 295954
rect 6326 295398 6562 295634
rect 6646 295398 6882 295634
rect 6326 259718 6562 259954
rect 6646 259718 6882 259954
rect 6326 259398 6562 259634
rect 6646 259398 6882 259634
rect 6326 223718 6562 223954
rect 6646 223718 6882 223954
rect 6326 223398 6562 223634
rect 6646 223398 6882 223634
rect 6326 187718 6562 187954
rect 6646 187718 6882 187954
rect 6326 187398 6562 187634
rect 6646 187398 6882 187634
rect 6326 151718 6562 151954
rect 6646 151718 6882 151954
rect 6326 151398 6562 151634
rect 6646 151398 6882 151634
rect 6326 115718 6562 115954
rect 6646 115718 6882 115954
rect 6326 115398 6562 115634
rect 6646 115398 6882 115634
rect 6326 79718 6562 79954
rect 6646 79718 6882 79954
rect 6326 79398 6562 79634
rect 6646 79398 6882 79634
rect 6326 43718 6562 43954
rect 6646 43718 6882 43954
rect 6326 43398 6562 43634
rect 6646 43398 6882 43634
rect 6326 7718 6562 7954
rect 6646 7718 6882 7954
rect 6326 7398 6562 7634
rect 6646 7398 6882 7634
rect 6326 -1542 6562 -1306
rect 6646 -1542 6882 -1306
rect 6326 -1862 6562 -1626
rect 6646 -1862 6882 -1626
rect 10826 706522 11062 706758
rect 11146 706522 11382 706758
rect 10826 706202 11062 706438
rect 11146 706202 11382 706438
rect 10826 696218 11062 696454
rect 11146 696218 11382 696454
rect 10826 695898 11062 696134
rect 11146 695898 11382 696134
rect 10826 660218 11062 660454
rect 11146 660218 11382 660454
rect 10826 659898 11062 660134
rect 11146 659898 11382 660134
rect 10826 624218 11062 624454
rect 11146 624218 11382 624454
rect 10826 623898 11062 624134
rect 11146 623898 11382 624134
rect 10826 588218 11062 588454
rect 11146 588218 11382 588454
rect 10826 587898 11062 588134
rect 11146 587898 11382 588134
rect 10826 552218 11062 552454
rect 11146 552218 11382 552454
rect 10826 551898 11062 552134
rect 11146 551898 11382 552134
rect 10826 516218 11062 516454
rect 11146 516218 11382 516454
rect 10826 515898 11062 516134
rect 11146 515898 11382 516134
rect 10826 480218 11062 480454
rect 11146 480218 11382 480454
rect 10826 479898 11062 480134
rect 11146 479898 11382 480134
rect 10826 444218 11062 444454
rect 11146 444218 11382 444454
rect 10826 443898 11062 444134
rect 11146 443898 11382 444134
rect 10826 408218 11062 408454
rect 11146 408218 11382 408454
rect 10826 407898 11062 408134
rect 11146 407898 11382 408134
rect 10826 372218 11062 372454
rect 11146 372218 11382 372454
rect 10826 371898 11062 372134
rect 11146 371898 11382 372134
rect 10826 336218 11062 336454
rect 11146 336218 11382 336454
rect 10826 335898 11062 336134
rect 11146 335898 11382 336134
rect 10826 300218 11062 300454
rect 11146 300218 11382 300454
rect 10826 299898 11062 300134
rect 11146 299898 11382 300134
rect 10826 264218 11062 264454
rect 11146 264218 11382 264454
rect 10826 263898 11062 264134
rect 11146 263898 11382 264134
rect 10826 228218 11062 228454
rect 11146 228218 11382 228454
rect 10826 227898 11062 228134
rect 11146 227898 11382 228134
rect 10826 192218 11062 192454
rect 11146 192218 11382 192454
rect 10826 191898 11062 192134
rect 11146 191898 11382 192134
rect 10826 156218 11062 156454
rect 11146 156218 11382 156454
rect 10826 155898 11062 156134
rect 11146 155898 11382 156134
rect 10826 120218 11062 120454
rect 11146 120218 11382 120454
rect 10826 119898 11062 120134
rect 11146 119898 11382 120134
rect 10826 84218 11062 84454
rect 11146 84218 11382 84454
rect 10826 83898 11062 84134
rect 11146 83898 11382 84134
rect 10826 48218 11062 48454
rect 11146 48218 11382 48454
rect 10826 47898 11062 48134
rect 11146 47898 11382 48134
rect 10826 12218 11062 12454
rect 11146 12218 11382 12454
rect 10826 11898 11062 12134
rect 11146 11898 11382 12134
rect 10826 -2502 11062 -2266
rect 11146 -2502 11382 -2266
rect 10826 -2822 11062 -2586
rect 11146 -2822 11382 -2586
rect 15326 707482 15562 707718
rect 15646 707482 15882 707718
rect 15326 707162 15562 707398
rect 15646 707162 15882 707398
rect 15326 700718 15562 700954
rect 15646 700718 15882 700954
rect 15326 700398 15562 700634
rect 15646 700398 15882 700634
rect 15326 664718 15562 664954
rect 15646 664718 15882 664954
rect 15326 664398 15562 664634
rect 15646 664398 15882 664634
rect 15326 628718 15562 628954
rect 15646 628718 15882 628954
rect 15326 628398 15562 628634
rect 15646 628398 15882 628634
rect 15326 592718 15562 592954
rect 15646 592718 15882 592954
rect 15326 592398 15562 592634
rect 15646 592398 15882 592634
rect 15326 556718 15562 556954
rect 15646 556718 15882 556954
rect 15326 556398 15562 556634
rect 15646 556398 15882 556634
rect 15326 520718 15562 520954
rect 15646 520718 15882 520954
rect 15326 520398 15562 520634
rect 15646 520398 15882 520634
rect 15326 484718 15562 484954
rect 15646 484718 15882 484954
rect 15326 484398 15562 484634
rect 15646 484398 15882 484634
rect 15326 448718 15562 448954
rect 15646 448718 15882 448954
rect 15326 448398 15562 448634
rect 15646 448398 15882 448634
rect 15326 412718 15562 412954
rect 15646 412718 15882 412954
rect 15326 412398 15562 412634
rect 15646 412398 15882 412634
rect 15326 376718 15562 376954
rect 15646 376718 15882 376954
rect 15326 376398 15562 376634
rect 15646 376398 15882 376634
rect 15326 340718 15562 340954
rect 15646 340718 15882 340954
rect 15326 340398 15562 340634
rect 15646 340398 15882 340634
rect 15326 304718 15562 304954
rect 15646 304718 15882 304954
rect 15326 304398 15562 304634
rect 15646 304398 15882 304634
rect 15326 268718 15562 268954
rect 15646 268718 15882 268954
rect 15326 268398 15562 268634
rect 15646 268398 15882 268634
rect 15326 232718 15562 232954
rect 15646 232718 15882 232954
rect 15326 232398 15562 232634
rect 15646 232398 15882 232634
rect 15326 196718 15562 196954
rect 15646 196718 15882 196954
rect 15326 196398 15562 196634
rect 15646 196398 15882 196634
rect 15326 160718 15562 160954
rect 15646 160718 15882 160954
rect 15326 160398 15562 160634
rect 15646 160398 15882 160634
rect 15326 124718 15562 124954
rect 15646 124718 15882 124954
rect 15326 124398 15562 124634
rect 15646 124398 15882 124634
rect 15326 88718 15562 88954
rect 15646 88718 15882 88954
rect 15326 88398 15562 88634
rect 15646 88398 15882 88634
rect 15326 52718 15562 52954
rect 15646 52718 15882 52954
rect 15326 52398 15562 52634
rect 15646 52398 15882 52634
rect 15326 16718 15562 16954
rect 15646 16718 15882 16954
rect 15326 16398 15562 16634
rect 15646 16398 15882 16634
rect 15326 -3462 15562 -3226
rect 15646 -3462 15882 -3226
rect 15326 -3782 15562 -3546
rect 15646 -3782 15882 -3546
rect 19826 708442 20062 708678
rect 20146 708442 20382 708678
rect 19826 708122 20062 708358
rect 20146 708122 20382 708358
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -4422 20062 -4186
rect 20146 -4422 20382 -4186
rect 19826 -4742 20062 -4506
rect 20146 -4742 20382 -4506
rect 24326 709402 24562 709638
rect 24646 709402 24882 709638
rect 24326 709082 24562 709318
rect 24646 709082 24882 709318
rect 24326 673718 24562 673954
rect 24646 673718 24882 673954
rect 24326 673398 24562 673634
rect 24646 673398 24882 673634
rect 24326 637718 24562 637954
rect 24646 637718 24882 637954
rect 24326 637398 24562 637634
rect 24646 637398 24882 637634
rect 24326 601718 24562 601954
rect 24646 601718 24882 601954
rect 24326 601398 24562 601634
rect 24646 601398 24882 601634
rect 24326 565718 24562 565954
rect 24646 565718 24882 565954
rect 24326 565398 24562 565634
rect 24646 565398 24882 565634
rect 24326 529718 24562 529954
rect 24646 529718 24882 529954
rect 24326 529398 24562 529634
rect 24646 529398 24882 529634
rect 24326 493718 24562 493954
rect 24646 493718 24882 493954
rect 24326 493398 24562 493634
rect 24646 493398 24882 493634
rect 24326 457718 24562 457954
rect 24646 457718 24882 457954
rect 24326 457398 24562 457634
rect 24646 457398 24882 457634
rect 24326 421718 24562 421954
rect 24646 421718 24882 421954
rect 24326 421398 24562 421634
rect 24646 421398 24882 421634
rect 24326 385718 24562 385954
rect 24646 385718 24882 385954
rect 24326 385398 24562 385634
rect 24646 385398 24882 385634
rect 24326 349718 24562 349954
rect 24646 349718 24882 349954
rect 24326 349398 24562 349634
rect 24646 349398 24882 349634
rect 24326 313718 24562 313954
rect 24646 313718 24882 313954
rect 24326 313398 24562 313634
rect 24646 313398 24882 313634
rect 24326 277718 24562 277954
rect 24646 277718 24882 277954
rect 24326 277398 24562 277634
rect 24646 277398 24882 277634
rect 24326 241718 24562 241954
rect 24646 241718 24882 241954
rect 24326 241398 24562 241634
rect 24646 241398 24882 241634
rect 24326 205718 24562 205954
rect 24646 205718 24882 205954
rect 24326 205398 24562 205634
rect 24646 205398 24882 205634
rect 24326 169718 24562 169954
rect 24646 169718 24882 169954
rect 24326 169398 24562 169634
rect 24646 169398 24882 169634
rect 24326 133718 24562 133954
rect 24646 133718 24882 133954
rect 24326 133398 24562 133634
rect 24646 133398 24882 133634
rect 24326 97718 24562 97954
rect 24646 97718 24882 97954
rect 24326 97398 24562 97634
rect 24646 97398 24882 97634
rect 24326 61718 24562 61954
rect 24646 61718 24882 61954
rect 24326 61398 24562 61634
rect 24646 61398 24882 61634
rect 24326 25718 24562 25954
rect 24646 25718 24882 25954
rect 24326 25398 24562 25634
rect 24646 25398 24882 25634
rect 24326 -5382 24562 -5146
rect 24646 -5382 24882 -5146
rect 24326 -5702 24562 -5466
rect 24646 -5702 24882 -5466
rect 28826 710362 29062 710598
rect 29146 710362 29382 710598
rect 28826 710042 29062 710278
rect 29146 710042 29382 710278
rect 28826 678218 29062 678454
rect 29146 678218 29382 678454
rect 28826 677898 29062 678134
rect 29146 677898 29382 678134
rect 28826 642218 29062 642454
rect 29146 642218 29382 642454
rect 28826 641898 29062 642134
rect 29146 641898 29382 642134
rect 28826 606218 29062 606454
rect 29146 606218 29382 606454
rect 28826 605898 29062 606134
rect 29146 605898 29382 606134
rect 28826 570218 29062 570454
rect 29146 570218 29382 570454
rect 28826 569898 29062 570134
rect 29146 569898 29382 570134
rect 28826 534218 29062 534454
rect 29146 534218 29382 534454
rect 28826 533898 29062 534134
rect 29146 533898 29382 534134
rect 28826 498218 29062 498454
rect 29146 498218 29382 498454
rect 28826 497898 29062 498134
rect 29146 497898 29382 498134
rect 28826 462218 29062 462454
rect 29146 462218 29382 462454
rect 28826 461898 29062 462134
rect 29146 461898 29382 462134
rect 28826 426218 29062 426454
rect 29146 426218 29382 426454
rect 28826 425898 29062 426134
rect 29146 425898 29382 426134
rect 28826 390218 29062 390454
rect 29146 390218 29382 390454
rect 28826 389898 29062 390134
rect 29146 389898 29382 390134
rect 28826 354218 29062 354454
rect 29146 354218 29382 354454
rect 28826 353898 29062 354134
rect 29146 353898 29382 354134
rect 28826 318218 29062 318454
rect 29146 318218 29382 318454
rect 28826 317898 29062 318134
rect 29146 317898 29382 318134
rect 28826 282218 29062 282454
rect 29146 282218 29382 282454
rect 28826 281898 29062 282134
rect 29146 281898 29382 282134
rect 28826 246218 29062 246454
rect 29146 246218 29382 246454
rect 28826 245898 29062 246134
rect 29146 245898 29382 246134
rect 28826 210218 29062 210454
rect 29146 210218 29382 210454
rect 28826 209898 29062 210134
rect 29146 209898 29382 210134
rect 28826 174218 29062 174454
rect 29146 174218 29382 174454
rect 28826 173898 29062 174134
rect 29146 173898 29382 174134
rect 28826 138218 29062 138454
rect 29146 138218 29382 138454
rect 28826 137898 29062 138134
rect 29146 137898 29382 138134
rect 28826 102218 29062 102454
rect 29146 102218 29382 102454
rect 28826 101898 29062 102134
rect 29146 101898 29382 102134
rect 28826 66218 29062 66454
rect 29146 66218 29382 66454
rect 28826 65898 29062 66134
rect 29146 65898 29382 66134
rect 28826 30218 29062 30454
rect 29146 30218 29382 30454
rect 28826 29898 29062 30134
rect 29146 29898 29382 30134
rect 28826 -6342 29062 -6106
rect 29146 -6342 29382 -6106
rect 28826 -6662 29062 -6426
rect 29146 -6662 29382 -6426
rect 33326 711322 33562 711558
rect 33646 711322 33882 711558
rect 33326 711002 33562 711238
rect 33646 711002 33882 711238
rect 33326 682718 33562 682954
rect 33646 682718 33882 682954
rect 33326 682398 33562 682634
rect 33646 682398 33882 682634
rect 33326 646718 33562 646954
rect 33646 646718 33882 646954
rect 33326 646398 33562 646634
rect 33646 646398 33882 646634
rect 33326 610718 33562 610954
rect 33646 610718 33882 610954
rect 33326 610398 33562 610634
rect 33646 610398 33882 610634
rect 33326 574718 33562 574954
rect 33646 574718 33882 574954
rect 33326 574398 33562 574634
rect 33646 574398 33882 574634
rect 33326 538718 33562 538954
rect 33646 538718 33882 538954
rect 33326 538398 33562 538634
rect 33646 538398 33882 538634
rect 33326 502718 33562 502954
rect 33646 502718 33882 502954
rect 33326 502398 33562 502634
rect 33646 502398 33882 502634
rect 33326 466718 33562 466954
rect 33646 466718 33882 466954
rect 33326 466398 33562 466634
rect 33646 466398 33882 466634
rect 33326 430718 33562 430954
rect 33646 430718 33882 430954
rect 33326 430398 33562 430634
rect 33646 430398 33882 430634
rect 33326 394718 33562 394954
rect 33646 394718 33882 394954
rect 33326 394398 33562 394634
rect 33646 394398 33882 394634
rect 33326 358718 33562 358954
rect 33646 358718 33882 358954
rect 33326 358398 33562 358634
rect 33646 358398 33882 358634
rect 33326 322718 33562 322954
rect 33646 322718 33882 322954
rect 33326 322398 33562 322634
rect 33646 322398 33882 322634
rect 33326 286718 33562 286954
rect 33646 286718 33882 286954
rect 33326 286398 33562 286634
rect 33646 286398 33882 286634
rect 33326 250718 33562 250954
rect 33646 250718 33882 250954
rect 33326 250398 33562 250634
rect 33646 250398 33882 250634
rect 33326 214718 33562 214954
rect 33646 214718 33882 214954
rect 33326 214398 33562 214634
rect 33646 214398 33882 214634
rect 33326 178718 33562 178954
rect 33646 178718 33882 178954
rect 33326 178398 33562 178634
rect 33646 178398 33882 178634
rect 33326 142718 33562 142954
rect 33646 142718 33882 142954
rect 33326 142398 33562 142634
rect 33646 142398 33882 142634
rect 33326 106718 33562 106954
rect 33646 106718 33882 106954
rect 33326 106398 33562 106634
rect 33646 106398 33882 106634
rect 33326 70718 33562 70954
rect 33646 70718 33882 70954
rect 33326 70398 33562 70634
rect 33646 70398 33882 70634
rect 33326 34718 33562 34954
rect 33646 34718 33882 34954
rect 33326 34398 33562 34634
rect 33646 34398 33882 34634
rect 33326 -7302 33562 -7066
rect 33646 -7302 33882 -7066
rect 33326 -7622 33562 -7386
rect 33646 -7622 33882 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 42326 705562 42562 705798
rect 42646 705562 42882 705798
rect 42326 705242 42562 705478
rect 42646 705242 42882 705478
rect 42326 691718 42562 691954
rect 42646 691718 42882 691954
rect 42326 691398 42562 691634
rect 42646 691398 42882 691634
rect 42326 655718 42562 655954
rect 42646 655718 42882 655954
rect 42326 655398 42562 655634
rect 42646 655398 42882 655634
rect 42326 619718 42562 619954
rect 42646 619718 42882 619954
rect 42326 619398 42562 619634
rect 42646 619398 42882 619634
rect 42326 583718 42562 583954
rect 42646 583718 42882 583954
rect 42326 583398 42562 583634
rect 42646 583398 42882 583634
rect 42326 547718 42562 547954
rect 42646 547718 42882 547954
rect 42326 547398 42562 547634
rect 42646 547398 42882 547634
rect 42326 511718 42562 511954
rect 42646 511718 42882 511954
rect 42326 511398 42562 511634
rect 42646 511398 42882 511634
rect 42326 475718 42562 475954
rect 42646 475718 42882 475954
rect 42326 475398 42562 475634
rect 42646 475398 42882 475634
rect 42326 439718 42562 439954
rect 42646 439718 42882 439954
rect 42326 439398 42562 439634
rect 42646 439398 42882 439634
rect 42326 403718 42562 403954
rect 42646 403718 42882 403954
rect 42326 403398 42562 403634
rect 42646 403398 42882 403634
rect 42326 367718 42562 367954
rect 42646 367718 42882 367954
rect 42326 367398 42562 367634
rect 42646 367398 42882 367634
rect 42326 331718 42562 331954
rect 42646 331718 42882 331954
rect 42326 331398 42562 331634
rect 42646 331398 42882 331634
rect 42326 295718 42562 295954
rect 42646 295718 42882 295954
rect 42326 295398 42562 295634
rect 42646 295398 42882 295634
rect 42326 259718 42562 259954
rect 42646 259718 42882 259954
rect 42326 259398 42562 259634
rect 42646 259398 42882 259634
rect 42326 223718 42562 223954
rect 42646 223718 42882 223954
rect 42326 223398 42562 223634
rect 42646 223398 42882 223634
rect 42326 187718 42562 187954
rect 42646 187718 42882 187954
rect 42326 187398 42562 187634
rect 42646 187398 42882 187634
rect 42326 151718 42562 151954
rect 42646 151718 42882 151954
rect 42326 151398 42562 151634
rect 42646 151398 42882 151634
rect 42326 115718 42562 115954
rect 42646 115718 42882 115954
rect 42326 115398 42562 115634
rect 42646 115398 42882 115634
rect 42326 79718 42562 79954
rect 42646 79718 42882 79954
rect 42326 79398 42562 79634
rect 42646 79398 42882 79634
rect 42326 43718 42562 43954
rect 42646 43718 42882 43954
rect 42326 43398 42562 43634
rect 42646 43398 42882 43634
rect 42326 7718 42562 7954
rect 42646 7718 42882 7954
rect 42326 7398 42562 7634
rect 42646 7398 42882 7634
rect 42326 -1542 42562 -1306
rect 42646 -1542 42882 -1306
rect 42326 -1862 42562 -1626
rect 42646 -1862 42882 -1626
rect 46826 706522 47062 706758
rect 47146 706522 47382 706758
rect 46826 706202 47062 706438
rect 47146 706202 47382 706438
rect 46826 696218 47062 696454
rect 47146 696218 47382 696454
rect 46826 695898 47062 696134
rect 47146 695898 47382 696134
rect 51326 707482 51562 707718
rect 51646 707482 51882 707718
rect 51326 707162 51562 707398
rect 51646 707162 51882 707398
rect 51326 700718 51562 700954
rect 51646 700718 51882 700954
rect 51326 700398 51562 700634
rect 51646 700398 51882 700634
rect 51326 664718 51562 664954
rect 51646 664718 51882 664954
rect 51326 664398 51562 664634
rect 51646 664398 51882 664634
rect 55826 708442 56062 708678
rect 56146 708442 56382 708678
rect 55826 708122 56062 708358
rect 56146 708122 56382 708358
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 60326 709402 60562 709638
rect 60646 709402 60882 709638
rect 60326 709082 60562 709318
rect 60646 709082 60882 709318
rect 60326 673718 60562 673954
rect 60646 673718 60882 673954
rect 60326 673398 60562 673634
rect 60646 673398 60882 673634
rect 64826 710362 65062 710598
rect 65146 710362 65382 710598
rect 64826 710042 65062 710278
rect 65146 710042 65382 710278
rect 64826 678218 65062 678454
rect 65146 678218 65382 678454
rect 64826 677898 65062 678134
rect 65146 677898 65382 678134
rect 69326 711322 69562 711558
rect 69646 711322 69882 711558
rect 69326 711002 69562 711238
rect 69646 711002 69882 711238
rect 69326 682718 69562 682954
rect 69646 682718 69882 682954
rect 69326 682398 69562 682634
rect 69646 682398 69882 682634
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 78326 705562 78562 705798
rect 78646 705562 78882 705798
rect 78326 705242 78562 705478
rect 78646 705242 78882 705478
rect 78326 691718 78562 691954
rect 78646 691718 78882 691954
rect 78326 691398 78562 691634
rect 78646 691398 78882 691634
rect 82826 706522 83062 706758
rect 83146 706522 83382 706758
rect 82826 706202 83062 706438
rect 83146 706202 83382 706438
rect 82826 696218 83062 696454
rect 83146 696218 83382 696454
rect 82826 695898 83062 696134
rect 83146 695898 83382 696134
rect 87326 707482 87562 707718
rect 87646 707482 87882 707718
rect 87326 707162 87562 707398
rect 87646 707162 87882 707398
rect 87326 700718 87562 700954
rect 87646 700718 87882 700954
rect 87326 700398 87562 700634
rect 87646 700398 87882 700634
rect 87326 664718 87562 664954
rect 87646 664718 87882 664954
rect 87326 664398 87562 664634
rect 87646 664398 87882 664634
rect 91826 708442 92062 708678
rect 92146 708442 92382 708678
rect 91826 708122 92062 708358
rect 92146 708122 92382 708358
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 96326 709402 96562 709638
rect 96646 709402 96882 709638
rect 96326 709082 96562 709318
rect 96646 709082 96882 709318
rect 96326 673718 96562 673954
rect 96646 673718 96882 673954
rect 96326 673398 96562 673634
rect 96646 673398 96882 673634
rect 100826 710362 101062 710598
rect 101146 710362 101382 710598
rect 100826 710042 101062 710278
rect 101146 710042 101382 710278
rect 100826 678218 101062 678454
rect 101146 678218 101382 678454
rect 100826 677898 101062 678134
rect 101146 677898 101382 678134
rect 105326 711322 105562 711558
rect 105646 711322 105882 711558
rect 105326 711002 105562 711238
rect 105646 711002 105882 711238
rect 105326 682718 105562 682954
rect 105646 682718 105882 682954
rect 105326 682398 105562 682634
rect 105646 682398 105882 682634
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 114326 705562 114562 705798
rect 114646 705562 114882 705798
rect 114326 705242 114562 705478
rect 114646 705242 114882 705478
rect 114326 691718 114562 691954
rect 114646 691718 114882 691954
rect 114326 691398 114562 691634
rect 114646 691398 114882 691634
rect 118826 706522 119062 706758
rect 119146 706522 119382 706758
rect 118826 706202 119062 706438
rect 119146 706202 119382 706438
rect 118826 696218 119062 696454
rect 119146 696218 119382 696454
rect 118826 695898 119062 696134
rect 119146 695898 119382 696134
rect 123326 707482 123562 707718
rect 123646 707482 123882 707718
rect 123326 707162 123562 707398
rect 123646 707162 123882 707398
rect 123326 700718 123562 700954
rect 123646 700718 123882 700954
rect 123326 700398 123562 700634
rect 123646 700398 123882 700634
rect 123326 664718 123562 664954
rect 123646 664718 123882 664954
rect 123326 664398 123562 664634
rect 123646 664398 123882 664634
rect 127826 708442 128062 708678
rect 128146 708442 128382 708678
rect 127826 708122 128062 708358
rect 128146 708122 128382 708358
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 132326 709402 132562 709638
rect 132646 709402 132882 709638
rect 132326 709082 132562 709318
rect 132646 709082 132882 709318
rect 132326 673718 132562 673954
rect 132646 673718 132882 673954
rect 132326 673398 132562 673634
rect 132646 673398 132882 673634
rect 136826 710362 137062 710598
rect 137146 710362 137382 710598
rect 136826 710042 137062 710278
rect 137146 710042 137382 710278
rect 136826 678218 137062 678454
rect 137146 678218 137382 678454
rect 136826 677898 137062 678134
rect 137146 677898 137382 678134
rect 141326 711322 141562 711558
rect 141646 711322 141882 711558
rect 141326 711002 141562 711238
rect 141646 711002 141882 711238
rect 141326 682718 141562 682954
rect 141646 682718 141882 682954
rect 141326 682398 141562 682634
rect 141646 682398 141882 682634
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 150326 705562 150562 705798
rect 150646 705562 150882 705798
rect 150326 705242 150562 705478
rect 150646 705242 150882 705478
rect 150326 691718 150562 691954
rect 150646 691718 150882 691954
rect 150326 691398 150562 691634
rect 150646 691398 150882 691634
rect 154826 706522 155062 706758
rect 155146 706522 155382 706758
rect 154826 706202 155062 706438
rect 155146 706202 155382 706438
rect 154826 696218 155062 696454
rect 155146 696218 155382 696454
rect 154826 695898 155062 696134
rect 155146 695898 155382 696134
rect 159326 707482 159562 707718
rect 159646 707482 159882 707718
rect 159326 707162 159562 707398
rect 159646 707162 159882 707398
rect 159326 700718 159562 700954
rect 159646 700718 159882 700954
rect 159326 700398 159562 700634
rect 159646 700398 159882 700634
rect 159326 664718 159562 664954
rect 159646 664718 159882 664954
rect 159326 664398 159562 664634
rect 159646 664398 159882 664634
rect 163826 708442 164062 708678
rect 164146 708442 164382 708678
rect 163826 708122 164062 708358
rect 164146 708122 164382 708358
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 168326 709402 168562 709638
rect 168646 709402 168882 709638
rect 168326 709082 168562 709318
rect 168646 709082 168882 709318
rect 168326 673718 168562 673954
rect 168646 673718 168882 673954
rect 168326 673398 168562 673634
rect 168646 673398 168882 673634
rect 172826 710362 173062 710598
rect 173146 710362 173382 710598
rect 172826 710042 173062 710278
rect 173146 710042 173382 710278
rect 172826 678218 173062 678454
rect 173146 678218 173382 678454
rect 172826 677898 173062 678134
rect 173146 677898 173382 678134
rect 177326 711322 177562 711558
rect 177646 711322 177882 711558
rect 177326 711002 177562 711238
rect 177646 711002 177882 711238
rect 177326 682718 177562 682954
rect 177646 682718 177882 682954
rect 177326 682398 177562 682634
rect 177646 682398 177882 682634
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 186326 705562 186562 705798
rect 186646 705562 186882 705798
rect 186326 705242 186562 705478
rect 186646 705242 186882 705478
rect 186326 691718 186562 691954
rect 186646 691718 186882 691954
rect 186326 691398 186562 691634
rect 186646 691398 186882 691634
rect 190826 706522 191062 706758
rect 191146 706522 191382 706758
rect 190826 706202 191062 706438
rect 191146 706202 191382 706438
rect 190826 696218 191062 696454
rect 191146 696218 191382 696454
rect 190826 695898 191062 696134
rect 191146 695898 191382 696134
rect 195326 707482 195562 707718
rect 195646 707482 195882 707718
rect 195326 707162 195562 707398
rect 195646 707162 195882 707398
rect 195326 700718 195562 700954
rect 195646 700718 195882 700954
rect 195326 700398 195562 700634
rect 195646 700398 195882 700634
rect 195326 664718 195562 664954
rect 195646 664718 195882 664954
rect 195326 664398 195562 664634
rect 195646 664398 195882 664634
rect 199826 708442 200062 708678
rect 200146 708442 200382 708678
rect 199826 708122 200062 708358
rect 200146 708122 200382 708358
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 204326 709402 204562 709638
rect 204646 709402 204882 709638
rect 204326 709082 204562 709318
rect 204646 709082 204882 709318
rect 204326 673718 204562 673954
rect 204646 673718 204882 673954
rect 204326 673398 204562 673634
rect 204646 673398 204882 673634
rect 208826 710362 209062 710598
rect 209146 710362 209382 710598
rect 208826 710042 209062 710278
rect 209146 710042 209382 710278
rect 208826 678218 209062 678454
rect 209146 678218 209382 678454
rect 208826 677898 209062 678134
rect 209146 677898 209382 678134
rect 213326 711322 213562 711558
rect 213646 711322 213882 711558
rect 213326 711002 213562 711238
rect 213646 711002 213882 711238
rect 213326 682718 213562 682954
rect 213646 682718 213882 682954
rect 213326 682398 213562 682634
rect 213646 682398 213882 682634
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 222326 705562 222562 705798
rect 222646 705562 222882 705798
rect 222326 705242 222562 705478
rect 222646 705242 222882 705478
rect 222326 691718 222562 691954
rect 222646 691718 222882 691954
rect 222326 691398 222562 691634
rect 222646 691398 222882 691634
rect 226826 706522 227062 706758
rect 227146 706522 227382 706758
rect 226826 706202 227062 706438
rect 227146 706202 227382 706438
rect 226826 696218 227062 696454
rect 227146 696218 227382 696454
rect 226826 695898 227062 696134
rect 227146 695898 227382 696134
rect 231326 707482 231562 707718
rect 231646 707482 231882 707718
rect 231326 707162 231562 707398
rect 231646 707162 231882 707398
rect 231326 700718 231562 700954
rect 231646 700718 231882 700954
rect 231326 700398 231562 700634
rect 231646 700398 231882 700634
rect 231326 664718 231562 664954
rect 231646 664718 231882 664954
rect 231326 664398 231562 664634
rect 231646 664398 231882 664634
rect 235826 708442 236062 708678
rect 236146 708442 236382 708678
rect 235826 708122 236062 708358
rect 236146 708122 236382 708358
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 240326 709402 240562 709638
rect 240646 709402 240882 709638
rect 240326 709082 240562 709318
rect 240646 709082 240882 709318
rect 240326 673718 240562 673954
rect 240646 673718 240882 673954
rect 240326 673398 240562 673634
rect 240646 673398 240882 673634
rect 244826 710362 245062 710598
rect 245146 710362 245382 710598
rect 244826 710042 245062 710278
rect 245146 710042 245382 710278
rect 244826 678218 245062 678454
rect 245146 678218 245382 678454
rect 244826 677898 245062 678134
rect 245146 677898 245382 678134
rect 249326 711322 249562 711558
rect 249646 711322 249882 711558
rect 249326 711002 249562 711238
rect 249646 711002 249882 711238
rect 249326 682718 249562 682954
rect 249646 682718 249882 682954
rect 249326 682398 249562 682634
rect 249646 682398 249882 682634
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 258326 705562 258562 705798
rect 258646 705562 258882 705798
rect 258326 705242 258562 705478
rect 258646 705242 258882 705478
rect 258326 691718 258562 691954
rect 258646 691718 258882 691954
rect 258326 691398 258562 691634
rect 258646 691398 258882 691634
rect 46826 660218 47062 660454
rect 47146 660218 47382 660454
rect 46826 659898 47062 660134
rect 47146 659898 47382 660134
rect 46826 624218 47062 624454
rect 47146 624218 47382 624454
rect 46826 623898 47062 624134
rect 47146 623898 47382 624134
rect 46826 588218 47062 588454
rect 47146 588218 47382 588454
rect 46826 587898 47062 588134
rect 47146 587898 47382 588134
rect 46826 552218 47062 552454
rect 47146 552218 47382 552454
rect 46826 551898 47062 552134
rect 47146 551898 47382 552134
rect 46826 516218 47062 516454
rect 47146 516218 47382 516454
rect 46826 515898 47062 516134
rect 47146 515898 47382 516134
rect 46826 480218 47062 480454
rect 47146 480218 47382 480454
rect 46826 479898 47062 480134
rect 47146 479898 47382 480134
rect 71610 655718 71846 655954
rect 71610 655398 71846 655634
rect 102330 655718 102566 655954
rect 102330 655398 102566 655634
rect 133050 655718 133286 655954
rect 133050 655398 133286 655634
rect 163770 655718 164006 655954
rect 163770 655398 164006 655634
rect 194490 655718 194726 655954
rect 194490 655398 194726 655634
rect 225210 655718 225446 655954
rect 225210 655398 225446 655634
rect 258326 655718 258562 655954
rect 258646 655718 258882 655954
rect 258326 655398 258562 655634
rect 258646 655398 258882 655634
rect 56250 651218 56486 651454
rect 56250 650898 56486 651134
rect 86970 651218 87206 651454
rect 86970 650898 87206 651134
rect 117690 651218 117926 651454
rect 117690 650898 117926 651134
rect 148410 651218 148646 651454
rect 148410 650898 148646 651134
rect 179130 651218 179366 651454
rect 179130 650898 179366 651134
rect 209850 651218 210086 651454
rect 209850 650898 210086 651134
rect 240570 651218 240806 651454
rect 240570 650898 240806 651134
rect 71610 619718 71846 619954
rect 71610 619398 71846 619634
rect 102330 619718 102566 619954
rect 102330 619398 102566 619634
rect 133050 619718 133286 619954
rect 133050 619398 133286 619634
rect 163770 619718 164006 619954
rect 163770 619398 164006 619634
rect 194490 619718 194726 619954
rect 194490 619398 194726 619634
rect 225210 619718 225446 619954
rect 225210 619398 225446 619634
rect 258326 619718 258562 619954
rect 258646 619718 258882 619954
rect 258326 619398 258562 619634
rect 258646 619398 258882 619634
rect 56250 615218 56486 615454
rect 56250 614898 56486 615134
rect 86970 615218 87206 615454
rect 86970 614898 87206 615134
rect 117690 615218 117926 615454
rect 117690 614898 117926 615134
rect 148410 615218 148646 615454
rect 148410 614898 148646 615134
rect 179130 615218 179366 615454
rect 179130 614898 179366 615134
rect 209850 615218 210086 615454
rect 209850 614898 210086 615134
rect 240570 615218 240806 615454
rect 240570 614898 240806 615134
rect 71610 583718 71846 583954
rect 71610 583398 71846 583634
rect 102330 583718 102566 583954
rect 102330 583398 102566 583634
rect 133050 583718 133286 583954
rect 133050 583398 133286 583634
rect 163770 583718 164006 583954
rect 163770 583398 164006 583634
rect 194490 583718 194726 583954
rect 194490 583398 194726 583634
rect 225210 583718 225446 583954
rect 225210 583398 225446 583634
rect 258326 583718 258562 583954
rect 258646 583718 258882 583954
rect 258326 583398 258562 583634
rect 258646 583398 258882 583634
rect 56250 579218 56486 579454
rect 56250 578898 56486 579134
rect 86970 579218 87206 579454
rect 86970 578898 87206 579134
rect 117690 579218 117926 579454
rect 117690 578898 117926 579134
rect 148410 579218 148646 579454
rect 148410 578898 148646 579134
rect 179130 579218 179366 579454
rect 179130 578898 179366 579134
rect 209850 579218 210086 579454
rect 209850 578898 210086 579134
rect 240570 579218 240806 579454
rect 240570 578898 240806 579134
rect 71610 547718 71846 547954
rect 71610 547398 71846 547634
rect 102330 547718 102566 547954
rect 102330 547398 102566 547634
rect 133050 547718 133286 547954
rect 133050 547398 133286 547634
rect 163770 547718 164006 547954
rect 163770 547398 164006 547634
rect 194490 547718 194726 547954
rect 194490 547398 194726 547634
rect 225210 547718 225446 547954
rect 225210 547398 225446 547634
rect 258326 547718 258562 547954
rect 258646 547718 258882 547954
rect 258326 547398 258562 547634
rect 258646 547398 258882 547634
rect 56250 543218 56486 543454
rect 56250 542898 56486 543134
rect 86970 543218 87206 543454
rect 86970 542898 87206 543134
rect 117690 543218 117926 543454
rect 117690 542898 117926 543134
rect 148410 543218 148646 543454
rect 148410 542898 148646 543134
rect 179130 543218 179366 543454
rect 179130 542898 179366 543134
rect 209850 543218 210086 543454
rect 209850 542898 210086 543134
rect 240570 543218 240806 543454
rect 240570 542898 240806 543134
rect 71610 511718 71846 511954
rect 71610 511398 71846 511634
rect 102330 511718 102566 511954
rect 102330 511398 102566 511634
rect 133050 511718 133286 511954
rect 133050 511398 133286 511634
rect 163770 511718 164006 511954
rect 163770 511398 164006 511634
rect 194490 511718 194726 511954
rect 194490 511398 194726 511634
rect 225210 511718 225446 511954
rect 225210 511398 225446 511634
rect 258326 511718 258562 511954
rect 258646 511718 258882 511954
rect 258326 511398 258562 511634
rect 258646 511398 258882 511634
rect 56250 507218 56486 507454
rect 56250 506898 56486 507134
rect 86970 507218 87206 507454
rect 86970 506898 87206 507134
rect 117690 507218 117926 507454
rect 117690 506898 117926 507134
rect 148410 507218 148646 507454
rect 148410 506898 148646 507134
rect 179130 507218 179366 507454
rect 179130 506898 179366 507134
rect 209850 507218 210086 507454
rect 209850 506898 210086 507134
rect 240570 507218 240806 507454
rect 240570 506898 240806 507134
rect 46826 444218 47062 444454
rect 47146 444218 47382 444454
rect 46826 443898 47062 444134
rect 47146 443898 47382 444134
rect 46826 408218 47062 408454
rect 47146 408218 47382 408454
rect 46826 407898 47062 408134
rect 47146 407898 47382 408134
rect 46826 372218 47062 372454
rect 47146 372218 47382 372454
rect 46826 371898 47062 372134
rect 47146 371898 47382 372134
rect 46826 336218 47062 336454
rect 47146 336218 47382 336454
rect 46826 335898 47062 336134
rect 47146 335898 47382 336134
rect 46826 300218 47062 300454
rect 47146 300218 47382 300454
rect 46826 299898 47062 300134
rect 47146 299898 47382 300134
rect 46826 264218 47062 264454
rect 47146 264218 47382 264454
rect 46826 263898 47062 264134
rect 47146 263898 47382 264134
rect 46826 228218 47062 228454
rect 47146 228218 47382 228454
rect 46826 227898 47062 228134
rect 47146 227898 47382 228134
rect 71610 475718 71846 475954
rect 71610 475398 71846 475634
rect 102330 475718 102566 475954
rect 102330 475398 102566 475634
rect 133050 475718 133286 475954
rect 133050 475398 133286 475634
rect 163770 475718 164006 475954
rect 163770 475398 164006 475634
rect 194490 475718 194726 475954
rect 194490 475398 194726 475634
rect 225210 475718 225446 475954
rect 225210 475398 225446 475634
rect 258326 475718 258562 475954
rect 258646 475718 258882 475954
rect 258326 475398 258562 475634
rect 258646 475398 258882 475634
rect 56250 471218 56486 471454
rect 56250 470898 56486 471134
rect 86970 471218 87206 471454
rect 86970 470898 87206 471134
rect 117690 471218 117926 471454
rect 117690 470898 117926 471134
rect 148410 471218 148646 471454
rect 148410 470898 148646 471134
rect 179130 471218 179366 471454
rect 179130 470898 179366 471134
rect 209850 471218 210086 471454
rect 209850 470898 210086 471134
rect 240570 471218 240806 471454
rect 240570 470898 240806 471134
rect 71610 439718 71846 439954
rect 71610 439398 71846 439634
rect 102330 439718 102566 439954
rect 102330 439398 102566 439634
rect 133050 439718 133286 439954
rect 133050 439398 133286 439634
rect 163770 439718 164006 439954
rect 163770 439398 164006 439634
rect 194490 439718 194726 439954
rect 194490 439398 194726 439634
rect 225210 439718 225446 439954
rect 225210 439398 225446 439634
rect 258326 439718 258562 439954
rect 258646 439718 258882 439954
rect 258326 439398 258562 439634
rect 258646 439398 258882 439634
rect 56250 435218 56486 435454
rect 56250 434898 56486 435134
rect 86970 435218 87206 435454
rect 86970 434898 87206 435134
rect 117690 435218 117926 435454
rect 117690 434898 117926 435134
rect 148410 435218 148646 435454
rect 148410 434898 148646 435134
rect 179130 435218 179366 435454
rect 179130 434898 179366 435134
rect 209850 435218 210086 435454
rect 209850 434898 210086 435134
rect 240570 435218 240806 435454
rect 240570 434898 240806 435134
rect 71610 403718 71846 403954
rect 71610 403398 71846 403634
rect 102330 403718 102566 403954
rect 102330 403398 102566 403634
rect 133050 403718 133286 403954
rect 133050 403398 133286 403634
rect 163770 403718 164006 403954
rect 163770 403398 164006 403634
rect 194490 403718 194726 403954
rect 194490 403398 194726 403634
rect 225210 403718 225446 403954
rect 225210 403398 225446 403634
rect 258326 403718 258562 403954
rect 258646 403718 258882 403954
rect 258326 403398 258562 403634
rect 258646 403398 258882 403634
rect 56250 399218 56486 399454
rect 56250 398898 56486 399134
rect 86970 399218 87206 399454
rect 86970 398898 87206 399134
rect 117690 399218 117926 399454
rect 117690 398898 117926 399134
rect 148410 399218 148646 399454
rect 148410 398898 148646 399134
rect 179130 399218 179366 399454
rect 179130 398898 179366 399134
rect 209850 399218 210086 399454
rect 209850 398898 210086 399134
rect 240570 399218 240806 399454
rect 240570 398898 240806 399134
rect 71610 367718 71846 367954
rect 71610 367398 71846 367634
rect 102330 367718 102566 367954
rect 102330 367398 102566 367634
rect 133050 367718 133286 367954
rect 133050 367398 133286 367634
rect 163770 367718 164006 367954
rect 163770 367398 164006 367634
rect 194490 367718 194726 367954
rect 194490 367398 194726 367634
rect 225210 367718 225446 367954
rect 225210 367398 225446 367634
rect 258326 367718 258562 367954
rect 258646 367718 258882 367954
rect 258326 367398 258562 367634
rect 258646 367398 258882 367634
rect 56250 363218 56486 363454
rect 56250 362898 56486 363134
rect 86970 363218 87206 363454
rect 86970 362898 87206 363134
rect 117690 363218 117926 363454
rect 117690 362898 117926 363134
rect 148410 363218 148646 363454
rect 148410 362898 148646 363134
rect 179130 363218 179366 363454
rect 179130 362898 179366 363134
rect 209850 363218 210086 363454
rect 209850 362898 210086 363134
rect 240570 363218 240806 363454
rect 240570 362898 240806 363134
rect 71610 331718 71846 331954
rect 71610 331398 71846 331634
rect 102330 331718 102566 331954
rect 102330 331398 102566 331634
rect 133050 331718 133286 331954
rect 133050 331398 133286 331634
rect 163770 331718 164006 331954
rect 163770 331398 164006 331634
rect 194490 331718 194726 331954
rect 194490 331398 194726 331634
rect 225210 331718 225446 331954
rect 225210 331398 225446 331634
rect 258326 331718 258562 331954
rect 258646 331718 258882 331954
rect 258326 331398 258562 331634
rect 258646 331398 258882 331634
rect 56250 327218 56486 327454
rect 56250 326898 56486 327134
rect 86970 327218 87206 327454
rect 86970 326898 87206 327134
rect 117690 327218 117926 327454
rect 117690 326898 117926 327134
rect 148410 327218 148646 327454
rect 148410 326898 148646 327134
rect 179130 327218 179366 327454
rect 179130 326898 179366 327134
rect 209850 327218 210086 327454
rect 209850 326898 210086 327134
rect 240570 327218 240806 327454
rect 240570 326898 240806 327134
rect 71610 295718 71846 295954
rect 71610 295398 71846 295634
rect 102330 295718 102566 295954
rect 102330 295398 102566 295634
rect 133050 295718 133286 295954
rect 133050 295398 133286 295634
rect 163770 295718 164006 295954
rect 163770 295398 164006 295634
rect 194490 295718 194726 295954
rect 194490 295398 194726 295634
rect 225210 295718 225446 295954
rect 225210 295398 225446 295634
rect 258326 295718 258562 295954
rect 258646 295718 258882 295954
rect 258326 295398 258562 295634
rect 258646 295398 258882 295634
rect 56250 291218 56486 291454
rect 56250 290898 56486 291134
rect 86970 291218 87206 291454
rect 86970 290898 87206 291134
rect 117690 291218 117926 291454
rect 117690 290898 117926 291134
rect 148410 291218 148646 291454
rect 148410 290898 148646 291134
rect 179130 291218 179366 291454
rect 179130 290898 179366 291134
rect 209850 291218 210086 291454
rect 209850 290898 210086 291134
rect 240570 291218 240806 291454
rect 240570 290898 240806 291134
rect 51326 268718 51562 268954
rect 51646 268718 51882 268954
rect 51326 268398 51562 268634
rect 51646 268398 51882 268634
rect 51326 232718 51562 232954
rect 51646 232718 51882 232954
rect 51326 232398 51562 232634
rect 51646 232398 51882 232634
rect 46826 192218 47062 192454
rect 47146 192218 47382 192454
rect 46826 191898 47062 192134
rect 47146 191898 47382 192134
rect 46826 156218 47062 156454
rect 47146 156218 47382 156454
rect 46826 155898 47062 156134
rect 47146 155898 47382 156134
rect 46826 120218 47062 120454
rect 47146 120218 47382 120454
rect 46826 119898 47062 120134
rect 47146 119898 47382 120134
rect 46826 84218 47062 84454
rect 47146 84218 47382 84454
rect 46826 83898 47062 84134
rect 47146 83898 47382 84134
rect 46826 48218 47062 48454
rect 47146 48218 47382 48454
rect 46826 47898 47062 48134
rect 47146 47898 47382 48134
rect 46826 12218 47062 12454
rect 47146 12218 47382 12454
rect 46826 11898 47062 12134
rect 47146 11898 47382 12134
rect 46826 -2502 47062 -2266
rect 47146 -2502 47382 -2266
rect 46826 -2822 47062 -2586
rect 47146 -2822 47382 -2586
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 60326 277718 60562 277954
rect 60646 277718 60882 277954
rect 60326 277398 60562 277634
rect 60646 277398 60882 277634
rect 60326 241718 60562 241954
rect 60646 241718 60882 241954
rect 60326 241398 60562 241634
rect 60646 241398 60882 241634
rect 51326 196718 51562 196954
rect 51646 196718 51882 196954
rect 51326 196398 51562 196634
rect 51646 196398 51882 196634
rect 51326 160718 51562 160954
rect 51646 160718 51882 160954
rect 51326 160398 51562 160634
rect 51646 160398 51882 160634
rect 78326 259718 78562 259954
rect 78646 259718 78882 259954
rect 78326 259398 78562 259634
rect 78646 259398 78882 259634
rect 78326 223718 78562 223954
rect 78646 223718 78882 223954
rect 78326 223398 78562 223634
rect 78646 223398 78882 223634
rect 82826 264218 83062 264454
rect 83146 264218 83382 264454
rect 82826 263898 83062 264134
rect 83146 263898 83382 264134
rect 82826 228218 83062 228454
rect 83146 228218 83382 228454
rect 82826 227898 83062 228134
rect 83146 227898 83382 228134
rect 87326 268718 87562 268954
rect 87646 268718 87882 268954
rect 87326 268398 87562 268634
rect 87646 268398 87882 268634
rect 87326 232718 87562 232954
rect 87646 232718 87882 232954
rect 87326 232398 87562 232634
rect 87646 232398 87882 232634
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 96326 277718 96562 277954
rect 96646 277718 96882 277954
rect 96326 277398 96562 277634
rect 96646 277398 96882 277634
rect 96326 241718 96562 241954
rect 96646 241718 96882 241954
rect 96326 241398 96562 241634
rect 96646 241398 96882 241634
rect 114326 259718 114562 259954
rect 114646 259718 114882 259954
rect 114326 259398 114562 259634
rect 114646 259398 114882 259634
rect 114326 223718 114562 223954
rect 114646 223718 114882 223954
rect 114326 223398 114562 223634
rect 114646 223398 114882 223634
rect 118826 264218 119062 264454
rect 119146 264218 119382 264454
rect 118826 263898 119062 264134
rect 119146 263898 119382 264134
rect 118826 228218 119062 228454
rect 119146 228218 119382 228454
rect 118826 227898 119062 228134
rect 119146 227898 119382 228134
rect 123326 268718 123562 268954
rect 123646 268718 123882 268954
rect 123326 268398 123562 268634
rect 123646 268398 123882 268634
rect 123326 232718 123562 232954
rect 123646 232718 123882 232954
rect 123326 232398 123562 232634
rect 123646 232398 123882 232634
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 132326 277718 132562 277954
rect 132646 277718 132882 277954
rect 132326 277398 132562 277634
rect 132646 277398 132882 277634
rect 132326 241718 132562 241954
rect 132646 241718 132882 241954
rect 132326 241398 132562 241634
rect 132646 241398 132882 241634
rect 150326 259718 150562 259954
rect 150646 259718 150882 259954
rect 150326 259398 150562 259634
rect 150646 259398 150882 259634
rect 150326 223718 150562 223954
rect 150646 223718 150882 223954
rect 150326 223398 150562 223634
rect 150646 223398 150882 223634
rect 154826 264218 155062 264454
rect 155146 264218 155382 264454
rect 154826 263898 155062 264134
rect 155146 263898 155382 264134
rect 154826 228218 155062 228454
rect 155146 228218 155382 228454
rect 154826 227898 155062 228134
rect 155146 227898 155382 228134
rect 159326 268718 159562 268954
rect 159646 268718 159882 268954
rect 159326 268398 159562 268634
rect 159646 268398 159882 268634
rect 159326 232718 159562 232954
rect 159646 232718 159882 232954
rect 159326 232398 159562 232634
rect 159646 232398 159882 232634
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 168326 277718 168562 277954
rect 168646 277718 168882 277954
rect 168326 277398 168562 277634
rect 168646 277398 168882 277634
rect 168326 241718 168562 241954
rect 168646 241718 168882 241954
rect 168326 241398 168562 241634
rect 168646 241398 168882 241634
rect 186326 259718 186562 259954
rect 186646 259718 186882 259954
rect 186326 259398 186562 259634
rect 186646 259398 186882 259634
rect 186326 223718 186562 223954
rect 186646 223718 186882 223954
rect 186326 223398 186562 223634
rect 186646 223398 186882 223634
rect 190826 264218 191062 264454
rect 191146 264218 191382 264454
rect 190826 263898 191062 264134
rect 191146 263898 191382 264134
rect 190826 228218 191062 228454
rect 191146 228218 191382 228454
rect 190826 227898 191062 228134
rect 191146 227898 191382 228134
rect 195326 268718 195562 268954
rect 195646 268718 195882 268954
rect 195326 268398 195562 268634
rect 195646 268398 195882 268634
rect 195326 232718 195562 232954
rect 195646 232718 195882 232954
rect 195326 232398 195562 232634
rect 195646 232398 195882 232634
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 204326 277718 204562 277954
rect 204646 277718 204882 277954
rect 204326 277398 204562 277634
rect 204646 277398 204882 277634
rect 204326 241718 204562 241954
rect 204646 241718 204882 241954
rect 204326 241398 204562 241634
rect 204646 241398 204882 241634
rect 222326 259718 222562 259954
rect 222646 259718 222882 259954
rect 222326 259398 222562 259634
rect 222646 259398 222882 259634
rect 222326 223718 222562 223954
rect 222646 223718 222882 223954
rect 222326 223398 222562 223634
rect 222646 223398 222882 223634
rect 226826 264218 227062 264454
rect 227146 264218 227382 264454
rect 226826 263898 227062 264134
rect 227146 263898 227382 264134
rect 226826 228218 227062 228454
rect 227146 228218 227382 228454
rect 226826 227898 227062 228134
rect 227146 227898 227382 228134
rect 226826 192218 227062 192454
rect 227146 192218 227382 192454
rect 226826 191898 227062 192134
rect 227146 191898 227382 192134
rect 79610 187718 79846 187954
rect 79610 187398 79846 187634
rect 110330 187718 110566 187954
rect 110330 187398 110566 187634
rect 141050 187718 141286 187954
rect 141050 187398 141286 187634
rect 171770 187718 172006 187954
rect 171770 187398 172006 187634
rect 202490 187718 202726 187954
rect 202490 187398 202726 187634
rect 64250 183218 64486 183454
rect 64250 182898 64486 183134
rect 94970 183218 95206 183454
rect 94970 182898 95206 183134
rect 125690 183218 125926 183454
rect 125690 182898 125926 183134
rect 156410 183218 156646 183454
rect 156410 182898 156646 183134
rect 187130 183218 187366 183454
rect 187130 182898 187366 183134
rect 217850 183218 218086 183454
rect 217850 182898 218086 183134
rect 226826 156218 227062 156454
rect 227146 156218 227382 156454
rect 226826 155898 227062 156134
rect 227146 155898 227382 156134
rect 79610 151718 79846 151954
rect 79610 151398 79846 151634
rect 110330 151718 110566 151954
rect 110330 151398 110566 151634
rect 141050 151718 141286 151954
rect 141050 151398 141286 151634
rect 171770 151718 172006 151954
rect 171770 151398 172006 151634
rect 202490 151718 202726 151954
rect 202490 151398 202726 151634
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 51326 124718 51562 124954
rect 51646 124718 51882 124954
rect 51326 124398 51562 124634
rect 51646 124398 51882 124634
rect 226826 120218 227062 120454
rect 227146 120218 227382 120454
rect 226826 119898 227062 120134
rect 227146 119898 227382 120134
rect 79610 115718 79846 115954
rect 79610 115398 79846 115634
rect 110330 115718 110566 115954
rect 110330 115398 110566 115634
rect 141050 115718 141286 115954
rect 141050 115398 141286 115634
rect 171770 115718 172006 115954
rect 171770 115398 172006 115634
rect 202490 115718 202726 115954
rect 202490 115398 202726 115634
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 51326 88718 51562 88954
rect 51646 88718 51882 88954
rect 51326 88398 51562 88634
rect 51646 88398 51882 88634
rect 226826 84218 227062 84454
rect 227146 84218 227382 84454
rect 226826 83898 227062 84134
rect 227146 83898 227382 84134
rect 79610 79718 79846 79954
rect 79610 79398 79846 79634
rect 110330 79718 110566 79954
rect 110330 79398 110566 79634
rect 141050 79718 141286 79954
rect 141050 79398 141286 79634
rect 171770 79718 172006 79954
rect 171770 79398 172006 79634
rect 202490 79718 202726 79954
rect 202490 79398 202726 79634
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 51326 52718 51562 52954
rect 51646 52718 51882 52954
rect 51326 52398 51562 52634
rect 51646 52398 51882 52634
rect 51326 16718 51562 16954
rect 51646 16718 51882 16954
rect 51326 16398 51562 16634
rect 51646 16398 51882 16634
rect 51326 -3462 51562 -3226
rect 51646 -3462 51882 -3226
rect 51326 -3782 51562 -3546
rect 51646 -3782 51882 -3546
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -4422 56062 -4186
rect 56146 -4422 56382 -4186
rect 55826 -4742 56062 -4506
rect 56146 -4742 56382 -4506
rect 60326 25718 60562 25954
rect 60646 25718 60882 25954
rect 60326 25398 60562 25634
rect 60646 25398 60882 25634
rect 60326 -5382 60562 -5146
rect 60646 -5382 60882 -5146
rect 60326 -5702 60562 -5466
rect 60646 -5702 60882 -5466
rect 64826 30218 65062 30454
rect 65146 30218 65382 30454
rect 64826 29898 65062 30134
rect 65146 29898 65382 30134
rect 64826 -6342 65062 -6106
rect 65146 -6342 65382 -6106
rect 64826 -6662 65062 -6426
rect 65146 -6662 65382 -6426
rect 69326 34718 69562 34954
rect 69646 34718 69882 34954
rect 69326 34398 69562 34634
rect 69646 34398 69882 34634
rect 69326 -7302 69562 -7066
rect 69646 -7302 69882 -7066
rect 69326 -7622 69562 -7386
rect 69646 -7622 69882 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 78326 43718 78562 43954
rect 78646 43718 78882 43954
rect 78326 43398 78562 43634
rect 78646 43398 78882 43634
rect 78326 7718 78562 7954
rect 78646 7718 78882 7954
rect 78326 7398 78562 7634
rect 78646 7398 78882 7634
rect 78326 -1542 78562 -1306
rect 78646 -1542 78882 -1306
rect 78326 -1862 78562 -1626
rect 78646 -1862 78882 -1626
rect 82826 48218 83062 48454
rect 83146 48218 83382 48454
rect 82826 47898 83062 48134
rect 83146 47898 83382 48134
rect 82826 12218 83062 12454
rect 83146 12218 83382 12454
rect 82826 11898 83062 12134
rect 83146 11898 83382 12134
rect 82826 -2502 83062 -2266
rect 83146 -2502 83382 -2266
rect 82826 -2822 83062 -2586
rect 83146 -2822 83382 -2586
rect 87326 52718 87562 52954
rect 87646 52718 87882 52954
rect 87326 52398 87562 52634
rect 87646 52398 87882 52634
rect 87326 16718 87562 16954
rect 87646 16718 87882 16954
rect 87326 16398 87562 16634
rect 87646 16398 87882 16634
rect 87326 -3462 87562 -3226
rect 87646 -3462 87882 -3226
rect 87326 -3782 87562 -3546
rect 87646 -3782 87882 -3546
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -4422 92062 -4186
rect 92146 -4422 92382 -4186
rect 91826 -4742 92062 -4506
rect 92146 -4742 92382 -4506
rect 96326 25718 96562 25954
rect 96646 25718 96882 25954
rect 96326 25398 96562 25634
rect 96646 25398 96882 25634
rect 96326 -5382 96562 -5146
rect 96646 -5382 96882 -5146
rect 96326 -5702 96562 -5466
rect 96646 -5702 96882 -5466
rect 100826 30218 101062 30454
rect 101146 30218 101382 30454
rect 100826 29898 101062 30134
rect 101146 29898 101382 30134
rect 100826 -6342 101062 -6106
rect 101146 -6342 101382 -6106
rect 100826 -6662 101062 -6426
rect 101146 -6662 101382 -6426
rect 105326 34718 105562 34954
rect 105646 34718 105882 34954
rect 105326 34398 105562 34634
rect 105646 34398 105882 34634
rect 105326 -7302 105562 -7066
rect 105646 -7302 105882 -7066
rect 105326 -7622 105562 -7386
rect 105646 -7622 105882 -7386
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 114326 43718 114562 43954
rect 114646 43718 114882 43954
rect 114326 43398 114562 43634
rect 114646 43398 114882 43634
rect 114326 7718 114562 7954
rect 114646 7718 114882 7954
rect 114326 7398 114562 7634
rect 114646 7398 114882 7634
rect 114326 -1542 114562 -1306
rect 114646 -1542 114882 -1306
rect 114326 -1862 114562 -1626
rect 114646 -1862 114882 -1626
rect 118826 48218 119062 48454
rect 119146 48218 119382 48454
rect 118826 47898 119062 48134
rect 119146 47898 119382 48134
rect 118826 12218 119062 12454
rect 119146 12218 119382 12454
rect 118826 11898 119062 12134
rect 119146 11898 119382 12134
rect 118826 -2502 119062 -2266
rect 119146 -2502 119382 -2266
rect 118826 -2822 119062 -2586
rect 119146 -2822 119382 -2586
rect 123326 52718 123562 52954
rect 123646 52718 123882 52954
rect 123326 52398 123562 52634
rect 123646 52398 123882 52634
rect 123326 16718 123562 16954
rect 123646 16718 123882 16954
rect 123326 16398 123562 16634
rect 123646 16398 123882 16634
rect 123326 -3462 123562 -3226
rect 123646 -3462 123882 -3226
rect 123326 -3782 123562 -3546
rect 123646 -3782 123882 -3546
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -4422 128062 -4186
rect 128146 -4422 128382 -4186
rect 127826 -4742 128062 -4506
rect 128146 -4742 128382 -4506
rect 132326 25718 132562 25954
rect 132646 25718 132882 25954
rect 132326 25398 132562 25634
rect 132646 25398 132882 25634
rect 132326 -5382 132562 -5146
rect 132646 -5382 132882 -5146
rect 132326 -5702 132562 -5466
rect 132646 -5702 132882 -5466
rect 136826 30218 137062 30454
rect 137146 30218 137382 30454
rect 136826 29898 137062 30134
rect 137146 29898 137382 30134
rect 136826 -6342 137062 -6106
rect 137146 -6342 137382 -6106
rect 136826 -6662 137062 -6426
rect 137146 -6662 137382 -6426
rect 141326 34718 141562 34954
rect 141646 34718 141882 34954
rect 141326 34398 141562 34634
rect 141646 34398 141882 34634
rect 141326 -7302 141562 -7066
rect 141646 -7302 141882 -7066
rect 141326 -7622 141562 -7386
rect 141646 -7622 141882 -7386
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 150326 43718 150562 43954
rect 150646 43718 150882 43954
rect 150326 43398 150562 43634
rect 150646 43398 150882 43634
rect 150326 7718 150562 7954
rect 150646 7718 150882 7954
rect 150326 7398 150562 7634
rect 150646 7398 150882 7634
rect 150326 -1542 150562 -1306
rect 150646 -1542 150882 -1306
rect 150326 -1862 150562 -1626
rect 150646 -1862 150882 -1626
rect 154826 48218 155062 48454
rect 155146 48218 155382 48454
rect 154826 47898 155062 48134
rect 155146 47898 155382 48134
rect 154826 12218 155062 12454
rect 155146 12218 155382 12454
rect 154826 11898 155062 12134
rect 155146 11898 155382 12134
rect 154826 -2502 155062 -2266
rect 155146 -2502 155382 -2266
rect 154826 -2822 155062 -2586
rect 155146 -2822 155382 -2586
rect 159326 52718 159562 52954
rect 159646 52718 159882 52954
rect 159326 52398 159562 52634
rect 159646 52398 159882 52634
rect 159326 16718 159562 16954
rect 159646 16718 159882 16954
rect 159326 16398 159562 16634
rect 159646 16398 159882 16634
rect 159326 -3462 159562 -3226
rect 159646 -3462 159882 -3226
rect 159326 -3782 159562 -3546
rect 159646 -3782 159882 -3546
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -4422 164062 -4186
rect 164146 -4422 164382 -4186
rect 163826 -4742 164062 -4506
rect 164146 -4742 164382 -4506
rect 168326 25718 168562 25954
rect 168646 25718 168882 25954
rect 168326 25398 168562 25634
rect 168646 25398 168882 25634
rect 168326 -5382 168562 -5146
rect 168646 -5382 168882 -5146
rect 168326 -5702 168562 -5466
rect 168646 -5702 168882 -5466
rect 172826 30218 173062 30454
rect 173146 30218 173382 30454
rect 172826 29898 173062 30134
rect 173146 29898 173382 30134
rect 172826 -6342 173062 -6106
rect 173146 -6342 173382 -6106
rect 172826 -6662 173062 -6426
rect 173146 -6662 173382 -6426
rect 177326 34718 177562 34954
rect 177646 34718 177882 34954
rect 177326 34398 177562 34634
rect 177646 34398 177882 34634
rect 177326 -7302 177562 -7066
rect 177646 -7302 177882 -7066
rect 177326 -7622 177562 -7386
rect 177646 -7622 177882 -7386
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 186326 43718 186562 43954
rect 186646 43718 186882 43954
rect 186326 43398 186562 43634
rect 186646 43398 186882 43634
rect 186326 7718 186562 7954
rect 186646 7718 186882 7954
rect 186326 7398 186562 7634
rect 186646 7398 186882 7634
rect 186326 -1542 186562 -1306
rect 186646 -1542 186882 -1306
rect 186326 -1862 186562 -1626
rect 186646 -1862 186882 -1626
rect 190826 48218 191062 48454
rect 191146 48218 191382 48454
rect 190826 47898 191062 48134
rect 191146 47898 191382 48134
rect 190826 12218 191062 12454
rect 191146 12218 191382 12454
rect 190826 11898 191062 12134
rect 191146 11898 191382 12134
rect 190826 -2502 191062 -2266
rect 191146 -2502 191382 -2266
rect 190826 -2822 191062 -2586
rect 191146 -2822 191382 -2586
rect 195326 52718 195562 52954
rect 195646 52718 195882 52954
rect 195326 52398 195562 52634
rect 195646 52398 195882 52634
rect 195326 16718 195562 16954
rect 195646 16718 195882 16954
rect 195326 16398 195562 16634
rect 195646 16398 195882 16634
rect 195326 -3462 195562 -3226
rect 195646 -3462 195882 -3226
rect 195326 -3782 195562 -3546
rect 195646 -3782 195882 -3546
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -4422 200062 -4186
rect 200146 -4422 200382 -4186
rect 199826 -4742 200062 -4506
rect 200146 -4742 200382 -4506
rect 204326 25718 204562 25954
rect 204646 25718 204882 25954
rect 204326 25398 204562 25634
rect 204646 25398 204882 25634
rect 204326 -5382 204562 -5146
rect 204646 -5382 204882 -5146
rect 204326 -5702 204562 -5466
rect 204646 -5702 204882 -5466
rect 208826 30218 209062 30454
rect 209146 30218 209382 30454
rect 208826 29898 209062 30134
rect 209146 29898 209382 30134
rect 208826 -6342 209062 -6106
rect 209146 -6342 209382 -6106
rect 208826 -6662 209062 -6426
rect 209146 -6662 209382 -6426
rect 213326 34718 213562 34954
rect 213646 34718 213882 34954
rect 213326 34398 213562 34634
rect 213646 34398 213882 34634
rect 213326 -7302 213562 -7066
rect 213646 -7302 213882 -7066
rect 213326 -7622 213562 -7386
rect 213646 -7622 213882 -7386
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 222326 43718 222562 43954
rect 222646 43718 222882 43954
rect 222326 43398 222562 43634
rect 222646 43398 222882 43634
rect 222326 7718 222562 7954
rect 222646 7718 222882 7954
rect 222326 7398 222562 7634
rect 222646 7398 222882 7634
rect 222326 -1542 222562 -1306
rect 222646 -1542 222882 -1306
rect 222326 -1862 222562 -1626
rect 222646 -1862 222882 -1626
rect 226826 48218 227062 48454
rect 227146 48218 227382 48454
rect 226826 47898 227062 48134
rect 227146 47898 227382 48134
rect 226826 12218 227062 12454
rect 227146 12218 227382 12454
rect 226826 11898 227062 12134
rect 227146 11898 227382 12134
rect 226826 -2502 227062 -2266
rect 227146 -2502 227382 -2266
rect 226826 -2822 227062 -2586
rect 227146 -2822 227382 -2586
rect 231326 268718 231562 268954
rect 231646 268718 231882 268954
rect 231326 268398 231562 268634
rect 231646 268398 231882 268634
rect 231326 232718 231562 232954
rect 231646 232718 231882 232954
rect 231326 232398 231562 232634
rect 231646 232398 231882 232634
rect 231326 196718 231562 196954
rect 231646 196718 231882 196954
rect 231326 196398 231562 196634
rect 231646 196398 231882 196634
rect 231326 160718 231562 160954
rect 231646 160718 231882 160954
rect 231326 160398 231562 160634
rect 231646 160398 231882 160634
rect 231326 124718 231562 124954
rect 231646 124718 231882 124954
rect 231326 124398 231562 124634
rect 231646 124398 231882 124634
rect 231326 88718 231562 88954
rect 231646 88718 231882 88954
rect 231326 88398 231562 88634
rect 231646 88398 231882 88634
rect 231326 52718 231562 52954
rect 231646 52718 231882 52954
rect 231326 52398 231562 52634
rect 231646 52398 231882 52634
rect 231326 16718 231562 16954
rect 231646 16718 231882 16954
rect 231326 16398 231562 16634
rect 231646 16398 231882 16634
rect 231326 -3462 231562 -3226
rect 231646 -3462 231882 -3226
rect 231326 -3782 231562 -3546
rect 231646 -3782 231882 -3546
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -4422 236062 -4186
rect 236146 -4422 236382 -4186
rect 235826 -4742 236062 -4506
rect 236146 -4742 236382 -4506
rect 240326 277718 240562 277954
rect 240646 277718 240882 277954
rect 240326 277398 240562 277634
rect 240646 277398 240882 277634
rect 240326 241718 240562 241954
rect 240646 241718 240882 241954
rect 240326 241398 240562 241634
rect 240646 241398 240882 241634
rect 240326 205718 240562 205954
rect 240646 205718 240882 205954
rect 240326 205398 240562 205634
rect 240646 205398 240882 205634
rect 240326 169718 240562 169954
rect 240646 169718 240882 169954
rect 240326 169398 240562 169634
rect 240646 169398 240882 169634
rect 240326 133718 240562 133954
rect 240646 133718 240882 133954
rect 240326 133398 240562 133634
rect 240646 133398 240882 133634
rect 240326 97718 240562 97954
rect 240646 97718 240882 97954
rect 240326 97398 240562 97634
rect 240646 97398 240882 97634
rect 240326 61718 240562 61954
rect 240646 61718 240882 61954
rect 240326 61398 240562 61634
rect 240646 61398 240882 61634
rect 240326 25718 240562 25954
rect 240646 25718 240882 25954
rect 240326 25398 240562 25634
rect 240646 25398 240882 25634
rect 240326 -5382 240562 -5146
rect 240646 -5382 240882 -5146
rect 240326 -5702 240562 -5466
rect 240646 -5702 240882 -5466
rect 244826 246218 245062 246454
rect 245146 246218 245382 246454
rect 244826 245898 245062 246134
rect 245146 245898 245382 246134
rect 244826 210218 245062 210454
rect 245146 210218 245382 210454
rect 244826 209898 245062 210134
rect 245146 209898 245382 210134
rect 244826 174218 245062 174454
rect 245146 174218 245382 174454
rect 244826 173898 245062 174134
rect 245146 173898 245382 174134
rect 244826 138218 245062 138454
rect 245146 138218 245382 138454
rect 244826 137898 245062 138134
rect 245146 137898 245382 138134
rect 244826 102218 245062 102454
rect 245146 102218 245382 102454
rect 244826 101898 245062 102134
rect 245146 101898 245382 102134
rect 244826 66218 245062 66454
rect 245146 66218 245382 66454
rect 244826 65898 245062 66134
rect 245146 65898 245382 66134
rect 244826 30218 245062 30454
rect 245146 30218 245382 30454
rect 244826 29898 245062 30134
rect 245146 29898 245382 30134
rect 244826 -6342 245062 -6106
rect 245146 -6342 245382 -6106
rect 244826 -6662 245062 -6426
rect 245146 -6662 245382 -6426
rect 249326 250718 249562 250954
rect 249646 250718 249882 250954
rect 249326 250398 249562 250634
rect 249646 250398 249882 250634
rect 249326 214718 249562 214954
rect 249646 214718 249882 214954
rect 249326 214398 249562 214634
rect 249646 214398 249882 214634
rect 249326 178718 249562 178954
rect 249646 178718 249882 178954
rect 249326 178398 249562 178634
rect 249646 178398 249882 178634
rect 249326 142718 249562 142954
rect 249646 142718 249882 142954
rect 249326 142398 249562 142634
rect 249646 142398 249882 142634
rect 249326 106718 249562 106954
rect 249646 106718 249882 106954
rect 249326 106398 249562 106634
rect 249646 106398 249882 106634
rect 249326 70718 249562 70954
rect 249646 70718 249882 70954
rect 249326 70398 249562 70634
rect 249646 70398 249882 70634
rect 249326 34718 249562 34954
rect 249646 34718 249882 34954
rect 249326 34398 249562 34634
rect 249646 34398 249882 34634
rect 249326 -7302 249562 -7066
rect 249646 -7302 249882 -7066
rect 249326 -7622 249562 -7386
rect 249646 -7622 249882 -7386
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 258326 259718 258562 259954
rect 258646 259718 258882 259954
rect 258326 259398 258562 259634
rect 258646 259398 258882 259634
rect 258326 223718 258562 223954
rect 258646 223718 258882 223954
rect 258326 223398 258562 223634
rect 258646 223398 258882 223634
rect 258326 187718 258562 187954
rect 258646 187718 258882 187954
rect 258326 187398 258562 187634
rect 258646 187398 258882 187634
rect 258326 151718 258562 151954
rect 258646 151718 258882 151954
rect 258326 151398 258562 151634
rect 258646 151398 258882 151634
rect 258326 115718 258562 115954
rect 258646 115718 258882 115954
rect 258326 115398 258562 115634
rect 258646 115398 258882 115634
rect 258326 79718 258562 79954
rect 258646 79718 258882 79954
rect 258326 79398 258562 79634
rect 258646 79398 258882 79634
rect 258326 43718 258562 43954
rect 258646 43718 258882 43954
rect 258326 43398 258562 43634
rect 258646 43398 258882 43634
rect 258326 7718 258562 7954
rect 258646 7718 258882 7954
rect 258326 7398 258562 7634
rect 258646 7398 258882 7634
rect 258326 -1542 258562 -1306
rect 258646 -1542 258882 -1306
rect 258326 -1862 258562 -1626
rect 258646 -1862 258882 -1626
rect 262826 706522 263062 706758
rect 263146 706522 263382 706758
rect 262826 706202 263062 706438
rect 263146 706202 263382 706438
rect 262826 696218 263062 696454
rect 263146 696218 263382 696454
rect 262826 695898 263062 696134
rect 263146 695898 263382 696134
rect 262826 660218 263062 660454
rect 263146 660218 263382 660454
rect 262826 659898 263062 660134
rect 263146 659898 263382 660134
rect 262826 624218 263062 624454
rect 263146 624218 263382 624454
rect 262826 623898 263062 624134
rect 263146 623898 263382 624134
rect 262826 588218 263062 588454
rect 263146 588218 263382 588454
rect 262826 587898 263062 588134
rect 263146 587898 263382 588134
rect 262826 552218 263062 552454
rect 263146 552218 263382 552454
rect 262826 551898 263062 552134
rect 263146 551898 263382 552134
rect 262826 516218 263062 516454
rect 263146 516218 263382 516454
rect 262826 515898 263062 516134
rect 263146 515898 263382 516134
rect 262826 480218 263062 480454
rect 263146 480218 263382 480454
rect 262826 479898 263062 480134
rect 263146 479898 263382 480134
rect 262826 444218 263062 444454
rect 263146 444218 263382 444454
rect 262826 443898 263062 444134
rect 263146 443898 263382 444134
rect 262826 408218 263062 408454
rect 263146 408218 263382 408454
rect 262826 407898 263062 408134
rect 263146 407898 263382 408134
rect 262826 372218 263062 372454
rect 263146 372218 263382 372454
rect 262826 371898 263062 372134
rect 263146 371898 263382 372134
rect 262826 336218 263062 336454
rect 263146 336218 263382 336454
rect 262826 335898 263062 336134
rect 263146 335898 263382 336134
rect 262826 300218 263062 300454
rect 263146 300218 263382 300454
rect 262826 299898 263062 300134
rect 263146 299898 263382 300134
rect 262826 264218 263062 264454
rect 263146 264218 263382 264454
rect 262826 263898 263062 264134
rect 263146 263898 263382 264134
rect 262826 228218 263062 228454
rect 263146 228218 263382 228454
rect 262826 227898 263062 228134
rect 263146 227898 263382 228134
rect 262826 192218 263062 192454
rect 263146 192218 263382 192454
rect 262826 191898 263062 192134
rect 263146 191898 263382 192134
rect 262826 156218 263062 156454
rect 263146 156218 263382 156454
rect 262826 155898 263062 156134
rect 263146 155898 263382 156134
rect 262826 120218 263062 120454
rect 263146 120218 263382 120454
rect 262826 119898 263062 120134
rect 263146 119898 263382 120134
rect 262826 84218 263062 84454
rect 263146 84218 263382 84454
rect 262826 83898 263062 84134
rect 263146 83898 263382 84134
rect 262826 48218 263062 48454
rect 263146 48218 263382 48454
rect 262826 47898 263062 48134
rect 263146 47898 263382 48134
rect 262826 12218 263062 12454
rect 263146 12218 263382 12454
rect 262826 11898 263062 12134
rect 263146 11898 263382 12134
rect 262826 -2502 263062 -2266
rect 263146 -2502 263382 -2266
rect 262826 -2822 263062 -2586
rect 263146 -2822 263382 -2586
rect 267326 707482 267562 707718
rect 267646 707482 267882 707718
rect 267326 707162 267562 707398
rect 267646 707162 267882 707398
rect 267326 700718 267562 700954
rect 267646 700718 267882 700954
rect 267326 700398 267562 700634
rect 267646 700398 267882 700634
rect 267326 664718 267562 664954
rect 267646 664718 267882 664954
rect 267326 664398 267562 664634
rect 267646 664398 267882 664634
rect 267326 628718 267562 628954
rect 267646 628718 267882 628954
rect 267326 628398 267562 628634
rect 267646 628398 267882 628634
rect 267326 592718 267562 592954
rect 267646 592718 267882 592954
rect 267326 592398 267562 592634
rect 267646 592398 267882 592634
rect 267326 556718 267562 556954
rect 267646 556718 267882 556954
rect 267326 556398 267562 556634
rect 267646 556398 267882 556634
rect 267326 520718 267562 520954
rect 267646 520718 267882 520954
rect 267326 520398 267562 520634
rect 267646 520398 267882 520634
rect 267326 484718 267562 484954
rect 267646 484718 267882 484954
rect 267326 484398 267562 484634
rect 267646 484398 267882 484634
rect 267326 448718 267562 448954
rect 267646 448718 267882 448954
rect 267326 448398 267562 448634
rect 267646 448398 267882 448634
rect 267326 412718 267562 412954
rect 267646 412718 267882 412954
rect 267326 412398 267562 412634
rect 267646 412398 267882 412634
rect 267326 376718 267562 376954
rect 267646 376718 267882 376954
rect 267326 376398 267562 376634
rect 267646 376398 267882 376634
rect 267326 340718 267562 340954
rect 267646 340718 267882 340954
rect 267326 340398 267562 340634
rect 267646 340398 267882 340634
rect 267326 304718 267562 304954
rect 267646 304718 267882 304954
rect 267326 304398 267562 304634
rect 267646 304398 267882 304634
rect 267326 268718 267562 268954
rect 267646 268718 267882 268954
rect 267326 268398 267562 268634
rect 267646 268398 267882 268634
rect 267326 232718 267562 232954
rect 267646 232718 267882 232954
rect 267326 232398 267562 232634
rect 267646 232398 267882 232634
rect 267326 196718 267562 196954
rect 267646 196718 267882 196954
rect 267326 196398 267562 196634
rect 267646 196398 267882 196634
rect 267326 160718 267562 160954
rect 267646 160718 267882 160954
rect 267326 160398 267562 160634
rect 267646 160398 267882 160634
rect 267326 124718 267562 124954
rect 267646 124718 267882 124954
rect 267326 124398 267562 124634
rect 267646 124398 267882 124634
rect 267326 88718 267562 88954
rect 267646 88718 267882 88954
rect 267326 88398 267562 88634
rect 267646 88398 267882 88634
rect 267326 52718 267562 52954
rect 267646 52718 267882 52954
rect 267326 52398 267562 52634
rect 267646 52398 267882 52634
rect 267326 16718 267562 16954
rect 267646 16718 267882 16954
rect 267326 16398 267562 16634
rect 267646 16398 267882 16634
rect 267326 -3462 267562 -3226
rect 267646 -3462 267882 -3226
rect 267326 -3782 267562 -3546
rect 267646 -3782 267882 -3546
rect 271826 708442 272062 708678
rect 272146 708442 272382 708678
rect 271826 708122 272062 708358
rect 272146 708122 272382 708358
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 276326 709402 276562 709638
rect 276646 709402 276882 709638
rect 276326 709082 276562 709318
rect 276646 709082 276882 709318
rect 276326 673718 276562 673954
rect 276646 673718 276882 673954
rect 276326 673398 276562 673634
rect 276646 673398 276882 673634
rect 280826 710362 281062 710598
rect 281146 710362 281382 710598
rect 280826 710042 281062 710278
rect 281146 710042 281382 710278
rect 280826 678218 281062 678454
rect 281146 678218 281382 678454
rect 280826 677898 281062 678134
rect 281146 677898 281382 678134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 285326 711322 285562 711558
rect 285646 711322 285882 711558
rect 285326 711002 285562 711238
rect 285646 711002 285882 711238
rect 285326 682718 285562 682954
rect 285646 682718 285882 682954
rect 285326 682398 285562 682634
rect 285646 682398 285882 682634
rect 280826 642125 281062 642361
rect 281146 642125 281382 642361
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 285326 646718 285562 646954
rect 285646 646718 285882 646954
rect 285326 646398 285562 646634
rect 285646 646398 285882 646634
rect 284250 615218 284486 615454
rect 284250 614898 284486 615134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 294326 705562 294562 705798
rect 294646 705562 294882 705798
rect 294326 705242 294562 705478
rect 294646 705242 294882 705478
rect 294326 691718 294562 691954
rect 294646 691718 294882 691954
rect 294326 691398 294562 691634
rect 294646 691398 294882 691634
rect 298826 706522 299062 706758
rect 299146 706522 299382 706758
rect 298826 706202 299062 706438
rect 299146 706202 299382 706438
rect 298826 696218 299062 696454
rect 299146 696218 299382 696454
rect 298826 695898 299062 696134
rect 299146 695898 299382 696134
rect 294326 655718 294562 655954
rect 294646 655718 294882 655954
rect 294326 655398 294562 655634
rect 294646 655398 294882 655634
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 294326 583718 294562 583954
rect 294646 583718 294882 583954
rect 294326 583398 294562 583634
rect 294646 583398 294882 583634
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -4422 272062 -4186
rect 272146 -4422 272382 -4186
rect 271826 -4742 272062 -4506
rect 272146 -4742 272382 -4506
rect 276326 493718 276562 493954
rect 276646 493718 276882 493954
rect 276326 493398 276562 493634
rect 276646 493398 276882 493634
rect 276326 457718 276562 457954
rect 276646 457718 276882 457954
rect 276326 457398 276562 457634
rect 276646 457398 276882 457634
rect 276326 421718 276562 421954
rect 276646 421718 276882 421954
rect 276326 421398 276562 421634
rect 276646 421398 276882 421634
rect 276326 385718 276562 385954
rect 276646 385718 276882 385954
rect 276326 385398 276562 385634
rect 276646 385398 276882 385634
rect 276326 349718 276562 349954
rect 276646 349718 276882 349954
rect 276326 349398 276562 349634
rect 276646 349398 276882 349634
rect 276326 313718 276562 313954
rect 276646 313718 276882 313954
rect 276326 313398 276562 313634
rect 276646 313398 276882 313634
rect 276326 277718 276562 277954
rect 276646 277718 276882 277954
rect 276326 277398 276562 277634
rect 276646 277398 276882 277634
rect 276326 241718 276562 241954
rect 276646 241718 276882 241954
rect 276326 241398 276562 241634
rect 276646 241398 276882 241634
rect 276326 205718 276562 205954
rect 276646 205718 276882 205954
rect 276326 205398 276562 205634
rect 276646 205398 276882 205634
rect 276326 169718 276562 169954
rect 276646 169718 276882 169954
rect 276326 169398 276562 169634
rect 276646 169398 276882 169634
rect 276326 133718 276562 133954
rect 276646 133718 276882 133954
rect 276326 133398 276562 133634
rect 276646 133398 276882 133634
rect 276326 97718 276562 97954
rect 276646 97718 276882 97954
rect 276326 97398 276562 97634
rect 276646 97398 276882 97634
rect 276326 61718 276562 61954
rect 276646 61718 276882 61954
rect 276326 61398 276562 61634
rect 276646 61398 276882 61634
rect 276326 25718 276562 25954
rect 276646 25718 276882 25954
rect 276326 25398 276562 25634
rect 276646 25398 276882 25634
rect 276326 -5382 276562 -5146
rect 276646 -5382 276882 -5146
rect 276326 -5702 276562 -5466
rect 276646 -5702 276882 -5466
rect 280826 462218 281062 462454
rect 281146 462218 281382 462454
rect 280826 461898 281062 462134
rect 281146 461898 281382 462134
rect 280826 426218 281062 426454
rect 281146 426218 281382 426454
rect 280826 425898 281062 426134
rect 281146 425898 281382 426134
rect 280826 390218 281062 390454
rect 281146 390218 281382 390454
rect 280826 389898 281062 390134
rect 281146 389898 281382 390134
rect 280826 354218 281062 354454
rect 281146 354218 281382 354454
rect 280826 353898 281062 354134
rect 281146 353898 281382 354134
rect 280826 318218 281062 318454
rect 281146 318218 281382 318454
rect 280826 317898 281062 318134
rect 281146 317898 281382 318134
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 294326 547718 294562 547954
rect 294646 547718 294882 547954
rect 294326 547398 294562 547634
rect 294646 547398 294882 547634
rect 298826 660218 299062 660454
rect 299146 660218 299382 660454
rect 298826 659898 299062 660134
rect 299146 659898 299382 660134
rect 303326 707482 303562 707718
rect 303646 707482 303882 707718
rect 303326 707162 303562 707398
rect 303646 707162 303882 707398
rect 303326 700718 303562 700954
rect 303646 700718 303882 700954
rect 303326 700398 303562 700634
rect 303646 700398 303882 700634
rect 303326 664718 303562 664954
rect 303646 664718 303882 664954
rect 303326 664398 303562 664634
rect 303646 664398 303882 664634
rect 307826 708442 308062 708678
rect 308146 708442 308382 708678
rect 307826 708122 308062 708358
rect 308146 708122 308382 708358
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 312326 709402 312562 709638
rect 312646 709402 312882 709638
rect 312326 709082 312562 709318
rect 312646 709082 312882 709318
rect 312326 673718 312562 673954
rect 312646 673718 312882 673954
rect 312326 673398 312562 673634
rect 312646 673398 312882 673634
rect 299610 619718 299846 619954
rect 299610 619398 299846 619634
rect 298826 588218 299062 588454
rect 299146 588218 299382 588454
rect 298826 587898 299062 588134
rect 299146 587898 299382 588134
rect 298826 552218 299062 552454
rect 299146 552218 299382 552454
rect 298826 551898 299062 552134
rect 299146 551898 299382 552134
rect 303326 592718 303562 592954
rect 303646 592718 303882 592954
rect 303326 592398 303562 592634
rect 303646 592398 303882 592634
rect 303326 556718 303562 556954
rect 303646 556718 303882 556954
rect 303326 556398 303562 556634
rect 303646 556398 303882 556634
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 316826 710362 317062 710598
rect 317146 710362 317382 710598
rect 316826 710042 317062 710278
rect 317146 710042 317382 710278
rect 316826 678218 317062 678454
rect 317146 678218 317382 678454
rect 316826 677898 317062 678134
rect 317146 677898 317382 678134
rect 321326 711322 321562 711558
rect 321646 711322 321882 711558
rect 321326 711002 321562 711238
rect 321646 711002 321882 711238
rect 321326 682718 321562 682954
rect 321646 682718 321882 682954
rect 321326 682398 321562 682634
rect 321646 682398 321882 682634
rect 316826 642125 317062 642361
rect 317146 642125 317382 642361
rect 314970 615218 315206 615454
rect 314970 614898 315206 615134
rect 321326 646718 321562 646954
rect 321646 646718 321882 646954
rect 321326 646398 321562 646634
rect 321646 646398 321882 646634
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 284250 507218 284486 507454
rect 284250 506898 284486 507134
rect 285326 466718 285562 466954
rect 285646 466718 285882 466954
rect 285326 466398 285562 466634
rect 285646 466398 285882 466634
rect 285326 430718 285562 430954
rect 285646 430718 285882 430954
rect 285326 430398 285562 430634
rect 285646 430398 285882 430634
rect 285326 394718 285562 394954
rect 285646 394718 285882 394954
rect 285326 394398 285562 394634
rect 285646 394398 285882 394634
rect 285326 358718 285562 358954
rect 285646 358718 285882 358954
rect 285326 358398 285562 358634
rect 285646 358398 285882 358634
rect 285326 322718 285562 322954
rect 285646 322718 285882 322954
rect 285326 322398 285562 322634
rect 285646 322398 285882 322634
rect 285326 286718 285562 286954
rect 285646 286718 285882 286954
rect 285326 286398 285562 286634
rect 285646 286398 285882 286634
rect 280826 246218 281062 246454
rect 281146 246218 281382 246454
rect 280826 245898 281062 246134
rect 281146 245898 281382 246134
rect 280826 210218 281062 210454
rect 281146 210218 281382 210454
rect 280826 209898 281062 210134
rect 281146 209898 281382 210134
rect 280826 174218 281062 174454
rect 281146 174218 281382 174454
rect 280826 173898 281062 174134
rect 281146 173898 281382 174134
rect 280826 138218 281062 138454
rect 281146 138218 281382 138454
rect 280826 137898 281062 138134
rect 281146 137898 281382 138134
rect 280826 102218 281062 102454
rect 281146 102218 281382 102454
rect 280826 101898 281062 102134
rect 281146 101898 281382 102134
rect 280826 66218 281062 66454
rect 281146 66218 281382 66454
rect 280826 65898 281062 66134
rect 281146 65898 281382 66134
rect 280826 30218 281062 30454
rect 281146 30218 281382 30454
rect 280826 29898 281062 30134
rect 281146 29898 281382 30134
rect 280826 -6342 281062 -6106
rect 281146 -6342 281382 -6106
rect 280826 -6662 281062 -6426
rect 281146 -6662 281382 -6426
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 285326 250718 285562 250954
rect 285646 250718 285882 250954
rect 285326 250398 285562 250634
rect 285646 250398 285882 250634
rect 285326 214718 285562 214954
rect 285646 214718 285882 214954
rect 285326 214398 285562 214634
rect 285646 214398 285882 214634
rect 285326 178718 285562 178954
rect 285646 178718 285882 178954
rect 285326 178398 285562 178634
rect 285646 178398 285882 178634
rect 285326 142718 285562 142954
rect 285646 142718 285882 142954
rect 285326 142398 285562 142634
rect 285646 142398 285882 142634
rect 285326 106718 285562 106954
rect 285646 106718 285882 106954
rect 285326 106398 285562 106634
rect 285646 106398 285882 106634
rect 285326 70718 285562 70954
rect 285646 70718 285882 70954
rect 285326 70398 285562 70634
rect 285646 70398 285882 70634
rect 285326 34718 285562 34954
rect 285646 34718 285882 34954
rect 285326 34398 285562 34634
rect 285646 34398 285882 34634
rect 285326 -7302 285562 -7066
rect 285646 -7302 285882 -7066
rect 285326 -7622 285562 -7386
rect 285646 -7622 285882 -7386
rect 294326 475718 294562 475954
rect 294646 475718 294882 475954
rect 294326 475398 294562 475634
rect 294646 475398 294882 475634
rect 294326 439718 294562 439954
rect 294646 439718 294882 439954
rect 294326 439398 294562 439634
rect 294646 439398 294882 439634
rect 294326 403718 294562 403954
rect 294646 403718 294882 403954
rect 294326 403398 294562 403634
rect 294646 403398 294882 403634
rect 294326 367718 294562 367954
rect 294646 367718 294882 367954
rect 294326 367398 294562 367634
rect 294646 367398 294882 367634
rect 294326 331718 294562 331954
rect 294646 331718 294882 331954
rect 294326 331398 294562 331634
rect 294646 331398 294882 331634
rect 294326 295718 294562 295954
rect 294646 295718 294882 295954
rect 294326 295398 294562 295634
rect 294646 295398 294882 295634
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 299610 511718 299846 511954
rect 299610 511398 299846 511634
rect 314970 507218 315206 507454
rect 314970 506898 315206 507134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 298826 480218 299062 480454
rect 299146 480218 299382 480454
rect 298826 479898 299062 480134
rect 299146 479898 299382 480134
rect 298826 444218 299062 444454
rect 299146 444218 299382 444454
rect 298826 443898 299062 444134
rect 299146 443898 299382 444134
rect 298826 408218 299062 408454
rect 299146 408218 299382 408454
rect 298826 407898 299062 408134
rect 299146 407898 299382 408134
rect 298826 372218 299062 372454
rect 299146 372218 299382 372454
rect 298826 371898 299062 372134
rect 299146 371898 299382 372134
rect 294326 259718 294562 259954
rect 294646 259718 294882 259954
rect 294326 259398 294562 259634
rect 294646 259398 294882 259634
rect 294326 223718 294562 223954
rect 294646 223718 294882 223954
rect 294326 223398 294562 223634
rect 294646 223398 294882 223634
rect 294326 187718 294562 187954
rect 294646 187718 294882 187954
rect 294326 187398 294562 187634
rect 294646 187398 294882 187634
rect 294326 151718 294562 151954
rect 294646 151718 294882 151954
rect 294326 151398 294562 151634
rect 294646 151398 294882 151634
rect 294326 115718 294562 115954
rect 294646 115718 294882 115954
rect 294326 115398 294562 115634
rect 294646 115398 294882 115634
rect 294326 79718 294562 79954
rect 294646 79718 294882 79954
rect 294326 79398 294562 79634
rect 294646 79398 294882 79634
rect 294326 43718 294562 43954
rect 294646 43718 294882 43954
rect 294326 43398 294562 43634
rect 294646 43398 294882 43634
rect 294326 7718 294562 7954
rect 294646 7718 294882 7954
rect 294326 7398 294562 7634
rect 294646 7398 294882 7634
rect 298826 336218 299062 336454
rect 299146 336218 299382 336454
rect 298826 335898 299062 336134
rect 299146 335898 299382 336134
rect 303326 484718 303562 484954
rect 303646 484718 303882 484954
rect 303326 484398 303562 484634
rect 303646 484398 303882 484634
rect 303326 448718 303562 448954
rect 303646 448718 303882 448954
rect 303326 448398 303562 448634
rect 303646 448398 303882 448634
rect 303326 412718 303562 412954
rect 303646 412718 303882 412954
rect 303326 412398 303562 412634
rect 303646 412398 303882 412634
rect 303326 376718 303562 376954
rect 303646 376718 303882 376954
rect 303326 376398 303562 376634
rect 303646 376398 303882 376634
rect 303326 340718 303562 340954
rect 303646 340718 303882 340954
rect 303326 340398 303562 340634
rect 303646 340398 303882 340634
rect 298826 264218 299062 264454
rect 299146 264218 299382 264454
rect 298826 263898 299062 264134
rect 299146 263898 299382 264134
rect 298826 228218 299062 228454
rect 299146 228218 299382 228454
rect 298826 227898 299062 228134
rect 299146 227898 299382 228134
rect 298826 48218 299062 48454
rect 299146 48218 299382 48454
rect 298826 47898 299062 48134
rect 299146 47898 299382 48134
rect 298826 12218 299062 12454
rect 299146 12218 299382 12454
rect 298826 11898 299062 12134
rect 299146 11898 299382 12134
rect 294326 -1542 294562 -1306
rect 294646 -1542 294882 -1306
rect 294326 -1862 294562 -1626
rect 294646 -1862 294882 -1626
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 312326 493718 312562 493954
rect 312646 493718 312882 493954
rect 312326 493398 312562 493634
rect 312646 493398 312882 493634
rect 312326 457718 312562 457954
rect 312646 457718 312882 457954
rect 312326 457398 312562 457634
rect 312646 457398 312882 457634
rect 312326 421718 312562 421954
rect 312646 421718 312882 421954
rect 312326 421398 312562 421634
rect 312646 421398 312882 421634
rect 312326 385718 312562 385954
rect 312646 385718 312882 385954
rect 312326 385398 312562 385634
rect 312646 385398 312882 385634
rect 312326 349718 312562 349954
rect 312646 349718 312882 349954
rect 312326 349398 312562 349634
rect 312646 349398 312882 349634
rect 316826 462218 317062 462454
rect 317146 462218 317382 462454
rect 316826 461898 317062 462134
rect 317146 461898 317382 462134
rect 316826 426218 317062 426454
rect 317146 426218 317382 426454
rect 316826 425898 317062 426134
rect 317146 425898 317382 426134
rect 316826 390218 317062 390454
rect 317146 390218 317382 390454
rect 316826 389898 317062 390134
rect 317146 389898 317382 390134
rect 316826 354218 317062 354454
rect 317146 354218 317382 354454
rect 316826 353898 317062 354134
rect 317146 353898 317382 354134
rect 321326 466718 321562 466954
rect 321646 466718 321882 466954
rect 321326 466398 321562 466634
rect 321646 466398 321882 466634
rect 321326 430718 321562 430954
rect 321646 430718 321882 430954
rect 321326 430398 321562 430634
rect 321646 430398 321882 430634
rect 321326 394718 321562 394954
rect 321646 394718 321882 394954
rect 321326 394398 321562 394634
rect 321646 394398 321882 394634
rect 321326 358718 321562 358954
rect 321646 358718 321882 358954
rect 321326 358398 321562 358634
rect 321646 358398 321882 358634
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 330326 705562 330562 705798
rect 330646 705562 330882 705798
rect 330326 705242 330562 705478
rect 330646 705242 330882 705478
rect 330326 691718 330562 691954
rect 330646 691718 330882 691954
rect 330326 691398 330562 691634
rect 330646 691398 330882 691634
rect 330326 655718 330562 655954
rect 330646 655718 330882 655954
rect 330326 655398 330562 655634
rect 330646 655398 330882 655634
rect 330326 619718 330562 619954
rect 330646 619718 330882 619954
rect 330326 619398 330562 619634
rect 330646 619398 330882 619634
rect 330326 583718 330562 583954
rect 330646 583718 330882 583954
rect 330326 583398 330562 583634
rect 330646 583398 330882 583634
rect 330326 547718 330562 547954
rect 330646 547718 330882 547954
rect 330326 547398 330562 547634
rect 330646 547398 330882 547634
rect 330326 511718 330562 511954
rect 330646 511718 330882 511954
rect 330326 511398 330562 511634
rect 330646 511398 330882 511634
rect 330326 475718 330562 475954
rect 330646 475718 330882 475954
rect 330326 475398 330562 475634
rect 330646 475398 330882 475634
rect 330326 439718 330562 439954
rect 330646 439718 330882 439954
rect 330326 439398 330562 439634
rect 330646 439398 330882 439634
rect 330326 403718 330562 403954
rect 330646 403718 330882 403954
rect 330326 403398 330562 403634
rect 330646 403398 330882 403634
rect 330326 367718 330562 367954
rect 330646 367718 330882 367954
rect 330326 367398 330562 367634
rect 330646 367398 330882 367634
rect 334826 706522 335062 706758
rect 335146 706522 335382 706758
rect 334826 706202 335062 706438
rect 335146 706202 335382 706438
rect 334826 696218 335062 696454
rect 335146 696218 335382 696454
rect 334826 695898 335062 696134
rect 335146 695898 335382 696134
rect 334826 660218 335062 660454
rect 335146 660218 335382 660454
rect 334826 659898 335062 660134
rect 335146 659898 335382 660134
rect 334826 624218 335062 624454
rect 335146 624218 335382 624454
rect 334826 623898 335062 624134
rect 335146 623898 335382 624134
rect 334826 588218 335062 588454
rect 335146 588218 335382 588454
rect 334826 587898 335062 588134
rect 335146 587898 335382 588134
rect 334826 552218 335062 552454
rect 335146 552218 335382 552454
rect 334826 551898 335062 552134
rect 335146 551898 335382 552134
rect 334826 516218 335062 516454
rect 335146 516218 335382 516454
rect 334826 515898 335062 516134
rect 335146 515898 335382 516134
rect 334826 480218 335062 480454
rect 335146 480218 335382 480454
rect 334826 479898 335062 480134
rect 335146 479898 335382 480134
rect 334826 444218 335062 444454
rect 335146 444218 335382 444454
rect 334826 443898 335062 444134
rect 335146 443898 335382 444134
rect 334826 408218 335062 408454
rect 335146 408218 335382 408454
rect 334826 407898 335062 408134
rect 335146 407898 335382 408134
rect 334826 372218 335062 372454
rect 335146 372218 335382 372454
rect 334826 371898 335062 372134
rect 335146 371898 335382 372134
rect 334826 336218 335062 336454
rect 335146 336218 335382 336454
rect 334826 335898 335062 336134
rect 335146 335898 335382 336134
rect 339326 707482 339562 707718
rect 339646 707482 339882 707718
rect 339326 707162 339562 707398
rect 339646 707162 339882 707398
rect 339326 700718 339562 700954
rect 339646 700718 339882 700954
rect 339326 700398 339562 700634
rect 339646 700398 339882 700634
rect 339326 664718 339562 664954
rect 339646 664718 339882 664954
rect 339326 664398 339562 664634
rect 339646 664398 339882 664634
rect 339326 628718 339562 628954
rect 339646 628718 339882 628954
rect 339326 628398 339562 628634
rect 339646 628398 339882 628634
rect 339326 592718 339562 592954
rect 339646 592718 339882 592954
rect 339326 592398 339562 592634
rect 339646 592398 339882 592634
rect 339326 556718 339562 556954
rect 339646 556718 339882 556954
rect 339326 556398 339562 556634
rect 339646 556398 339882 556634
rect 339326 520718 339562 520954
rect 339646 520718 339882 520954
rect 339326 520398 339562 520634
rect 339646 520398 339882 520634
rect 339326 484718 339562 484954
rect 339646 484718 339882 484954
rect 339326 484398 339562 484634
rect 339646 484398 339882 484634
rect 339326 448718 339562 448954
rect 339646 448718 339882 448954
rect 339326 448398 339562 448634
rect 339646 448398 339882 448634
rect 339326 412718 339562 412954
rect 339646 412718 339882 412954
rect 339326 412398 339562 412634
rect 339646 412398 339882 412634
rect 339326 376718 339562 376954
rect 339646 376718 339882 376954
rect 339326 376398 339562 376634
rect 339646 376398 339882 376634
rect 339326 340718 339562 340954
rect 339646 340718 339882 340954
rect 339326 340398 339562 340634
rect 339646 340398 339882 340634
rect 343826 708442 344062 708678
rect 344146 708442 344382 708678
rect 343826 708122 344062 708358
rect 344146 708122 344382 708358
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 348326 709402 348562 709638
rect 348646 709402 348882 709638
rect 348326 709082 348562 709318
rect 348646 709082 348882 709318
rect 348326 673718 348562 673954
rect 348646 673718 348882 673954
rect 348326 673398 348562 673634
rect 348646 673398 348882 673634
rect 352826 710362 353062 710598
rect 353146 710362 353382 710598
rect 352826 710042 353062 710278
rect 353146 710042 353382 710278
rect 352826 678218 353062 678454
rect 353146 678218 353382 678454
rect 352826 677898 353062 678134
rect 353146 677898 353382 678134
rect 352826 642218 353062 642454
rect 353146 642218 353382 642454
rect 352826 641898 353062 642134
rect 353146 641898 353382 642134
rect 357326 711322 357562 711558
rect 357646 711322 357882 711558
rect 357326 711002 357562 711238
rect 357646 711002 357882 711238
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 357326 682718 357562 682954
rect 357646 682718 357882 682954
rect 357326 682398 357562 682634
rect 357646 682398 357882 682634
rect 357326 646718 357562 646954
rect 357646 646718 357882 646954
rect 357326 646398 357562 646634
rect 357646 646398 357882 646634
rect 348326 637718 348562 637954
rect 348646 637718 348882 637954
rect 348326 637398 348562 637634
rect 348646 637398 348882 637634
rect 348326 601718 348562 601954
rect 348646 601718 348882 601954
rect 348326 601398 348562 601634
rect 348646 601398 348882 601634
rect 348326 565718 348562 565954
rect 348646 565718 348882 565954
rect 348326 565398 348562 565634
rect 348646 565398 348882 565634
rect 348326 529718 348562 529954
rect 348646 529718 348882 529954
rect 348326 529398 348562 529634
rect 348646 529398 348882 529634
rect 348326 493718 348562 493954
rect 348646 493718 348882 493954
rect 348326 493398 348562 493634
rect 348646 493398 348882 493634
rect 348326 457718 348562 457954
rect 348646 457718 348882 457954
rect 348326 457398 348562 457634
rect 348646 457398 348882 457634
rect 348326 421718 348562 421954
rect 348646 421718 348882 421954
rect 348326 421398 348562 421634
rect 348646 421398 348882 421634
rect 348326 385718 348562 385954
rect 348646 385718 348882 385954
rect 348326 385398 348562 385634
rect 348646 385398 348882 385634
rect 348326 349718 348562 349954
rect 348646 349718 348882 349954
rect 348326 349398 348562 349634
rect 348646 349398 348882 349634
rect 304250 327003 304486 327239
rect 334970 327003 335206 327239
rect 319610 295718 319846 295954
rect 319610 295398 319846 295634
rect 304250 291218 304486 291454
rect 304250 290898 304486 291134
rect 334970 291218 335206 291454
rect 334970 290898 335206 291134
rect 303326 268718 303562 268954
rect 303646 268718 303882 268954
rect 303326 268398 303562 268634
rect 303646 268398 303882 268634
rect 303326 232718 303562 232954
rect 303646 232718 303882 232954
rect 303326 232398 303562 232634
rect 303646 232398 303882 232634
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 312326 277718 312562 277954
rect 312646 277718 312882 277954
rect 312326 277398 312562 277634
rect 312646 277398 312882 277634
rect 312326 241718 312562 241954
rect 312646 241718 312882 241954
rect 312326 241398 312562 241634
rect 312646 241398 312882 241634
rect 330326 259718 330562 259954
rect 330646 259718 330882 259954
rect 330326 259398 330562 259634
rect 330646 259398 330882 259634
rect 330326 223718 330562 223954
rect 330646 223718 330882 223954
rect 330326 223398 330562 223634
rect 330646 223398 330882 223634
rect 334826 264218 335062 264454
rect 335146 264218 335382 264454
rect 334826 263898 335062 264134
rect 335146 263898 335382 264134
rect 334826 228218 335062 228454
rect 335146 228218 335382 228454
rect 334826 227898 335062 228134
rect 335146 227898 335382 228134
rect 339326 268718 339562 268954
rect 339646 268718 339882 268954
rect 339326 268398 339562 268634
rect 339646 268398 339882 268634
rect 339326 232718 339562 232954
rect 339646 232718 339882 232954
rect 339326 232398 339562 232634
rect 339646 232398 339882 232634
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 348326 277718 348562 277954
rect 348646 277718 348882 277954
rect 348326 277398 348562 277634
rect 348646 277398 348882 277634
rect 348326 241718 348562 241954
rect 348646 241718 348882 241954
rect 348326 241398 348562 241634
rect 348646 241398 348882 241634
rect 348326 205718 348562 205954
rect 348646 205718 348882 205954
rect 348326 205398 348562 205634
rect 348646 205398 348882 205634
rect 319610 187718 319846 187954
rect 319610 187398 319846 187634
rect 304250 183218 304486 183454
rect 304250 182898 304486 183134
rect 334970 183218 335206 183454
rect 334970 182898 335206 183134
rect 348326 169718 348562 169954
rect 348646 169718 348882 169954
rect 348326 169398 348562 169634
rect 348646 169398 348882 169634
rect 319610 151718 319846 151954
rect 319610 151398 319846 151634
rect 304250 147218 304486 147454
rect 304250 146898 304486 147134
rect 334970 147218 335206 147454
rect 334970 146898 335206 147134
rect 348326 133718 348562 133954
rect 348646 133718 348882 133954
rect 348326 133398 348562 133634
rect 348646 133398 348882 133634
rect 319610 115718 319846 115954
rect 319610 115398 319846 115634
rect 304250 111218 304486 111454
rect 304250 110898 304486 111134
rect 334970 111218 335206 111454
rect 334970 110898 335206 111134
rect 319610 79718 319846 79954
rect 319610 79398 319846 79634
rect 304250 75218 304486 75454
rect 304250 74898 304486 75134
rect 334970 75218 335206 75454
rect 334970 74898 335206 75134
rect 303326 52718 303562 52954
rect 303646 52718 303882 52954
rect 303326 52398 303562 52634
rect 303646 52398 303882 52634
rect 303326 16718 303562 16954
rect 303646 16718 303882 16954
rect 303326 16398 303562 16634
rect 303646 16398 303882 16634
rect 298826 -2502 299062 -2266
rect 299146 -2502 299382 -2266
rect 298826 -2822 299062 -2586
rect 299146 -2822 299382 -2586
rect 303326 -3462 303562 -3226
rect 303646 -3462 303882 -3226
rect 303326 -3782 303562 -3546
rect 303646 -3782 303882 -3546
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -4422 308062 -4186
rect 308146 -4422 308382 -4186
rect 307826 -4742 308062 -4506
rect 308146 -4742 308382 -4506
rect 312326 25718 312562 25954
rect 312646 25718 312882 25954
rect 312326 25398 312562 25634
rect 312646 25398 312882 25634
rect 312326 -5382 312562 -5146
rect 312646 -5382 312882 -5146
rect 312326 -5702 312562 -5466
rect 312646 -5702 312882 -5466
rect 316826 30218 317062 30454
rect 317146 30218 317382 30454
rect 316826 29898 317062 30134
rect 317146 29898 317382 30134
rect 316826 -6342 317062 -6106
rect 317146 -6342 317382 -6106
rect 316826 -6662 317062 -6426
rect 317146 -6662 317382 -6426
rect 321326 34718 321562 34954
rect 321646 34718 321882 34954
rect 321326 34398 321562 34634
rect 321646 34398 321882 34634
rect 321326 -7302 321562 -7066
rect 321646 -7302 321882 -7066
rect 321326 -7622 321562 -7386
rect 321646 -7622 321882 -7386
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 330326 43718 330562 43954
rect 330646 43718 330882 43954
rect 330326 43398 330562 43634
rect 330646 43398 330882 43634
rect 330326 7718 330562 7954
rect 330646 7718 330882 7954
rect 330326 7398 330562 7634
rect 330646 7398 330882 7634
rect 330326 -1542 330562 -1306
rect 330646 -1542 330882 -1306
rect 330326 -1862 330562 -1626
rect 330646 -1862 330882 -1626
rect 334826 48218 335062 48454
rect 335146 48218 335382 48454
rect 334826 47898 335062 48134
rect 335146 47898 335382 48134
rect 334826 12218 335062 12454
rect 335146 12218 335382 12454
rect 334826 11898 335062 12134
rect 335146 11898 335382 12134
rect 334826 -2502 335062 -2266
rect 335146 -2502 335382 -2266
rect 334826 -2822 335062 -2586
rect 335146 -2822 335382 -2586
rect 339326 52718 339562 52954
rect 339646 52718 339882 52954
rect 339326 52398 339562 52634
rect 339646 52398 339882 52634
rect 339326 16718 339562 16954
rect 339646 16718 339882 16954
rect 339326 16398 339562 16634
rect 339646 16398 339882 16634
rect 348326 97718 348562 97954
rect 348646 97718 348882 97954
rect 348326 97398 348562 97634
rect 348646 97398 348882 97634
rect 348326 61718 348562 61954
rect 348646 61718 348882 61954
rect 348326 61398 348562 61634
rect 348646 61398 348882 61634
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 339326 -3462 339562 -3226
rect 339646 -3462 339882 -3226
rect 339326 -3782 339562 -3546
rect 339646 -3782 339882 -3546
rect 343826 -4422 344062 -4186
rect 344146 -4422 344382 -4186
rect 343826 -4742 344062 -4506
rect 344146 -4742 344382 -4506
rect 348326 25718 348562 25954
rect 348646 25718 348882 25954
rect 348326 25398 348562 25634
rect 348646 25398 348882 25634
rect 352826 606218 353062 606454
rect 353146 606218 353382 606454
rect 352826 605898 353062 606134
rect 353146 605898 353382 606134
rect 352826 570218 353062 570454
rect 353146 570218 353382 570454
rect 352826 569898 353062 570134
rect 353146 569898 353382 570134
rect 352826 534218 353062 534454
rect 353146 534218 353382 534454
rect 352826 533898 353062 534134
rect 353146 533898 353382 534134
rect 352826 498218 353062 498454
rect 353146 498218 353382 498454
rect 352826 497898 353062 498134
rect 353146 497898 353382 498134
rect 352826 462218 353062 462454
rect 353146 462218 353382 462454
rect 352826 461898 353062 462134
rect 353146 461898 353382 462134
rect 352826 426218 353062 426454
rect 353146 426218 353382 426454
rect 352826 425898 353062 426134
rect 353146 425898 353382 426134
rect 352826 390218 353062 390454
rect 353146 390218 353382 390454
rect 352826 389898 353062 390134
rect 353146 389898 353382 390134
rect 352826 354218 353062 354454
rect 353146 354218 353382 354454
rect 352826 353898 353062 354134
rect 353146 353898 353382 354134
rect 352826 246218 353062 246454
rect 353146 246218 353382 246454
rect 352826 245898 353062 246134
rect 353146 245898 353382 246134
rect 352826 210218 353062 210454
rect 353146 210218 353382 210454
rect 352826 209898 353062 210134
rect 353146 209898 353382 210134
rect 352826 174218 353062 174454
rect 353146 174218 353382 174454
rect 352826 173898 353062 174134
rect 353146 173898 353382 174134
rect 352826 138218 353062 138454
rect 353146 138218 353382 138454
rect 352826 137898 353062 138134
rect 353146 137898 353382 138134
rect 352826 102218 353062 102454
rect 353146 102218 353382 102454
rect 352826 101898 353062 102134
rect 353146 101898 353382 102134
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 366326 705562 366562 705798
rect 366646 705562 366882 705798
rect 366326 705242 366562 705478
rect 366646 705242 366882 705478
rect 366326 691718 366562 691954
rect 366646 691718 366882 691954
rect 366326 691398 366562 691634
rect 366646 691398 366882 691634
rect 366326 655718 366562 655954
rect 366646 655718 366882 655954
rect 366326 655398 366562 655634
rect 366646 655398 366882 655634
rect 370826 706522 371062 706758
rect 371146 706522 371382 706758
rect 370826 706202 371062 706438
rect 371146 706202 371382 706438
rect 370826 696218 371062 696454
rect 371146 696218 371382 696454
rect 370826 695898 371062 696134
rect 371146 695898 371382 696134
rect 370826 660218 371062 660454
rect 371146 660218 371382 660454
rect 370826 659898 371062 660134
rect 371146 659898 371382 660134
rect 375326 707482 375562 707718
rect 375646 707482 375882 707718
rect 375326 707162 375562 707398
rect 375646 707162 375882 707398
rect 375326 700718 375562 700954
rect 375646 700718 375882 700954
rect 375326 700398 375562 700634
rect 375646 700398 375882 700634
rect 375326 664718 375562 664954
rect 375646 664718 375882 664954
rect 375326 664398 375562 664634
rect 375646 664398 375882 664634
rect 379826 708442 380062 708678
rect 380146 708442 380382 708678
rect 379826 708122 380062 708358
rect 380146 708122 380382 708358
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 384326 709402 384562 709638
rect 384646 709402 384882 709638
rect 384326 709082 384562 709318
rect 384646 709082 384882 709318
rect 384326 673718 384562 673954
rect 384646 673718 384882 673954
rect 384326 673398 384562 673634
rect 384646 673398 384882 673634
rect 388826 710362 389062 710598
rect 389146 710362 389382 710598
rect 388826 710042 389062 710278
rect 389146 710042 389382 710278
rect 388826 678218 389062 678454
rect 389146 678218 389382 678454
rect 388826 677898 389062 678134
rect 389146 677898 389382 678134
rect 388826 642125 389062 642361
rect 389146 642125 389382 642361
rect 393326 711322 393562 711558
rect 393646 711322 393882 711558
rect 393326 711002 393562 711238
rect 393646 711002 393882 711238
rect 393326 682718 393562 682954
rect 393646 682718 393882 682954
rect 393326 682398 393562 682634
rect 393646 682398 393882 682634
rect 393326 646718 393562 646954
rect 393646 646718 393882 646954
rect 393326 646398 393562 646634
rect 393646 646398 393882 646634
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 402326 705562 402562 705798
rect 402646 705562 402882 705798
rect 402326 705242 402562 705478
rect 402646 705242 402882 705478
rect 402326 691718 402562 691954
rect 402646 691718 402882 691954
rect 402326 691398 402562 691634
rect 402646 691398 402882 691634
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 379610 619718 379846 619954
rect 379610 619398 379846 619634
rect 364250 615218 364486 615454
rect 364250 614898 364486 615134
rect 394970 615218 395206 615454
rect 394970 614898 395206 615134
rect 364250 543218 364486 543454
rect 364250 542898 364486 543134
rect 364250 507218 364486 507454
rect 364250 506898 364486 507134
rect 370826 588218 371062 588454
rect 371146 588218 371382 588454
rect 370826 587898 371062 588134
rect 371146 587898 371382 588134
rect 375326 592718 375562 592954
rect 375646 592718 375882 592954
rect 375326 592398 375562 592634
rect 375646 592398 375882 592634
rect 370826 552125 371062 552361
rect 371146 552125 371382 552361
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 375326 556718 375562 556954
rect 375646 556718 375882 556954
rect 375326 556398 375562 556634
rect 375646 556398 375882 556634
rect 357326 466718 357562 466954
rect 357646 466718 357882 466954
rect 357326 466398 357562 466634
rect 357646 466398 357882 466634
rect 357326 430718 357562 430954
rect 357646 430718 357882 430954
rect 357326 430398 357562 430634
rect 357646 430398 357882 430634
rect 357326 394718 357562 394954
rect 357646 394718 357882 394954
rect 357326 394398 357562 394634
rect 357646 394398 357882 394634
rect 357326 358718 357562 358954
rect 357646 358718 357882 358954
rect 357326 358398 357562 358634
rect 357646 358398 357882 358634
rect 357326 322718 357562 322954
rect 357646 322718 357882 322954
rect 357326 322398 357562 322634
rect 357646 322398 357882 322634
rect 357326 286718 357562 286954
rect 357646 286718 357882 286954
rect 357326 286398 357562 286634
rect 357646 286398 357882 286634
rect 357326 250718 357562 250954
rect 357646 250718 357882 250954
rect 357326 250398 357562 250634
rect 357646 250398 357882 250634
rect 357326 214718 357562 214954
rect 357646 214718 357882 214954
rect 357326 214398 357562 214634
rect 357646 214398 357882 214634
rect 357326 178718 357562 178954
rect 357646 178718 357882 178954
rect 357326 178398 357562 178634
rect 357646 178398 357882 178634
rect 357326 142718 357562 142954
rect 357646 142718 357882 142954
rect 357326 142398 357562 142634
rect 357646 142398 357882 142634
rect 357326 106718 357562 106954
rect 357646 106718 357882 106954
rect 357326 106398 357562 106634
rect 357646 106398 357882 106634
rect 352826 66218 353062 66454
rect 353146 66218 353382 66454
rect 352826 65898 353062 66134
rect 353146 65898 353382 66134
rect 352826 30218 353062 30454
rect 353146 30218 353382 30454
rect 352826 29898 353062 30134
rect 353146 29898 353382 30134
rect 348326 -5382 348562 -5146
rect 348646 -5382 348882 -5146
rect 348326 -5702 348562 -5466
rect 348646 -5702 348882 -5466
rect 352826 -6342 353062 -6106
rect 353146 -6342 353382 -6106
rect 352826 -6662 353062 -6426
rect 353146 -6662 353382 -6426
rect 357326 70718 357562 70954
rect 357646 70718 357882 70954
rect 357326 70398 357562 70634
rect 357646 70398 357882 70634
rect 357326 34718 357562 34954
rect 357646 34718 357882 34954
rect 357326 34398 357562 34634
rect 357646 34398 357882 34634
rect 357326 -7302 357562 -7066
rect 357646 -7302 357882 -7066
rect 357326 -7622 357562 -7386
rect 357646 -7622 357882 -7386
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 366326 475718 366562 475954
rect 366646 475718 366882 475954
rect 366326 475398 366562 475634
rect 366646 475398 366882 475634
rect 366326 439718 366562 439954
rect 366646 439718 366882 439954
rect 366326 439398 366562 439634
rect 366646 439398 366882 439634
rect 366326 403718 366562 403954
rect 366646 403718 366882 403954
rect 366326 403398 366562 403634
rect 366646 403398 366882 403634
rect 366326 367718 366562 367954
rect 366646 367718 366882 367954
rect 366326 367398 366562 367634
rect 366646 367398 366882 367634
rect 366326 331718 366562 331954
rect 366646 331718 366882 331954
rect 366326 331398 366562 331634
rect 366646 331398 366882 331634
rect 366326 295718 366562 295954
rect 366646 295718 366882 295954
rect 366326 295398 366562 295634
rect 366646 295398 366882 295634
rect 366326 259718 366562 259954
rect 366646 259718 366882 259954
rect 366326 259398 366562 259634
rect 366646 259398 366882 259634
rect 366326 223718 366562 223954
rect 366646 223718 366882 223954
rect 366326 223398 366562 223634
rect 366646 223398 366882 223634
rect 366326 187718 366562 187954
rect 366646 187718 366882 187954
rect 366326 187398 366562 187634
rect 366646 187398 366882 187634
rect 366326 151718 366562 151954
rect 366646 151718 366882 151954
rect 366326 151398 366562 151634
rect 366646 151398 366882 151634
rect 366326 115718 366562 115954
rect 366646 115718 366882 115954
rect 366326 115398 366562 115634
rect 366646 115398 366882 115634
rect 366326 79718 366562 79954
rect 366646 79718 366882 79954
rect 366326 79398 366562 79634
rect 366646 79398 366882 79634
rect 366326 43718 366562 43954
rect 366646 43718 366882 43954
rect 366326 43398 366562 43634
rect 366646 43398 366882 43634
rect 366326 7718 366562 7954
rect 366646 7718 366882 7954
rect 366326 7398 366562 7634
rect 366646 7398 366882 7634
rect 366326 -1542 366562 -1306
rect 366646 -1542 366882 -1306
rect 366326 -1862 366562 -1626
rect 366646 -1862 366882 -1626
rect 370826 480218 371062 480454
rect 371146 480218 371382 480454
rect 370826 479898 371062 480134
rect 371146 479898 371382 480134
rect 370826 444218 371062 444454
rect 371146 444218 371382 444454
rect 370826 443898 371062 444134
rect 371146 443898 371382 444134
rect 370826 408218 371062 408454
rect 371146 408218 371382 408454
rect 370826 407898 371062 408134
rect 371146 407898 371382 408134
rect 370826 372218 371062 372454
rect 371146 372218 371382 372454
rect 370826 371898 371062 372134
rect 371146 371898 371382 372134
rect 370826 336218 371062 336454
rect 371146 336218 371382 336454
rect 370826 335898 371062 336134
rect 371146 335898 371382 336134
rect 370826 300218 371062 300454
rect 371146 300218 371382 300454
rect 370826 299898 371062 300134
rect 371146 299898 371382 300134
rect 370826 264218 371062 264454
rect 371146 264218 371382 264454
rect 370826 263898 371062 264134
rect 371146 263898 371382 264134
rect 370826 228218 371062 228454
rect 371146 228218 371382 228454
rect 370826 227898 371062 228134
rect 371146 227898 371382 228134
rect 370826 192218 371062 192454
rect 371146 192218 371382 192454
rect 370826 191898 371062 192134
rect 371146 191898 371382 192134
rect 370826 156218 371062 156454
rect 371146 156218 371382 156454
rect 370826 155898 371062 156134
rect 371146 155898 371382 156134
rect 370826 120218 371062 120454
rect 371146 120218 371382 120454
rect 370826 119898 371062 120134
rect 371146 119898 371382 120134
rect 370826 84218 371062 84454
rect 371146 84218 371382 84454
rect 370826 83898 371062 84134
rect 371146 83898 371382 84134
rect 370826 48218 371062 48454
rect 371146 48218 371382 48454
rect 370826 47898 371062 48134
rect 371146 47898 371382 48134
rect 370826 12218 371062 12454
rect 371146 12218 371382 12454
rect 370826 11898 371062 12134
rect 371146 11898 371382 12134
rect 370826 -2502 371062 -2266
rect 371146 -2502 371382 -2266
rect 370826 -2822 371062 -2586
rect 371146 -2822 371382 -2586
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379610 511718 379846 511954
rect 379610 511398 379846 511634
rect 375326 484718 375562 484954
rect 375646 484718 375882 484954
rect 375326 484398 375562 484634
rect 375646 484398 375882 484634
rect 375326 448718 375562 448954
rect 375646 448718 375882 448954
rect 375326 448398 375562 448634
rect 375646 448398 375882 448634
rect 375326 412718 375562 412954
rect 375646 412718 375882 412954
rect 375326 412398 375562 412634
rect 375646 412398 375882 412634
rect 375326 376718 375562 376954
rect 375646 376718 375882 376954
rect 375326 376398 375562 376634
rect 375646 376398 375882 376634
rect 375326 340718 375562 340954
rect 375646 340718 375882 340954
rect 375326 340398 375562 340634
rect 375646 340398 375882 340634
rect 375326 304718 375562 304954
rect 375646 304718 375882 304954
rect 375326 304398 375562 304634
rect 375646 304398 375882 304634
rect 375326 268718 375562 268954
rect 375646 268718 375882 268954
rect 375326 268398 375562 268634
rect 375646 268398 375882 268634
rect 375326 232718 375562 232954
rect 375646 232718 375882 232954
rect 375326 232398 375562 232634
rect 375646 232398 375882 232634
rect 375326 196718 375562 196954
rect 375646 196718 375882 196954
rect 375326 196398 375562 196634
rect 375646 196398 375882 196634
rect 375326 160718 375562 160954
rect 375646 160718 375882 160954
rect 375326 160398 375562 160634
rect 375646 160398 375882 160634
rect 375326 124718 375562 124954
rect 375646 124718 375882 124954
rect 375326 124398 375562 124634
rect 375646 124398 375882 124634
rect 375326 88718 375562 88954
rect 375646 88718 375882 88954
rect 375326 88398 375562 88634
rect 375646 88398 375882 88634
rect 375326 52718 375562 52954
rect 375646 52718 375882 52954
rect 375326 52398 375562 52634
rect 375646 52398 375882 52634
rect 375326 16718 375562 16954
rect 375646 16718 375882 16954
rect 375326 16398 375562 16634
rect 375646 16398 375882 16634
rect 375326 -3462 375562 -3226
rect 375646 -3462 375882 -3226
rect 375326 -3782 375562 -3546
rect 375646 -3782 375882 -3546
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -4422 380062 -4186
rect 380146 -4422 380382 -4186
rect 379826 -4742 380062 -4506
rect 380146 -4742 380382 -4506
rect 384326 493718 384562 493954
rect 384646 493718 384882 493954
rect 384326 493398 384562 493634
rect 384646 493398 384882 493634
rect 384326 457718 384562 457954
rect 384646 457718 384882 457954
rect 384326 457398 384562 457634
rect 384646 457398 384882 457634
rect 384326 421718 384562 421954
rect 384646 421718 384882 421954
rect 384326 421398 384562 421634
rect 384646 421398 384882 421634
rect 384326 385718 384562 385954
rect 384646 385718 384882 385954
rect 384326 385398 384562 385634
rect 384646 385398 384882 385634
rect 384326 349718 384562 349954
rect 384646 349718 384882 349954
rect 384326 349398 384562 349634
rect 384646 349398 384882 349634
rect 384326 313718 384562 313954
rect 384646 313718 384882 313954
rect 384326 313398 384562 313634
rect 384646 313398 384882 313634
rect 384326 277718 384562 277954
rect 384646 277718 384882 277954
rect 384326 277398 384562 277634
rect 384646 277398 384882 277634
rect 384326 241718 384562 241954
rect 384646 241718 384882 241954
rect 384326 241398 384562 241634
rect 384646 241398 384882 241634
rect 384326 205718 384562 205954
rect 384646 205718 384882 205954
rect 384326 205398 384562 205634
rect 384646 205398 384882 205634
rect 384326 169718 384562 169954
rect 384646 169718 384882 169954
rect 384326 169398 384562 169634
rect 384646 169398 384882 169634
rect 384326 133718 384562 133954
rect 384646 133718 384882 133954
rect 384326 133398 384562 133634
rect 384646 133398 384882 133634
rect 384326 97718 384562 97954
rect 384646 97718 384882 97954
rect 384326 97398 384562 97634
rect 384646 97398 384882 97634
rect 384326 61718 384562 61954
rect 384646 61718 384882 61954
rect 384326 61398 384562 61634
rect 384646 61398 384882 61634
rect 384326 25718 384562 25954
rect 384646 25718 384882 25954
rect 384326 25398 384562 25634
rect 384646 25398 384882 25634
rect 384326 -5382 384562 -5146
rect 384646 -5382 384882 -5146
rect 384326 -5702 384562 -5466
rect 384646 -5702 384882 -5466
rect 388826 462218 389062 462454
rect 389146 462218 389382 462454
rect 388826 461898 389062 462134
rect 389146 461898 389382 462134
rect 388826 426218 389062 426454
rect 389146 426218 389382 426454
rect 388826 425898 389062 426134
rect 389146 425898 389382 426134
rect 388826 390218 389062 390454
rect 389146 390218 389382 390454
rect 388826 389898 389062 390134
rect 389146 389898 389382 390134
rect 388826 354218 389062 354454
rect 389146 354218 389382 354454
rect 388826 353898 389062 354134
rect 389146 353898 389382 354134
rect 388826 318218 389062 318454
rect 389146 318218 389382 318454
rect 388826 317898 389062 318134
rect 389146 317898 389382 318134
rect 388826 282218 389062 282454
rect 389146 282218 389382 282454
rect 388826 281898 389062 282134
rect 389146 281898 389382 282134
rect 388826 246218 389062 246454
rect 389146 246218 389382 246454
rect 388826 245898 389062 246134
rect 389146 245898 389382 246134
rect 388826 210218 389062 210454
rect 389146 210218 389382 210454
rect 388826 209898 389062 210134
rect 389146 209898 389382 210134
rect 388826 174218 389062 174454
rect 389146 174218 389382 174454
rect 388826 173898 389062 174134
rect 389146 173898 389382 174134
rect 388826 138218 389062 138454
rect 389146 138218 389382 138454
rect 388826 137898 389062 138134
rect 389146 137898 389382 138134
rect 388826 102218 389062 102454
rect 389146 102218 389382 102454
rect 388826 101898 389062 102134
rect 389146 101898 389382 102134
rect 388826 66218 389062 66454
rect 389146 66218 389382 66454
rect 388826 65898 389062 66134
rect 389146 65898 389382 66134
rect 388826 30218 389062 30454
rect 389146 30218 389382 30454
rect 388826 29898 389062 30134
rect 389146 29898 389382 30134
rect 388826 -6342 389062 -6106
rect 389146 -6342 389382 -6106
rect 388826 -6662 389062 -6426
rect 389146 -6662 389382 -6426
rect 394970 543218 395206 543454
rect 394970 542898 395206 543134
rect 394970 507218 395206 507454
rect 394970 506898 395206 507134
rect 406826 706522 407062 706758
rect 407146 706522 407382 706758
rect 406826 706202 407062 706438
rect 407146 706202 407382 706438
rect 406826 696218 407062 696454
rect 407146 696218 407382 696454
rect 406826 695898 407062 696134
rect 407146 695898 407382 696134
rect 402326 655718 402562 655954
rect 402646 655718 402882 655954
rect 402326 655398 402562 655634
rect 402646 655398 402882 655634
rect 393326 466718 393562 466954
rect 393646 466718 393882 466954
rect 393326 466398 393562 466634
rect 393646 466398 393882 466634
rect 393326 430718 393562 430954
rect 393646 430718 393882 430954
rect 393326 430398 393562 430634
rect 393646 430398 393882 430634
rect 393326 394718 393562 394954
rect 393646 394718 393882 394954
rect 393326 394398 393562 394634
rect 393646 394398 393882 394634
rect 393326 358718 393562 358954
rect 393646 358718 393882 358954
rect 393326 358398 393562 358634
rect 393646 358398 393882 358634
rect 393326 322718 393562 322954
rect 393646 322718 393882 322954
rect 393326 322398 393562 322634
rect 393646 322398 393882 322634
rect 393326 286718 393562 286954
rect 393646 286718 393882 286954
rect 393326 286398 393562 286634
rect 393646 286398 393882 286634
rect 393326 250718 393562 250954
rect 393646 250718 393882 250954
rect 393326 250398 393562 250634
rect 393646 250398 393882 250634
rect 393326 214718 393562 214954
rect 393646 214718 393882 214954
rect 393326 214398 393562 214634
rect 393646 214398 393882 214634
rect 393326 178718 393562 178954
rect 393646 178718 393882 178954
rect 393326 178398 393562 178634
rect 393646 178398 393882 178634
rect 393326 142718 393562 142954
rect 393646 142718 393882 142954
rect 393326 142398 393562 142634
rect 393646 142398 393882 142634
rect 393326 106718 393562 106954
rect 393646 106718 393882 106954
rect 393326 106398 393562 106634
rect 393646 106398 393882 106634
rect 393326 70718 393562 70954
rect 393646 70718 393882 70954
rect 393326 70398 393562 70634
rect 393646 70398 393882 70634
rect 393326 34718 393562 34954
rect 393646 34718 393882 34954
rect 393326 34398 393562 34634
rect 393646 34398 393882 34634
rect 393326 -7302 393562 -7066
rect 393646 -7302 393882 -7066
rect 393326 -7622 393562 -7386
rect 393646 -7622 393882 -7386
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 402326 475718 402562 475954
rect 402646 475718 402882 475954
rect 402326 475398 402562 475634
rect 402646 475398 402882 475634
rect 402326 439718 402562 439954
rect 402646 439718 402882 439954
rect 402326 439398 402562 439634
rect 402646 439398 402882 439634
rect 402326 403718 402562 403954
rect 402646 403718 402882 403954
rect 402326 403398 402562 403634
rect 402646 403398 402882 403634
rect 402326 367718 402562 367954
rect 402646 367718 402882 367954
rect 402326 367398 402562 367634
rect 402646 367398 402882 367634
rect 402326 331718 402562 331954
rect 402646 331718 402882 331954
rect 402326 331398 402562 331634
rect 402646 331398 402882 331634
rect 402326 295718 402562 295954
rect 402646 295718 402882 295954
rect 402326 295398 402562 295634
rect 402646 295398 402882 295634
rect 402326 259718 402562 259954
rect 402646 259718 402882 259954
rect 402326 259398 402562 259634
rect 402646 259398 402882 259634
rect 402326 223718 402562 223954
rect 402646 223718 402882 223954
rect 402326 223398 402562 223634
rect 402646 223398 402882 223634
rect 402326 187718 402562 187954
rect 402646 187718 402882 187954
rect 402326 187398 402562 187634
rect 402646 187398 402882 187634
rect 402326 151718 402562 151954
rect 402646 151718 402882 151954
rect 402326 151398 402562 151634
rect 402646 151398 402882 151634
rect 402326 115718 402562 115954
rect 402646 115718 402882 115954
rect 402326 115398 402562 115634
rect 402646 115398 402882 115634
rect 402326 79718 402562 79954
rect 402646 79718 402882 79954
rect 402326 79398 402562 79634
rect 402646 79398 402882 79634
rect 402326 43718 402562 43954
rect 402646 43718 402882 43954
rect 402326 43398 402562 43634
rect 402646 43398 402882 43634
rect 406826 660218 407062 660454
rect 407146 660218 407382 660454
rect 406826 659898 407062 660134
rect 407146 659898 407382 660134
rect 406826 624218 407062 624454
rect 407146 624218 407382 624454
rect 406826 623898 407062 624134
rect 407146 623898 407382 624134
rect 406826 588218 407062 588454
rect 407146 588218 407382 588454
rect 406826 587898 407062 588134
rect 407146 587898 407382 588134
rect 406826 552218 407062 552454
rect 407146 552218 407382 552454
rect 406826 551898 407062 552134
rect 407146 551898 407382 552134
rect 406826 516218 407062 516454
rect 407146 516218 407382 516454
rect 406826 515898 407062 516134
rect 407146 515898 407382 516134
rect 406826 480218 407062 480454
rect 407146 480218 407382 480454
rect 406826 479898 407062 480134
rect 407146 479898 407382 480134
rect 406826 444218 407062 444454
rect 407146 444218 407382 444454
rect 406826 443898 407062 444134
rect 407146 443898 407382 444134
rect 406826 408218 407062 408454
rect 407146 408218 407382 408454
rect 406826 407898 407062 408134
rect 407146 407898 407382 408134
rect 406826 372218 407062 372454
rect 407146 372218 407382 372454
rect 406826 371898 407062 372134
rect 407146 371898 407382 372134
rect 406826 336218 407062 336454
rect 407146 336218 407382 336454
rect 406826 335898 407062 336134
rect 407146 335898 407382 336134
rect 406826 300218 407062 300454
rect 407146 300218 407382 300454
rect 406826 299898 407062 300134
rect 407146 299898 407382 300134
rect 406826 264218 407062 264454
rect 407146 264218 407382 264454
rect 406826 263898 407062 264134
rect 407146 263898 407382 264134
rect 406826 228218 407062 228454
rect 407146 228218 407382 228454
rect 406826 227898 407062 228134
rect 407146 227898 407382 228134
rect 406826 192218 407062 192454
rect 407146 192218 407382 192454
rect 406826 191898 407062 192134
rect 407146 191898 407382 192134
rect 406826 156218 407062 156454
rect 407146 156218 407382 156454
rect 406826 155898 407062 156134
rect 407146 155898 407382 156134
rect 406826 120218 407062 120454
rect 407146 120218 407382 120454
rect 406826 119898 407062 120134
rect 407146 119898 407382 120134
rect 406826 84218 407062 84454
rect 407146 84218 407382 84454
rect 406826 83898 407062 84134
rect 407146 83898 407382 84134
rect 406826 48218 407062 48454
rect 407146 48218 407382 48454
rect 406826 47898 407062 48134
rect 407146 47898 407382 48134
rect 402326 7718 402562 7954
rect 402646 7718 402882 7954
rect 402326 7398 402562 7634
rect 402646 7398 402882 7634
rect 402326 -1542 402562 -1306
rect 402646 -1542 402882 -1306
rect 402326 -1862 402562 -1626
rect 402646 -1862 402882 -1626
rect 406826 12218 407062 12454
rect 407146 12218 407382 12454
rect 406826 11898 407062 12134
rect 407146 11898 407382 12134
rect 406826 -2502 407062 -2266
rect 407146 -2502 407382 -2266
rect 406826 -2822 407062 -2586
rect 407146 -2822 407382 -2586
rect 411326 707482 411562 707718
rect 411646 707482 411882 707718
rect 411326 707162 411562 707398
rect 411646 707162 411882 707398
rect 411326 700718 411562 700954
rect 411646 700718 411882 700954
rect 411326 700398 411562 700634
rect 411646 700398 411882 700634
rect 411326 664718 411562 664954
rect 411646 664718 411882 664954
rect 411326 664398 411562 664634
rect 411646 664398 411882 664634
rect 411326 628718 411562 628954
rect 411646 628718 411882 628954
rect 411326 628398 411562 628634
rect 411646 628398 411882 628634
rect 411326 592718 411562 592954
rect 411646 592718 411882 592954
rect 411326 592398 411562 592634
rect 411646 592398 411882 592634
rect 411326 556718 411562 556954
rect 411646 556718 411882 556954
rect 411326 556398 411562 556634
rect 411646 556398 411882 556634
rect 411326 520718 411562 520954
rect 411646 520718 411882 520954
rect 411326 520398 411562 520634
rect 411646 520398 411882 520634
rect 411326 484718 411562 484954
rect 411646 484718 411882 484954
rect 411326 484398 411562 484634
rect 411646 484398 411882 484634
rect 411326 448718 411562 448954
rect 411646 448718 411882 448954
rect 411326 448398 411562 448634
rect 411646 448398 411882 448634
rect 411326 412718 411562 412954
rect 411646 412718 411882 412954
rect 411326 412398 411562 412634
rect 411646 412398 411882 412634
rect 411326 376718 411562 376954
rect 411646 376718 411882 376954
rect 411326 376398 411562 376634
rect 411646 376398 411882 376634
rect 411326 340718 411562 340954
rect 411646 340718 411882 340954
rect 411326 340398 411562 340634
rect 411646 340398 411882 340634
rect 411326 304718 411562 304954
rect 411646 304718 411882 304954
rect 411326 304398 411562 304634
rect 411646 304398 411882 304634
rect 411326 268718 411562 268954
rect 411646 268718 411882 268954
rect 411326 268398 411562 268634
rect 411646 268398 411882 268634
rect 411326 232718 411562 232954
rect 411646 232718 411882 232954
rect 411326 232398 411562 232634
rect 411646 232398 411882 232634
rect 411326 196718 411562 196954
rect 411646 196718 411882 196954
rect 411326 196398 411562 196634
rect 411646 196398 411882 196634
rect 411326 160718 411562 160954
rect 411646 160718 411882 160954
rect 411326 160398 411562 160634
rect 411646 160398 411882 160634
rect 411326 124718 411562 124954
rect 411646 124718 411882 124954
rect 411326 124398 411562 124634
rect 411646 124398 411882 124634
rect 411326 88718 411562 88954
rect 411646 88718 411882 88954
rect 411326 88398 411562 88634
rect 411646 88398 411882 88634
rect 411326 52718 411562 52954
rect 411646 52718 411882 52954
rect 411326 52398 411562 52634
rect 411646 52398 411882 52634
rect 411326 16718 411562 16954
rect 411646 16718 411882 16954
rect 411326 16398 411562 16634
rect 411646 16398 411882 16634
rect 411326 -3462 411562 -3226
rect 411646 -3462 411882 -3226
rect 411326 -3782 411562 -3546
rect 411646 -3782 411882 -3546
rect 415826 708442 416062 708678
rect 416146 708442 416382 708678
rect 415826 708122 416062 708358
rect 416146 708122 416382 708358
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -4422 416062 -4186
rect 416146 -4422 416382 -4186
rect 415826 -4742 416062 -4506
rect 416146 -4742 416382 -4506
rect 420326 709402 420562 709638
rect 420646 709402 420882 709638
rect 420326 709082 420562 709318
rect 420646 709082 420882 709318
rect 420326 673718 420562 673954
rect 420646 673718 420882 673954
rect 420326 673398 420562 673634
rect 420646 673398 420882 673634
rect 420326 637718 420562 637954
rect 420646 637718 420882 637954
rect 420326 637398 420562 637634
rect 420646 637398 420882 637634
rect 420326 601718 420562 601954
rect 420646 601718 420882 601954
rect 420326 601398 420562 601634
rect 420646 601398 420882 601634
rect 420326 565718 420562 565954
rect 420646 565718 420882 565954
rect 420326 565398 420562 565634
rect 420646 565398 420882 565634
rect 420326 529718 420562 529954
rect 420646 529718 420882 529954
rect 420326 529398 420562 529634
rect 420646 529398 420882 529634
rect 420326 493718 420562 493954
rect 420646 493718 420882 493954
rect 420326 493398 420562 493634
rect 420646 493398 420882 493634
rect 420326 457718 420562 457954
rect 420646 457718 420882 457954
rect 420326 457398 420562 457634
rect 420646 457398 420882 457634
rect 420326 421718 420562 421954
rect 420646 421718 420882 421954
rect 420326 421398 420562 421634
rect 420646 421398 420882 421634
rect 420326 385718 420562 385954
rect 420646 385718 420882 385954
rect 420326 385398 420562 385634
rect 420646 385398 420882 385634
rect 420326 349718 420562 349954
rect 420646 349718 420882 349954
rect 420326 349398 420562 349634
rect 420646 349398 420882 349634
rect 420326 313718 420562 313954
rect 420646 313718 420882 313954
rect 420326 313398 420562 313634
rect 420646 313398 420882 313634
rect 420326 277718 420562 277954
rect 420646 277718 420882 277954
rect 420326 277398 420562 277634
rect 420646 277398 420882 277634
rect 420326 241718 420562 241954
rect 420646 241718 420882 241954
rect 420326 241398 420562 241634
rect 420646 241398 420882 241634
rect 420326 205718 420562 205954
rect 420646 205718 420882 205954
rect 420326 205398 420562 205634
rect 420646 205398 420882 205634
rect 420326 169718 420562 169954
rect 420646 169718 420882 169954
rect 420326 169398 420562 169634
rect 420646 169398 420882 169634
rect 420326 133718 420562 133954
rect 420646 133718 420882 133954
rect 420326 133398 420562 133634
rect 420646 133398 420882 133634
rect 420326 97718 420562 97954
rect 420646 97718 420882 97954
rect 420326 97398 420562 97634
rect 420646 97398 420882 97634
rect 420326 61718 420562 61954
rect 420646 61718 420882 61954
rect 420326 61398 420562 61634
rect 420646 61398 420882 61634
rect 420326 25718 420562 25954
rect 420646 25718 420882 25954
rect 420326 25398 420562 25634
rect 420646 25398 420882 25634
rect 420326 -5382 420562 -5146
rect 420646 -5382 420882 -5146
rect 420326 -5702 420562 -5466
rect 420646 -5702 420882 -5466
rect 424826 710362 425062 710598
rect 425146 710362 425382 710598
rect 424826 710042 425062 710278
rect 425146 710042 425382 710278
rect 424826 678218 425062 678454
rect 425146 678218 425382 678454
rect 424826 677898 425062 678134
rect 425146 677898 425382 678134
rect 424826 642218 425062 642454
rect 425146 642218 425382 642454
rect 424826 641898 425062 642134
rect 425146 641898 425382 642134
rect 424826 606218 425062 606454
rect 425146 606218 425382 606454
rect 424826 605898 425062 606134
rect 425146 605898 425382 606134
rect 424826 570218 425062 570454
rect 425146 570218 425382 570454
rect 424826 569898 425062 570134
rect 425146 569898 425382 570134
rect 424826 534218 425062 534454
rect 425146 534218 425382 534454
rect 424826 533898 425062 534134
rect 425146 533898 425382 534134
rect 424826 498218 425062 498454
rect 425146 498218 425382 498454
rect 424826 497898 425062 498134
rect 425146 497898 425382 498134
rect 424826 462218 425062 462454
rect 425146 462218 425382 462454
rect 424826 461898 425062 462134
rect 425146 461898 425382 462134
rect 424826 426218 425062 426454
rect 425146 426218 425382 426454
rect 424826 425898 425062 426134
rect 425146 425898 425382 426134
rect 424826 390218 425062 390454
rect 425146 390218 425382 390454
rect 424826 389898 425062 390134
rect 425146 389898 425382 390134
rect 424826 354218 425062 354454
rect 425146 354218 425382 354454
rect 424826 353898 425062 354134
rect 425146 353898 425382 354134
rect 424826 318218 425062 318454
rect 425146 318218 425382 318454
rect 424826 317898 425062 318134
rect 425146 317898 425382 318134
rect 424826 282218 425062 282454
rect 425146 282218 425382 282454
rect 424826 281898 425062 282134
rect 425146 281898 425382 282134
rect 424826 246218 425062 246454
rect 425146 246218 425382 246454
rect 424826 245898 425062 246134
rect 425146 245898 425382 246134
rect 424826 210218 425062 210454
rect 425146 210218 425382 210454
rect 424826 209898 425062 210134
rect 425146 209898 425382 210134
rect 424826 174218 425062 174454
rect 425146 174218 425382 174454
rect 424826 173898 425062 174134
rect 425146 173898 425382 174134
rect 424826 138218 425062 138454
rect 425146 138218 425382 138454
rect 424826 137898 425062 138134
rect 425146 137898 425382 138134
rect 424826 102218 425062 102454
rect 425146 102218 425382 102454
rect 424826 101898 425062 102134
rect 425146 101898 425382 102134
rect 424826 66218 425062 66454
rect 425146 66218 425382 66454
rect 424826 65898 425062 66134
rect 425146 65898 425382 66134
rect 424826 30218 425062 30454
rect 425146 30218 425382 30454
rect 424826 29898 425062 30134
rect 425146 29898 425382 30134
rect 424826 -6342 425062 -6106
rect 425146 -6342 425382 -6106
rect 424826 -6662 425062 -6426
rect 425146 -6662 425382 -6426
rect 429326 711322 429562 711558
rect 429646 711322 429882 711558
rect 429326 711002 429562 711238
rect 429646 711002 429882 711238
rect 429326 682718 429562 682954
rect 429646 682718 429882 682954
rect 429326 682398 429562 682634
rect 429646 682398 429882 682634
rect 429326 646718 429562 646954
rect 429646 646718 429882 646954
rect 429326 646398 429562 646634
rect 429646 646398 429882 646634
rect 429326 610718 429562 610954
rect 429646 610718 429882 610954
rect 429326 610398 429562 610634
rect 429646 610398 429882 610634
rect 429326 574718 429562 574954
rect 429646 574718 429882 574954
rect 429326 574398 429562 574634
rect 429646 574398 429882 574634
rect 429326 538718 429562 538954
rect 429646 538718 429882 538954
rect 429326 538398 429562 538634
rect 429646 538398 429882 538634
rect 429326 502718 429562 502954
rect 429646 502718 429882 502954
rect 429326 502398 429562 502634
rect 429646 502398 429882 502634
rect 429326 466718 429562 466954
rect 429646 466718 429882 466954
rect 429326 466398 429562 466634
rect 429646 466398 429882 466634
rect 429326 430718 429562 430954
rect 429646 430718 429882 430954
rect 429326 430398 429562 430634
rect 429646 430398 429882 430634
rect 429326 394718 429562 394954
rect 429646 394718 429882 394954
rect 429326 394398 429562 394634
rect 429646 394398 429882 394634
rect 429326 358718 429562 358954
rect 429646 358718 429882 358954
rect 429326 358398 429562 358634
rect 429646 358398 429882 358634
rect 429326 322718 429562 322954
rect 429646 322718 429882 322954
rect 429326 322398 429562 322634
rect 429646 322398 429882 322634
rect 429326 286718 429562 286954
rect 429646 286718 429882 286954
rect 429326 286398 429562 286634
rect 429646 286398 429882 286634
rect 429326 250718 429562 250954
rect 429646 250718 429882 250954
rect 429326 250398 429562 250634
rect 429646 250398 429882 250634
rect 429326 214718 429562 214954
rect 429646 214718 429882 214954
rect 429326 214398 429562 214634
rect 429646 214398 429882 214634
rect 429326 178718 429562 178954
rect 429646 178718 429882 178954
rect 429326 178398 429562 178634
rect 429646 178398 429882 178634
rect 429326 142718 429562 142954
rect 429646 142718 429882 142954
rect 429326 142398 429562 142634
rect 429646 142398 429882 142634
rect 429326 106718 429562 106954
rect 429646 106718 429882 106954
rect 429326 106398 429562 106634
rect 429646 106398 429882 106634
rect 429326 70718 429562 70954
rect 429646 70718 429882 70954
rect 429326 70398 429562 70634
rect 429646 70398 429882 70634
rect 429326 34718 429562 34954
rect 429646 34718 429882 34954
rect 429326 34398 429562 34634
rect 429646 34398 429882 34634
rect 429326 -7302 429562 -7066
rect 429646 -7302 429882 -7066
rect 429326 -7622 429562 -7386
rect 429646 -7622 429882 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 438326 705562 438562 705798
rect 438646 705562 438882 705798
rect 438326 705242 438562 705478
rect 438646 705242 438882 705478
rect 438326 691718 438562 691954
rect 438646 691718 438882 691954
rect 438326 691398 438562 691634
rect 438646 691398 438882 691634
rect 438326 655718 438562 655954
rect 438646 655718 438882 655954
rect 438326 655398 438562 655634
rect 438646 655398 438882 655634
rect 438326 619718 438562 619954
rect 438646 619718 438882 619954
rect 438326 619398 438562 619634
rect 438646 619398 438882 619634
rect 438326 583718 438562 583954
rect 438646 583718 438882 583954
rect 438326 583398 438562 583634
rect 438646 583398 438882 583634
rect 438326 547718 438562 547954
rect 438646 547718 438882 547954
rect 438326 547398 438562 547634
rect 438646 547398 438882 547634
rect 438326 511718 438562 511954
rect 438646 511718 438882 511954
rect 438326 511398 438562 511634
rect 438646 511398 438882 511634
rect 438326 475718 438562 475954
rect 438646 475718 438882 475954
rect 438326 475398 438562 475634
rect 438646 475398 438882 475634
rect 438326 439718 438562 439954
rect 438646 439718 438882 439954
rect 438326 439398 438562 439634
rect 438646 439398 438882 439634
rect 438326 403718 438562 403954
rect 438646 403718 438882 403954
rect 438326 403398 438562 403634
rect 438646 403398 438882 403634
rect 438326 367718 438562 367954
rect 438646 367718 438882 367954
rect 438326 367398 438562 367634
rect 438646 367398 438882 367634
rect 438326 331718 438562 331954
rect 438646 331718 438882 331954
rect 438326 331398 438562 331634
rect 438646 331398 438882 331634
rect 438326 295718 438562 295954
rect 438646 295718 438882 295954
rect 438326 295398 438562 295634
rect 438646 295398 438882 295634
rect 438326 259718 438562 259954
rect 438646 259718 438882 259954
rect 438326 259398 438562 259634
rect 438646 259398 438882 259634
rect 438326 223718 438562 223954
rect 438646 223718 438882 223954
rect 438326 223398 438562 223634
rect 438646 223398 438882 223634
rect 438326 187718 438562 187954
rect 438646 187718 438882 187954
rect 438326 187398 438562 187634
rect 438646 187398 438882 187634
rect 438326 151718 438562 151954
rect 438646 151718 438882 151954
rect 438326 151398 438562 151634
rect 438646 151398 438882 151634
rect 438326 115718 438562 115954
rect 438646 115718 438882 115954
rect 438326 115398 438562 115634
rect 438646 115398 438882 115634
rect 438326 79718 438562 79954
rect 438646 79718 438882 79954
rect 438326 79398 438562 79634
rect 438646 79398 438882 79634
rect 438326 43718 438562 43954
rect 438646 43718 438882 43954
rect 438326 43398 438562 43634
rect 438646 43398 438882 43634
rect 438326 7718 438562 7954
rect 438646 7718 438882 7954
rect 438326 7398 438562 7634
rect 438646 7398 438882 7634
rect 438326 -1542 438562 -1306
rect 438646 -1542 438882 -1306
rect 438326 -1862 438562 -1626
rect 438646 -1862 438882 -1626
rect 442826 706522 443062 706758
rect 443146 706522 443382 706758
rect 442826 706202 443062 706438
rect 443146 706202 443382 706438
rect 442826 696218 443062 696454
rect 443146 696218 443382 696454
rect 442826 695898 443062 696134
rect 443146 695898 443382 696134
rect 442826 660218 443062 660454
rect 443146 660218 443382 660454
rect 442826 659898 443062 660134
rect 443146 659898 443382 660134
rect 442826 624218 443062 624454
rect 443146 624218 443382 624454
rect 442826 623898 443062 624134
rect 443146 623898 443382 624134
rect 442826 588218 443062 588454
rect 443146 588218 443382 588454
rect 442826 587898 443062 588134
rect 443146 587898 443382 588134
rect 442826 552218 443062 552454
rect 443146 552218 443382 552454
rect 442826 551898 443062 552134
rect 443146 551898 443382 552134
rect 442826 516218 443062 516454
rect 443146 516218 443382 516454
rect 442826 515898 443062 516134
rect 443146 515898 443382 516134
rect 442826 480218 443062 480454
rect 443146 480218 443382 480454
rect 442826 479898 443062 480134
rect 443146 479898 443382 480134
rect 442826 444218 443062 444454
rect 443146 444218 443382 444454
rect 442826 443898 443062 444134
rect 443146 443898 443382 444134
rect 442826 408218 443062 408454
rect 443146 408218 443382 408454
rect 442826 407898 443062 408134
rect 443146 407898 443382 408134
rect 442826 372218 443062 372454
rect 443146 372218 443382 372454
rect 442826 371898 443062 372134
rect 443146 371898 443382 372134
rect 442826 336218 443062 336454
rect 443146 336218 443382 336454
rect 442826 335898 443062 336134
rect 443146 335898 443382 336134
rect 442826 300218 443062 300454
rect 443146 300218 443382 300454
rect 442826 299898 443062 300134
rect 443146 299898 443382 300134
rect 442826 264218 443062 264454
rect 443146 264218 443382 264454
rect 442826 263898 443062 264134
rect 443146 263898 443382 264134
rect 442826 228218 443062 228454
rect 443146 228218 443382 228454
rect 442826 227898 443062 228134
rect 443146 227898 443382 228134
rect 442826 192218 443062 192454
rect 443146 192218 443382 192454
rect 442826 191898 443062 192134
rect 443146 191898 443382 192134
rect 442826 156218 443062 156454
rect 443146 156218 443382 156454
rect 442826 155898 443062 156134
rect 443146 155898 443382 156134
rect 442826 120218 443062 120454
rect 443146 120218 443382 120454
rect 442826 119898 443062 120134
rect 443146 119898 443382 120134
rect 442826 84218 443062 84454
rect 443146 84218 443382 84454
rect 442826 83898 443062 84134
rect 443146 83898 443382 84134
rect 442826 48218 443062 48454
rect 443146 48218 443382 48454
rect 442826 47898 443062 48134
rect 443146 47898 443382 48134
rect 442826 12218 443062 12454
rect 443146 12218 443382 12454
rect 442826 11898 443062 12134
rect 443146 11898 443382 12134
rect 442826 -2502 443062 -2266
rect 443146 -2502 443382 -2266
rect 442826 -2822 443062 -2586
rect 443146 -2822 443382 -2586
rect 447326 707482 447562 707718
rect 447646 707482 447882 707718
rect 447326 707162 447562 707398
rect 447646 707162 447882 707398
rect 447326 700718 447562 700954
rect 447646 700718 447882 700954
rect 447326 700398 447562 700634
rect 447646 700398 447882 700634
rect 447326 664718 447562 664954
rect 447646 664718 447882 664954
rect 447326 664398 447562 664634
rect 447646 664398 447882 664634
rect 447326 628718 447562 628954
rect 447646 628718 447882 628954
rect 447326 628398 447562 628634
rect 447646 628398 447882 628634
rect 447326 592718 447562 592954
rect 447646 592718 447882 592954
rect 447326 592398 447562 592634
rect 447646 592398 447882 592634
rect 447326 556718 447562 556954
rect 447646 556718 447882 556954
rect 447326 556398 447562 556634
rect 447646 556398 447882 556634
rect 447326 520718 447562 520954
rect 447646 520718 447882 520954
rect 447326 520398 447562 520634
rect 447646 520398 447882 520634
rect 447326 484718 447562 484954
rect 447646 484718 447882 484954
rect 447326 484398 447562 484634
rect 447646 484398 447882 484634
rect 447326 448718 447562 448954
rect 447646 448718 447882 448954
rect 447326 448398 447562 448634
rect 447646 448398 447882 448634
rect 447326 412718 447562 412954
rect 447646 412718 447882 412954
rect 447326 412398 447562 412634
rect 447646 412398 447882 412634
rect 447326 376718 447562 376954
rect 447646 376718 447882 376954
rect 447326 376398 447562 376634
rect 447646 376398 447882 376634
rect 447326 340718 447562 340954
rect 447646 340718 447882 340954
rect 447326 340398 447562 340634
rect 447646 340398 447882 340634
rect 447326 304718 447562 304954
rect 447646 304718 447882 304954
rect 447326 304398 447562 304634
rect 447646 304398 447882 304634
rect 447326 268718 447562 268954
rect 447646 268718 447882 268954
rect 447326 268398 447562 268634
rect 447646 268398 447882 268634
rect 447326 232718 447562 232954
rect 447646 232718 447882 232954
rect 447326 232398 447562 232634
rect 447646 232398 447882 232634
rect 447326 196718 447562 196954
rect 447646 196718 447882 196954
rect 447326 196398 447562 196634
rect 447646 196398 447882 196634
rect 447326 160718 447562 160954
rect 447646 160718 447882 160954
rect 447326 160398 447562 160634
rect 447646 160398 447882 160634
rect 447326 124718 447562 124954
rect 447646 124718 447882 124954
rect 447326 124398 447562 124634
rect 447646 124398 447882 124634
rect 447326 88718 447562 88954
rect 447646 88718 447882 88954
rect 447326 88398 447562 88634
rect 447646 88398 447882 88634
rect 447326 52718 447562 52954
rect 447646 52718 447882 52954
rect 447326 52398 447562 52634
rect 447646 52398 447882 52634
rect 447326 16718 447562 16954
rect 447646 16718 447882 16954
rect 447326 16398 447562 16634
rect 447646 16398 447882 16634
rect 447326 -3462 447562 -3226
rect 447646 -3462 447882 -3226
rect 447326 -3782 447562 -3546
rect 447646 -3782 447882 -3546
rect 451826 708442 452062 708678
rect 452146 708442 452382 708678
rect 451826 708122 452062 708358
rect 452146 708122 452382 708358
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -4422 452062 -4186
rect 452146 -4422 452382 -4186
rect 451826 -4742 452062 -4506
rect 452146 -4742 452382 -4506
rect 456326 709402 456562 709638
rect 456646 709402 456882 709638
rect 456326 709082 456562 709318
rect 456646 709082 456882 709318
rect 456326 673718 456562 673954
rect 456646 673718 456882 673954
rect 456326 673398 456562 673634
rect 456646 673398 456882 673634
rect 456326 637718 456562 637954
rect 456646 637718 456882 637954
rect 456326 637398 456562 637634
rect 456646 637398 456882 637634
rect 456326 601718 456562 601954
rect 456646 601718 456882 601954
rect 456326 601398 456562 601634
rect 456646 601398 456882 601634
rect 456326 565718 456562 565954
rect 456646 565718 456882 565954
rect 456326 565398 456562 565634
rect 456646 565398 456882 565634
rect 456326 529718 456562 529954
rect 456646 529718 456882 529954
rect 456326 529398 456562 529634
rect 456646 529398 456882 529634
rect 456326 493718 456562 493954
rect 456646 493718 456882 493954
rect 456326 493398 456562 493634
rect 456646 493398 456882 493634
rect 456326 457718 456562 457954
rect 456646 457718 456882 457954
rect 456326 457398 456562 457634
rect 456646 457398 456882 457634
rect 456326 421718 456562 421954
rect 456646 421718 456882 421954
rect 456326 421398 456562 421634
rect 456646 421398 456882 421634
rect 456326 385718 456562 385954
rect 456646 385718 456882 385954
rect 456326 385398 456562 385634
rect 456646 385398 456882 385634
rect 456326 349718 456562 349954
rect 456646 349718 456882 349954
rect 456326 349398 456562 349634
rect 456646 349398 456882 349634
rect 456326 313718 456562 313954
rect 456646 313718 456882 313954
rect 456326 313398 456562 313634
rect 456646 313398 456882 313634
rect 456326 277718 456562 277954
rect 456646 277718 456882 277954
rect 456326 277398 456562 277634
rect 456646 277398 456882 277634
rect 456326 241718 456562 241954
rect 456646 241718 456882 241954
rect 456326 241398 456562 241634
rect 456646 241398 456882 241634
rect 456326 205718 456562 205954
rect 456646 205718 456882 205954
rect 456326 205398 456562 205634
rect 456646 205398 456882 205634
rect 456326 169718 456562 169954
rect 456646 169718 456882 169954
rect 456326 169398 456562 169634
rect 456646 169398 456882 169634
rect 456326 133718 456562 133954
rect 456646 133718 456882 133954
rect 456326 133398 456562 133634
rect 456646 133398 456882 133634
rect 456326 97718 456562 97954
rect 456646 97718 456882 97954
rect 456326 97398 456562 97634
rect 456646 97398 456882 97634
rect 456326 61718 456562 61954
rect 456646 61718 456882 61954
rect 456326 61398 456562 61634
rect 456646 61398 456882 61634
rect 456326 25718 456562 25954
rect 456646 25718 456882 25954
rect 456326 25398 456562 25634
rect 456646 25398 456882 25634
rect 456326 -5382 456562 -5146
rect 456646 -5382 456882 -5146
rect 456326 -5702 456562 -5466
rect 456646 -5702 456882 -5466
rect 460826 710362 461062 710598
rect 461146 710362 461382 710598
rect 460826 710042 461062 710278
rect 461146 710042 461382 710278
rect 460826 678218 461062 678454
rect 461146 678218 461382 678454
rect 460826 677898 461062 678134
rect 461146 677898 461382 678134
rect 460826 642218 461062 642454
rect 461146 642218 461382 642454
rect 460826 641898 461062 642134
rect 461146 641898 461382 642134
rect 460826 606218 461062 606454
rect 461146 606218 461382 606454
rect 460826 605898 461062 606134
rect 461146 605898 461382 606134
rect 460826 570218 461062 570454
rect 461146 570218 461382 570454
rect 460826 569898 461062 570134
rect 461146 569898 461382 570134
rect 460826 534218 461062 534454
rect 461146 534218 461382 534454
rect 460826 533898 461062 534134
rect 461146 533898 461382 534134
rect 460826 498218 461062 498454
rect 461146 498218 461382 498454
rect 460826 497898 461062 498134
rect 461146 497898 461382 498134
rect 460826 462218 461062 462454
rect 461146 462218 461382 462454
rect 460826 461898 461062 462134
rect 461146 461898 461382 462134
rect 460826 426218 461062 426454
rect 461146 426218 461382 426454
rect 460826 425898 461062 426134
rect 461146 425898 461382 426134
rect 460826 390218 461062 390454
rect 461146 390218 461382 390454
rect 460826 389898 461062 390134
rect 461146 389898 461382 390134
rect 460826 354218 461062 354454
rect 461146 354218 461382 354454
rect 460826 353898 461062 354134
rect 461146 353898 461382 354134
rect 460826 318218 461062 318454
rect 461146 318218 461382 318454
rect 460826 317898 461062 318134
rect 461146 317898 461382 318134
rect 460826 282218 461062 282454
rect 461146 282218 461382 282454
rect 460826 281898 461062 282134
rect 461146 281898 461382 282134
rect 460826 246218 461062 246454
rect 461146 246218 461382 246454
rect 460826 245898 461062 246134
rect 461146 245898 461382 246134
rect 460826 210218 461062 210454
rect 461146 210218 461382 210454
rect 460826 209898 461062 210134
rect 461146 209898 461382 210134
rect 460826 174218 461062 174454
rect 461146 174218 461382 174454
rect 460826 173898 461062 174134
rect 461146 173898 461382 174134
rect 460826 138218 461062 138454
rect 461146 138218 461382 138454
rect 460826 137898 461062 138134
rect 461146 137898 461382 138134
rect 460826 102218 461062 102454
rect 461146 102218 461382 102454
rect 460826 101898 461062 102134
rect 461146 101898 461382 102134
rect 460826 66218 461062 66454
rect 461146 66218 461382 66454
rect 460826 65898 461062 66134
rect 461146 65898 461382 66134
rect 460826 30218 461062 30454
rect 461146 30218 461382 30454
rect 460826 29898 461062 30134
rect 461146 29898 461382 30134
rect 460826 -6342 461062 -6106
rect 461146 -6342 461382 -6106
rect 460826 -6662 461062 -6426
rect 461146 -6662 461382 -6426
rect 465326 711322 465562 711558
rect 465646 711322 465882 711558
rect 465326 711002 465562 711238
rect 465646 711002 465882 711238
rect 465326 682718 465562 682954
rect 465646 682718 465882 682954
rect 465326 682398 465562 682634
rect 465646 682398 465882 682634
rect 465326 646718 465562 646954
rect 465646 646718 465882 646954
rect 465326 646398 465562 646634
rect 465646 646398 465882 646634
rect 465326 610718 465562 610954
rect 465646 610718 465882 610954
rect 465326 610398 465562 610634
rect 465646 610398 465882 610634
rect 465326 574718 465562 574954
rect 465646 574718 465882 574954
rect 465326 574398 465562 574634
rect 465646 574398 465882 574634
rect 465326 538718 465562 538954
rect 465646 538718 465882 538954
rect 465326 538398 465562 538634
rect 465646 538398 465882 538634
rect 465326 502718 465562 502954
rect 465646 502718 465882 502954
rect 465326 502398 465562 502634
rect 465646 502398 465882 502634
rect 465326 466718 465562 466954
rect 465646 466718 465882 466954
rect 465326 466398 465562 466634
rect 465646 466398 465882 466634
rect 465326 430718 465562 430954
rect 465646 430718 465882 430954
rect 465326 430398 465562 430634
rect 465646 430398 465882 430634
rect 465326 394718 465562 394954
rect 465646 394718 465882 394954
rect 465326 394398 465562 394634
rect 465646 394398 465882 394634
rect 465326 358718 465562 358954
rect 465646 358718 465882 358954
rect 465326 358398 465562 358634
rect 465646 358398 465882 358634
rect 465326 322718 465562 322954
rect 465646 322718 465882 322954
rect 465326 322398 465562 322634
rect 465646 322398 465882 322634
rect 465326 286718 465562 286954
rect 465646 286718 465882 286954
rect 465326 286398 465562 286634
rect 465646 286398 465882 286634
rect 465326 250718 465562 250954
rect 465646 250718 465882 250954
rect 465326 250398 465562 250634
rect 465646 250398 465882 250634
rect 465326 214718 465562 214954
rect 465646 214718 465882 214954
rect 465326 214398 465562 214634
rect 465646 214398 465882 214634
rect 465326 178718 465562 178954
rect 465646 178718 465882 178954
rect 465326 178398 465562 178634
rect 465646 178398 465882 178634
rect 465326 142718 465562 142954
rect 465646 142718 465882 142954
rect 465326 142398 465562 142634
rect 465646 142398 465882 142634
rect 465326 106718 465562 106954
rect 465646 106718 465882 106954
rect 465326 106398 465562 106634
rect 465646 106398 465882 106634
rect 465326 70718 465562 70954
rect 465646 70718 465882 70954
rect 465326 70398 465562 70634
rect 465646 70398 465882 70634
rect 465326 34718 465562 34954
rect 465646 34718 465882 34954
rect 465326 34398 465562 34634
rect 465646 34398 465882 34634
rect 465326 -7302 465562 -7066
rect 465646 -7302 465882 -7066
rect 465326 -7622 465562 -7386
rect 465646 -7622 465882 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 474326 705562 474562 705798
rect 474646 705562 474882 705798
rect 474326 705242 474562 705478
rect 474646 705242 474882 705478
rect 474326 691718 474562 691954
rect 474646 691718 474882 691954
rect 474326 691398 474562 691634
rect 474646 691398 474882 691634
rect 474326 655718 474562 655954
rect 474646 655718 474882 655954
rect 474326 655398 474562 655634
rect 474646 655398 474882 655634
rect 478826 706522 479062 706758
rect 479146 706522 479382 706758
rect 478826 706202 479062 706438
rect 479146 706202 479382 706438
rect 478826 696218 479062 696454
rect 479146 696218 479382 696454
rect 478826 695898 479062 696134
rect 479146 695898 479382 696134
rect 478826 660218 479062 660454
rect 479146 660218 479382 660454
rect 478826 659898 479062 660134
rect 479146 659898 479382 660134
rect 483326 707482 483562 707718
rect 483646 707482 483882 707718
rect 483326 707162 483562 707398
rect 483646 707162 483882 707398
rect 483326 700718 483562 700954
rect 483646 700718 483882 700954
rect 483326 700398 483562 700634
rect 483646 700398 483882 700634
rect 483326 664718 483562 664954
rect 483646 664718 483882 664954
rect 483326 664398 483562 664634
rect 483646 664398 483882 664634
rect 487826 708442 488062 708678
rect 488146 708442 488382 708678
rect 487826 708122 488062 708358
rect 488146 708122 488382 708358
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 492326 709402 492562 709638
rect 492646 709402 492882 709638
rect 492326 709082 492562 709318
rect 492646 709082 492882 709318
rect 492326 673718 492562 673954
rect 492646 673718 492882 673954
rect 492326 673398 492562 673634
rect 492646 673398 492882 673634
rect 474326 619718 474562 619954
rect 474646 619718 474882 619954
rect 474326 619398 474562 619634
rect 474646 619398 474882 619634
rect 484250 615218 484486 615454
rect 484250 614898 484486 615134
rect 474326 583718 474562 583954
rect 474646 583718 474882 583954
rect 474326 583398 474562 583634
rect 474646 583398 474882 583634
rect 474326 547718 474562 547954
rect 474646 547718 474882 547954
rect 474326 547398 474562 547634
rect 474646 547398 474882 547634
rect 478826 588218 479062 588454
rect 479146 588218 479382 588454
rect 478826 587898 479062 588134
rect 479146 587898 479382 588134
rect 478826 552218 479062 552454
rect 479146 552218 479382 552454
rect 478826 551898 479062 552134
rect 479146 551898 479382 552134
rect 483326 592718 483562 592954
rect 483646 592718 483882 592954
rect 483326 592398 483562 592634
rect 483646 592398 483882 592634
rect 483326 556718 483562 556954
rect 483646 556718 483882 556954
rect 483326 556398 483562 556634
rect 483646 556398 483882 556634
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 496826 710362 497062 710598
rect 497146 710362 497382 710598
rect 496826 710042 497062 710278
rect 497146 710042 497382 710278
rect 496826 678218 497062 678454
rect 497146 678218 497382 678454
rect 496826 677898 497062 678134
rect 497146 677898 497382 678134
rect 496826 642125 497062 642361
rect 497146 642125 497382 642361
rect 501326 711322 501562 711558
rect 501646 711322 501882 711558
rect 501326 711002 501562 711238
rect 501646 711002 501882 711238
rect 501326 682718 501562 682954
rect 501646 682718 501882 682954
rect 501326 682398 501562 682634
rect 501646 682398 501882 682634
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 501326 646718 501562 646954
rect 501646 646718 501882 646954
rect 501326 646398 501562 646634
rect 501646 646398 501882 646634
rect 499610 619718 499846 619954
rect 499610 619398 499846 619634
rect 474326 511718 474562 511954
rect 474646 511718 474882 511954
rect 474326 511398 474562 511634
rect 474646 511398 474882 511634
rect 484250 507218 484486 507454
rect 484250 506898 484486 507134
rect 474326 475718 474562 475954
rect 474646 475718 474882 475954
rect 474326 475398 474562 475634
rect 474646 475398 474882 475634
rect 474326 439718 474562 439954
rect 474646 439718 474882 439954
rect 474326 439398 474562 439634
rect 474646 439398 474882 439634
rect 474326 403718 474562 403954
rect 474646 403718 474882 403954
rect 474326 403398 474562 403634
rect 474646 403398 474882 403634
rect 474326 367718 474562 367954
rect 474646 367718 474882 367954
rect 474326 367398 474562 367634
rect 474646 367398 474882 367634
rect 474326 331718 474562 331954
rect 474646 331718 474882 331954
rect 474326 331398 474562 331634
rect 474646 331398 474882 331634
rect 474326 295718 474562 295954
rect 474646 295718 474882 295954
rect 474326 295398 474562 295634
rect 474646 295398 474882 295634
rect 474326 259718 474562 259954
rect 474646 259718 474882 259954
rect 474326 259398 474562 259634
rect 474646 259398 474882 259634
rect 474326 223718 474562 223954
rect 474646 223718 474882 223954
rect 474326 223398 474562 223634
rect 474646 223398 474882 223634
rect 474326 187718 474562 187954
rect 474646 187718 474882 187954
rect 474326 187398 474562 187634
rect 474646 187398 474882 187634
rect 474326 151718 474562 151954
rect 474646 151718 474882 151954
rect 474326 151398 474562 151634
rect 474646 151398 474882 151634
rect 474326 115718 474562 115954
rect 474646 115718 474882 115954
rect 474326 115398 474562 115634
rect 474646 115398 474882 115634
rect 474326 79718 474562 79954
rect 474646 79718 474882 79954
rect 474326 79398 474562 79634
rect 474646 79398 474882 79634
rect 474326 43718 474562 43954
rect 474646 43718 474882 43954
rect 474326 43398 474562 43634
rect 474646 43398 474882 43634
rect 474326 7718 474562 7954
rect 474646 7718 474882 7954
rect 474326 7398 474562 7634
rect 474646 7398 474882 7634
rect 474326 -1542 474562 -1306
rect 474646 -1542 474882 -1306
rect 474326 -1862 474562 -1626
rect 474646 -1862 474882 -1626
rect 478826 480218 479062 480454
rect 479146 480218 479382 480454
rect 478826 479898 479062 480134
rect 479146 479898 479382 480134
rect 478826 444218 479062 444454
rect 479146 444218 479382 444454
rect 478826 443898 479062 444134
rect 479146 443898 479382 444134
rect 478826 408218 479062 408454
rect 479146 408218 479382 408454
rect 478826 407898 479062 408134
rect 479146 407898 479382 408134
rect 478826 372218 479062 372454
rect 479146 372218 479382 372454
rect 478826 371898 479062 372134
rect 479146 371898 479382 372134
rect 478826 336218 479062 336454
rect 479146 336218 479382 336454
rect 478826 335898 479062 336134
rect 479146 335898 479382 336134
rect 478826 300218 479062 300454
rect 479146 300218 479382 300454
rect 478826 299898 479062 300134
rect 479146 299898 479382 300134
rect 478826 264218 479062 264454
rect 479146 264218 479382 264454
rect 478826 263898 479062 264134
rect 479146 263898 479382 264134
rect 478826 228218 479062 228454
rect 479146 228218 479382 228454
rect 478826 227898 479062 228134
rect 479146 227898 479382 228134
rect 478826 192218 479062 192454
rect 479146 192218 479382 192454
rect 478826 191898 479062 192134
rect 479146 191898 479382 192134
rect 478826 156218 479062 156454
rect 479146 156218 479382 156454
rect 478826 155898 479062 156134
rect 479146 155898 479382 156134
rect 478826 120218 479062 120454
rect 479146 120218 479382 120454
rect 478826 119898 479062 120134
rect 479146 119898 479382 120134
rect 478826 84218 479062 84454
rect 479146 84218 479382 84454
rect 478826 83898 479062 84134
rect 479146 83898 479382 84134
rect 478826 48218 479062 48454
rect 479146 48218 479382 48454
rect 478826 47898 479062 48134
rect 479146 47898 479382 48134
rect 478826 12218 479062 12454
rect 479146 12218 479382 12454
rect 478826 11898 479062 12134
rect 479146 11898 479382 12134
rect 478826 -2502 479062 -2266
rect 479146 -2502 479382 -2266
rect 478826 -2822 479062 -2586
rect 479146 -2822 479382 -2586
rect 483326 484718 483562 484954
rect 483646 484718 483882 484954
rect 483326 484398 483562 484634
rect 483646 484398 483882 484634
rect 483326 448718 483562 448954
rect 483646 448718 483882 448954
rect 483326 448398 483562 448634
rect 483646 448398 483882 448634
rect 483326 412718 483562 412954
rect 483646 412718 483882 412954
rect 483326 412398 483562 412634
rect 483646 412398 483882 412634
rect 483326 376718 483562 376954
rect 483646 376718 483882 376954
rect 483326 376398 483562 376634
rect 483646 376398 483882 376634
rect 483326 340718 483562 340954
rect 483646 340718 483882 340954
rect 483326 340398 483562 340634
rect 483646 340398 483882 340634
rect 483326 304718 483562 304954
rect 483646 304718 483882 304954
rect 483326 304398 483562 304634
rect 483646 304398 483882 304634
rect 483326 268718 483562 268954
rect 483646 268718 483882 268954
rect 483326 268398 483562 268634
rect 483646 268398 483882 268634
rect 483326 232718 483562 232954
rect 483646 232718 483882 232954
rect 483326 232398 483562 232634
rect 483646 232398 483882 232634
rect 483326 196718 483562 196954
rect 483646 196718 483882 196954
rect 483326 196398 483562 196634
rect 483646 196398 483882 196634
rect 483326 160718 483562 160954
rect 483646 160718 483882 160954
rect 483326 160398 483562 160634
rect 483646 160398 483882 160634
rect 483326 124718 483562 124954
rect 483646 124718 483882 124954
rect 483326 124398 483562 124634
rect 483646 124398 483882 124634
rect 483326 88718 483562 88954
rect 483646 88718 483882 88954
rect 483326 88398 483562 88634
rect 483646 88398 483882 88634
rect 483326 52718 483562 52954
rect 483646 52718 483882 52954
rect 483326 52398 483562 52634
rect 483646 52398 483882 52634
rect 483326 16718 483562 16954
rect 483646 16718 483882 16954
rect 483326 16398 483562 16634
rect 483646 16398 483882 16634
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 483326 -3462 483562 -3226
rect 483646 -3462 483882 -3226
rect 483326 -3782 483562 -3546
rect 483646 -3782 483882 -3546
rect 487826 -4422 488062 -4186
rect 488146 -4422 488382 -4186
rect 487826 -4742 488062 -4506
rect 488146 -4742 488382 -4506
rect 492326 493718 492562 493954
rect 492646 493718 492882 493954
rect 492326 493398 492562 493634
rect 492646 493398 492882 493634
rect 492326 457718 492562 457954
rect 492646 457718 492882 457954
rect 492326 457398 492562 457634
rect 492646 457398 492882 457634
rect 492326 421718 492562 421954
rect 492646 421718 492882 421954
rect 492326 421398 492562 421634
rect 492646 421398 492882 421634
rect 492326 385718 492562 385954
rect 492646 385718 492882 385954
rect 492326 385398 492562 385634
rect 492646 385398 492882 385634
rect 492326 349718 492562 349954
rect 492646 349718 492882 349954
rect 492326 349398 492562 349634
rect 492646 349398 492882 349634
rect 492326 313718 492562 313954
rect 492646 313718 492882 313954
rect 492326 313398 492562 313634
rect 492646 313398 492882 313634
rect 492326 277718 492562 277954
rect 492646 277718 492882 277954
rect 492326 277398 492562 277634
rect 492646 277398 492882 277634
rect 492326 241718 492562 241954
rect 492646 241718 492882 241954
rect 492326 241398 492562 241634
rect 492646 241398 492882 241634
rect 492326 205718 492562 205954
rect 492646 205718 492882 205954
rect 492326 205398 492562 205634
rect 492646 205398 492882 205634
rect 492326 169718 492562 169954
rect 492646 169718 492882 169954
rect 492326 169398 492562 169634
rect 492646 169398 492882 169634
rect 492326 133718 492562 133954
rect 492646 133718 492882 133954
rect 492326 133398 492562 133634
rect 492646 133398 492882 133634
rect 492326 97718 492562 97954
rect 492646 97718 492882 97954
rect 492326 97398 492562 97634
rect 492646 97398 492882 97634
rect 492326 61718 492562 61954
rect 492646 61718 492882 61954
rect 492326 61398 492562 61634
rect 492646 61398 492882 61634
rect 492326 25718 492562 25954
rect 492646 25718 492882 25954
rect 492326 25398 492562 25634
rect 492646 25398 492882 25634
rect 499610 511718 499846 511954
rect 499610 511398 499846 511634
rect 496826 462218 497062 462454
rect 497146 462218 497382 462454
rect 496826 461898 497062 462134
rect 497146 461898 497382 462134
rect 496826 426218 497062 426454
rect 497146 426218 497382 426454
rect 496826 425898 497062 426134
rect 497146 425898 497382 426134
rect 496826 390218 497062 390454
rect 497146 390218 497382 390454
rect 496826 389898 497062 390134
rect 497146 389898 497382 390134
rect 496826 354218 497062 354454
rect 497146 354218 497382 354454
rect 496826 353898 497062 354134
rect 497146 353898 497382 354134
rect 496826 318218 497062 318454
rect 497146 318218 497382 318454
rect 496826 317898 497062 318134
rect 497146 317898 497382 318134
rect 496826 282218 497062 282454
rect 497146 282218 497382 282454
rect 496826 281898 497062 282134
rect 497146 281898 497382 282134
rect 496826 246218 497062 246454
rect 497146 246218 497382 246454
rect 496826 245898 497062 246134
rect 497146 245898 497382 246134
rect 496826 210218 497062 210454
rect 497146 210218 497382 210454
rect 496826 209898 497062 210134
rect 497146 209898 497382 210134
rect 496826 174218 497062 174454
rect 497146 174218 497382 174454
rect 496826 173898 497062 174134
rect 497146 173898 497382 174134
rect 496826 138218 497062 138454
rect 497146 138218 497382 138454
rect 496826 137898 497062 138134
rect 497146 137898 497382 138134
rect 496826 102218 497062 102454
rect 497146 102218 497382 102454
rect 496826 101898 497062 102134
rect 497146 101898 497382 102134
rect 496826 66218 497062 66454
rect 497146 66218 497382 66454
rect 496826 65898 497062 66134
rect 497146 65898 497382 66134
rect 496826 30218 497062 30454
rect 497146 30218 497382 30454
rect 496826 29898 497062 30134
rect 497146 29898 497382 30134
rect 492326 -5382 492562 -5146
rect 492646 -5382 492882 -5146
rect 492326 -5702 492562 -5466
rect 492646 -5702 492882 -5466
rect 496826 -6342 497062 -6106
rect 497146 -6342 497382 -6106
rect 496826 -6662 497062 -6426
rect 497146 -6662 497382 -6426
rect 501326 466718 501562 466954
rect 501646 466718 501882 466954
rect 501326 466398 501562 466634
rect 501646 466398 501882 466634
rect 501326 430718 501562 430954
rect 501646 430718 501882 430954
rect 501326 430398 501562 430634
rect 501646 430398 501882 430634
rect 501326 394718 501562 394954
rect 501646 394718 501882 394954
rect 501326 394398 501562 394634
rect 501646 394398 501882 394634
rect 501326 358718 501562 358954
rect 501646 358718 501882 358954
rect 501326 358398 501562 358634
rect 501646 358398 501882 358634
rect 501326 322718 501562 322954
rect 501646 322718 501882 322954
rect 501326 322398 501562 322634
rect 501646 322398 501882 322634
rect 501326 286718 501562 286954
rect 501646 286718 501882 286954
rect 501326 286398 501562 286634
rect 501646 286398 501882 286634
rect 501326 250718 501562 250954
rect 501646 250718 501882 250954
rect 501326 250398 501562 250634
rect 501646 250398 501882 250634
rect 501326 214718 501562 214954
rect 501646 214718 501882 214954
rect 501326 214398 501562 214634
rect 501646 214398 501882 214634
rect 501326 178718 501562 178954
rect 501646 178718 501882 178954
rect 501326 178398 501562 178634
rect 501646 178398 501882 178634
rect 501326 142718 501562 142954
rect 501646 142718 501882 142954
rect 501326 142398 501562 142634
rect 501646 142398 501882 142634
rect 501326 106718 501562 106954
rect 501646 106718 501882 106954
rect 501326 106398 501562 106634
rect 501646 106398 501882 106634
rect 501326 70718 501562 70954
rect 501646 70718 501882 70954
rect 501326 70398 501562 70634
rect 501646 70398 501882 70634
rect 501326 34718 501562 34954
rect 501646 34718 501882 34954
rect 501326 34398 501562 34634
rect 501646 34398 501882 34634
rect 510326 705562 510562 705798
rect 510646 705562 510882 705798
rect 510326 705242 510562 705478
rect 510646 705242 510882 705478
rect 510326 691718 510562 691954
rect 510646 691718 510882 691954
rect 510326 691398 510562 691634
rect 510646 691398 510882 691634
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 510326 655718 510562 655954
rect 510646 655718 510882 655954
rect 510326 655398 510562 655634
rect 510646 655398 510882 655634
rect 514826 706522 515062 706758
rect 515146 706522 515382 706758
rect 514826 706202 515062 706438
rect 515146 706202 515382 706438
rect 514826 696218 515062 696454
rect 515146 696218 515382 696454
rect 514826 695898 515062 696134
rect 515146 695898 515382 696134
rect 514826 660218 515062 660454
rect 515146 660218 515382 660454
rect 514826 659898 515062 660134
rect 515146 659898 515382 660134
rect 519326 707482 519562 707718
rect 519646 707482 519882 707718
rect 519326 707162 519562 707398
rect 519646 707162 519882 707398
rect 519326 700718 519562 700954
rect 519646 700718 519882 700954
rect 519326 700398 519562 700634
rect 519646 700398 519882 700634
rect 519326 664718 519562 664954
rect 519646 664718 519882 664954
rect 519326 664398 519562 664634
rect 519646 664398 519882 664634
rect 523826 708442 524062 708678
rect 524146 708442 524382 708678
rect 523826 708122 524062 708358
rect 524146 708122 524382 708358
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 528326 709402 528562 709638
rect 528646 709402 528882 709638
rect 528326 709082 528562 709318
rect 528646 709082 528882 709318
rect 528326 673718 528562 673954
rect 528646 673718 528882 673954
rect 528326 673398 528562 673634
rect 528646 673398 528882 673634
rect 528326 637718 528562 637954
rect 528646 637718 528882 637954
rect 528326 637398 528562 637634
rect 528646 637398 528882 637634
rect 514970 615218 515206 615454
rect 514970 614898 515206 615134
rect 528326 601718 528562 601954
rect 528646 601718 528882 601954
rect 528326 601398 528562 601634
rect 528646 601398 528882 601634
rect 510326 583718 510562 583954
rect 510646 583718 510882 583954
rect 510326 583398 510562 583634
rect 510646 583398 510882 583634
rect 510326 547718 510562 547954
rect 510646 547718 510882 547954
rect 510326 547398 510562 547634
rect 510646 547398 510882 547634
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 514826 588218 515062 588454
rect 515146 588218 515382 588454
rect 514826 587898 515062 588134
rect 515146 587898 515382 588134
rect 514826 552218 515062 552454
rect 515146 552218 515382 552454
rect 514826 551898 515062 552134
rect 515146 551898 515382 552134
rect 519326 592718 519562 592954
rect 519646 592718 519882 592954
rect 519326 592398 519562 592634
rect 519646 592398 519882 592634
rect 519326 556718 519562 556954
rect 519646 556718 519882 556954
rect 519326 556398 519562 556634
rect 519646 556398 519882 556634
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 528326 565718 528562 565954
rect 528646 565718 528882 565954
rect 528326 565398 528562 565634
rect 528646 565398 528882 565634
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 501326 -7302 501562 -7066
rect 501646 -7302 501882 -7066
rect 501326 -7622 501562 -7386
rect 501646 -7622 501882 -7386
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 510326 475718 510562 475954
rect 510646 475718 510882 475954
rect 510326 475398 510562 475634
rect 510646 475398 510882 475634
rect 510326 439718 510562 439954
rect 510646 439718 510882 439954
rect 510326 439398 510562 439634
rect 510646 439398 510882 439634
rect 510326 403718 510562 403954
rect 510646 403718 510882 403954
rect 510326 403398 510562 403634
rect 510646 403398 510882 403634
rect 510326 367718 510562 367954
rect 510646 367718 510882 367954
rect 510326 367398 510562 367634
rect 510646 367398 510882 367634
rect 510326 331718 510562 331954
rect 510646 331718 510882 331954
rect 510326 331398 510562 331634
rect 510646 331398 510882 331634
rect 510326 295718 510562 295954
rect 510646 295718 510882 295954
rect 510326 295398 510562 295634
rect 510646 295398 510882 295634
rect 510326 259718 510562 259954
rect 510646 259718 510882 259954
rect 510326 259398 510562 259634
rect 510646 259398 510882 259634
rect 510326 223718 510562 223954
rect 510646 223718 510882 223954
rect 510326 223398 510562 223634
rect 510646 223398 510882 223634
rect 510326 187718 510562 187954
rect 510646 187718 510882 187954
rect 510326 187398 510562 187634
rect 510646 187398 510882 187634
rect 510326 151718 510562 151954
rect 510646 151718 510882 151954
rect 510326 151398 510562 151634
rect 510646 151398 510882 151634
rect 510326 115718 510562 115954
rect 510646 115718 510882 115954
rect 510326 115398 510562 115634
rect 510646 115398 510882 115634
rect 510326 79718 510562 79954
rect 510646 79718 510882 79954
rect 510326 79398 510562 79634
rect 510646 79398 510882 79634
rect 510326 43718 510562 43954
rect 510646 43718 510882 43954
rect 510326 43398 510562 43634
rect 510646 43398 510882 43634
rect 510326 7718 510562 7954
rect 510646 7718 510882 7954
rect 510326 7398 510562 7634
rect 510646 7398 510882 7634
rect 514970 507218 515206 507454
rect 514970 506898 515206 507134
rect 514826 480218 515062 480454
rect 515146 480218 515382 480454
rect 514826 479898 515062 480134
rect 515146 479898 515382 480134
rect 514826 444218 515062 444454
rect 515146 444218 515382 444454
rect 514826 443898 515062 444134
rect 515146 443898 515382 444134
rect 514826 408218 515062 408454
rect 515146 408218 515382 408454
rect 514826 407898 515062 408134
rect 515146 407898 515382 408134
rect 514826 372218 515062 372454
rect 515146 372218 515382 372454
rect 514826 371898 515062 372134
rect 515146 371898 515382 372134
rect 514826 336218 515062 336454
rect 515146 336218 515382 336454
rect 514826 335898 515062 336134
rect 515146 335898 515382 336134
rect 514826 300218 515062 300454
rect 515146 300218 515382 300454
rect 514826 299898 515062 300134
rect 515146 299898 515382 300134
rect 514826 264218 515062 264454
rect 515146 264218 515382 264454
rect 514826 263898 515062 264134
rect 515146 263898 515382 264134
rect 514826 228218 515062 228454
rect 515146 228218 515382 228454
rect 514826 227898 515062 228134
rect 515146 227898 515382 228134
rect 514826 192218 515062 192454
rect 515146 192218 515382 192454
rect 514826 191898 515062 192134
rect 515146 191898 515382 192134
rect 514826 156218 515062 156454
rect 515146 156218 515382 156454
rect 514826 155898 515062 156134
rect 515146 155898 515382 156134
rect 514826 120218 515062 120454
rect 515146 120218 515382 120454
rect 514826 119898 515062 120134
rect 515146 119898 515382 120134
rect 514826 84218 515062 84454
rect 515146 84218 515382 84454
rect 514826 83898 515062 84134
rect 515146 83898 515382 84134
rect 514826 48218 515062 48454
rect 515146 48218 515382 48454
rect 514826 47898 515062 48134
rect 515146 47898 515382 48134
rect 514826 12218 515062 12454
rect 515146 12218 515382 12454
rect 514826 11898 515062 12134
rect 515146 11898 515382 12134
rect 510326 -1542 510562 -1306
rect 510646 -1542 510882 -1306
rect 510326 -1862 510562 -1626
rect 510646 -1862 510882 -1626
rect 519326 484718 519562 484954
rect 519646 484718 519882 484954
rect 519326 484398 519562 484634
rect 519646 484398 519882 484634
rect 519326 448718 519562 448954
rect 519646 448718 519882 448954
rect 519326 448398 519562 448634
rect 519646 448398 519882 448634
rect 519326 412718 519562 412954
rect 519646 412718 519882 412954
rect 519326 412398 519562 412634
rect 519646 412398 519882 412634
rect 519326 376718 519562 376954
rect 519646 376718 519882 376954
rect 519326 376398 519562 376634
rect 519646 376398 519882 376634
rect 519326 340718 519562 340954
rect 519646 340718 519882 340954
rect 519326 340398 519562 340634
rect 519646 340398 519882 340634
rect 519326 304718 519562 304954
rect 519646 304718 519882 304954
rect 519326 304398 519562 304634
rect 519646 304398 519882 304634
rect 519326 268718 519562 268954
rect 519646 268718 519882 268954
rect 519326 268398 519562 268634
rect 519646 268398 519882 268634
rect 519326 232718 519562 232954
rect 519646 232718 519882 232954
rect 519326 232398 519562 232634
rect 519646 232398 519882 232634
rect 519326 196718 519562 196954
rect 519646 196718 519882 196954
rect 519326 196398 519562 196634
rect 519646 196398 519882 196634
rect 519326 160718 519562 160954
rect 519646 160718 519882 160954
rect 519326 160398 519562 160634
rect 519646 160398 519882 160634
rect 519326 124718 519562 124954
rect 519646 124718 519882 124954
rect 519326 124398 519562 124634
rect 519646 124398 519882 124634
rect 519326 88718 519562 88954
rect 519646 88718 519882 88954
rect 519326 88398 519562 88634
rect 519646 88398 519882 88634
rect 519326 52718 519562 52954
rect 519646 52718 519882 52954
rect 519326 52398 519562 52634
rect 519646 52398 519882 52634
rect 519326 16718 519562 16954
rect 519646 16718 519882 16954
rect 519326 16398 519562 16634
rect 519646 16398 519882 16634
rect 514826 -2502 515062 -2266
rect 515146 -2502 515382 -2266
rect 514826 -2822 515062 -2586
rect 515146 -2822 515382 -2586
rect 528326 529718 528562 529954
rect 528646 529718 528882 529954
rect 528326 529398 528562 529634
rect 528646 529398 528882 529634
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 519326 -3462 519562 -3226
rect 519646 -3462 519882 -3226
rect 519326 -3782 519562 -3546
rect 519646 -3782 519882 -3546
rect 523826 -4422 524062 -4186
rect 524146 -4422 524382 -4186
rect 523826 -4742 524062 -4506
rect 524146 -4742 524382 -4506
rect 528326 493718 528562 493954
rect 528646 493718 528882 493954
rect 528326 493398 528562 493634
rect 528646 493398 528882 493634
rect 528326 457718 528562 457954
rect 528646 457718 528882 457954
rect 528326 457398 528562 457634
rect 528646 457398 528882 457634
rect 528326 421718 528562 421954
rect 528646 421718 528882 421954
rect 528326 421398 528562 421634
rect 528646 421398 528882 421634
rect 528326 385718 528562 385954
rect 528646 385718 528882 385954
rect 528326 385398 528562 385634
rect 528646 385398 528882 385634
rect 528326 349718 528562 349954
rect 528646 349718 528882 349954
rect 528326 349398 528562 349634
rect 528646 349398 528882 349634
rect 528326 313718 528562 313954
rect 528646 313718 528882 313954
rect 528326 313398 528562 313634
rect 528646 313398 528882 313634
rect 528326 277718 528562 277954
rect 528646 277718 528882 277954
rect 528326 277398 528562 277634
rect 528646 277398 528882 277634
rect 528326 241718 528562 241954
rect 528646 241718 528882 241954
rect 528326 241398 528562 241634
rect 528646 241398 528882 241634
rect 528326 205718 528562 205954
rect 528646 205718 528882 205954
rect 528326 205398 528562 205634
rect 528646 205398 528882 205634
rect 528326 169718 528562 169954
rect 528646 169718 528882 169954
rect 528326 169398 528562 169634
rect 528646 169398 528882 169634
rect 528326 133718 528562 133954
rect 528646 133718 528882 133954
rect 528326 133398 528562 133634
rect 528646 133398 528882 133634
rect 528326 97718 528562 97954
rect 528646 97718 528882 97954
rect 528326 97398 528562 97634
rect 528646 97398 528882 97634
rect 528326 61718 528562 61954
rect 528646 61718 528882 61954
rect 528326 61398 528562 61634
rect 528646 61398 528882 61634
rect 528326 25718 528562 25954
rect 528646 25718 528882 25954
rect 528326 25398 528562 25634
rect 528646 25398 528882 25634
rect 528326 -5382 528562 -5146
rect 528646 -5382 528882 -5146
rect 528326 -5702 528562 -5466
rect 528646 -5702 528882 -5466
rect 532826 710362 533062 710598
rect 533146 710362 533382 710598
rect 532826 710042 533062 710278
rect 533146 710042 533382 710278
rect 532826 678218 533062 678454
rect 533146 678218 533382 678454
rect 532826 677898 533062 678134
rect 533146 677898 533382 678134
rect 532826 642218 533062 642454
rect 533146 642218 533382 642454
rect 532826 641898 533062 642134
rect 533146 641898 533382 642134
rect 532826 606218 533062 606454
rect 533146 606218 533382 606454
rect 532826 605898 533062 606134
rect 533146 605898 533382 606134
rect 532826 570218 533062 570454
rect 533146 570218 533382 570454
rect 532826 569898 533062 570134
rect 533146 569898 533382 570134
rect 532826 534218 533062 534454
rect 533146 534218 533382 534454
rect 532826 533898 533062 534134
rect 533146 533898 533382 534134
rect 532826 498218 533062 498454
rect 533146 498218 533382 498454
rect 532826 497898 533062 498134
rect 533146 497898 533382 498134
rect 532826 462218 533062 462454
rect 533146 462218 533382 462454
rect 532826 461898 533062 462134
rect 533146 461898 533382 462134
rect 532826 426218 533062 426454
rect 533146 426218 533382 426454
rect 532826 425898 533062 426134
rect 533146 425898 533382 426134
rect 532826 390218 533062 390454
rect 533146 390218 533382 390454
rect 532826 389898 533062 390134
rect 533146 389898 533382 390134
rect 532826 354218 533062 354454
rect 533146 354218 533382 354454
rect 532826 353898 533062 354134
rect 533146 353898 533382 354134
rect 532826 318218 533062 318454
rect 533146 318218 533382 318454
rect 532826 317898 533062 318134
rect 533146 317898 533382 318134
rect 532826 282218 533062 282454
rect 533146 282218 533382 282454
rect 532826 281898 533062 282134
rect 533146 281898 533382 282134
rect 532826 246218 533062 246454
rect 533146 246218 533382 246454
rect 532826 245898 533062 246134
rect 533146 245898 533382 246134
rect 532826 210218 533062 210454
rect 533146 210218 533382 210454
rect 532826 209898 533062 210134
rect 533146 209898 533382 210134
rect 532826 174218 533062 174454
rect 533146 174218 533382 174454
rect 532826 173898 533062 174134
rect 533146 173898 533382 174134
rect 532826 138218 533062 138454
rect 533146 138218 533382 138454
rect 532826 137898 533062 138134
rect 533146 137898 533382 138134
rect 532826 102218 533062 102454
rect 533146 102218 533382 102454
rect 532826 101898 533062 102134
rect 533146 101898 533382 102134
rect 532826 66218 533062 66454
rect 533146 66218 533382 66454
rect 532826 65898 533062 66134
rect 533146 65898 533382 66134
rect 532826 30218 533062 30454
rect 533146 30218 533382 30454
rect 532826 29898 533062 30134
rect 533146 29898 533382 30134
rect 532826 -6342 533062 -6106
rect 533146 -6342 533382 -6106
rect 532826 -6662 533062 -6426
rect 533146 -6662 533382 -6426
rect 537326 711322 537562 711558
rect 537646 711322 537882 711558
rect 537326 711002 537562 711238
rect 537646 711002 537882 711238
rect 537326 682718 537562 682954
rect 537646 682718 537882 682954
rect 537326 682398 537562 682634
rect 537646 682398 537882 682634
rect 537326 646718 537562 646954
rect 537646 646718 537882 646954
rect 537326 646398 537562 646634
rect 537646 646398 537882 646634
rect 537326 610718 537562 610954
rect 537646 610718 537882 610954
rect 537326 610398 537562 610634
rect 537646 610398 537882 610634
rect 537326 574718 537562 574954
rect 537646 574718 537882 574954
rect 537326 574398 537562 574634
rect 537646 574398 537882 574634
rect 537326 538718 537562 538954
rect 537646 538718 537882 538954
rect 537326 538398 537562 538634
rect 537646 538398 537882 538634
rect 537326 502718 537562 502954
rect 537646 502718 537882 502954
rect 537326 502398 537562 502634
rect 537646 502398 537882 502634
rect 537326 466718 537562 466954
rect 537646 466718 537882 466954
rect 537326 466398 537562 466634
rect 537646 466398 537882 466634
rect 537326 430718 537562 430954
rect 537646 430718 537882 430954
rect 537326 430398 537562 430634
rect 537646 430398 537882 430634
rect 537326 394718 537562 394954
rect 537646 394718 537882 394954
rect 537326 394398 537562 394634
rect 537646 394398 537882 394634
rect 537326 358718 537562 358954
rect 537646 358718 537882 358954
rect 537326 358398 537562 358634
rect 537646 358398 537882 358634
rect 537326 322718 537562 322954
rect 537646 322718 537882 322954
rect 537326 322398 537562 322634
rect 537646 322398 537882 322634
rect 537326 286718 537562 286954
rect 537646 286718 537882 286954
rect 537326 286398 537562 286634
rect 537646 286398 537882 286634
rect 537326 250718 537562 250954
rect 537646 250718 537882 250954
rect 537326 250398 537562 250634
rect 537646 250398 537882 250634
rect 537326 214718 537562 214954
rect 537646 214718 537882 214954
rect 537326 214398 537562 214634
rect 537646 214398 537882 214634
rect 537326 178718 537562 178954
rect 537646 178718 537882 178954
rect 537326 178398 537562 178634
rect 537646 178398 537882 178634
rect 537326 142718 537562 142954
rect 537646 142718 537882 142954
rect 537326 142398 537562 142634
rect 537646 142398 537882 142634
rect 537326 106718 537562 106954
rect 537646 106718 537882 106954
rect 537326 106398 537562 106634
rect 537646 106398 537882 106634
rect 537326 70718 537562 70954
rect 537646 70718 537882 70954
rect 537326 70398 537562 70634
rect 537646 70398 537882 70634
rect 537326 34718 537562 34954
rect 537646 34718 537882 34954
rect 537326 34398 537562 34634
rect 537646 34398 537882 34634
rect 537326 -7302 537562 -7066
rect 537646 -7302 537882 -7066
rect 537326 -7622 537562 -7386
rect 537646 -7622 537882 -7386
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 546326 705562 546562 705798
rect 546646 705562 546882 705798
rect 546326 705242 546562 705478
rect 546646 705242 546882 705478
rect 546326 691718 546562 691954
rect 546646 691718 546882 691954
rect 546326 691398 546562 691634
rect 546646 691398 546882 691634
rect 546326 655718 546562 655954
rect 546646 655718 546882 655954
rect 546326 655398 546562 655634
rect 546646 655398 546882 655634
rect 546326 619718 546562 619954
rect 546646 619718 546882 619954
rect 546326 619398 546562 619634
rect 546646 619398 546882 619634
rect 546326 583718 546562 583954
rect 546646 583718 546882 583954
rect 546326 583398 546562 583634
rect 546646 583398 546882 583634
rect 546326 547718 546562 547954
rect 546646 547718 546882 547954
rect 546326 547398 546562 547634
rect 546646 547398 546882 547634
rect 546326 511718 546562 511954
rect 546646 511718 546882 511954
rect 546326 511398 546562 511634
rect 546646 511398 546882 511634
rect 546326 475718 546562 475954
rect 546646 475718 546882 475954
rect 546326 475398 546562 475634
rect 546646 475398 546882 475634
rect 546326 439718 546562 439954
rect 546646 439718 546882 439954
rect 546326 439398 546562 439634
rect 546646 439398 546882 439634
rect 546326 403718 546562 403954
rect 546646 403718 546882 403954
rect 546326 403398 546562 403634
rect 546646 403398 546882 403634
rect 546326 367718 546562 367954
rect 546646 367718 546882 367954
rect 546326 367398 546562 367634
rect 546646 367398 546882 367634
rect 546326 331718 546562 331954
rect 546646 331718 546882 331954
rect 546326 331398 546562 331634
rect 546646 331398 546882 331634
rect 546326 295718 546562 295954
rect 546646 295718 546882 295954
rect 546326 295398 546562 295634
rect 546646 295398 546882 295634
rect 546326 259718 546562 259954
rect 546646 259718 546882 259954
rect 546326 259398 546562 259634
rect 546646 259398 546882 259634
rect 546326 223718 546562 223954
rect 546646 223718 546882 223954
rect 546326 223398 546562 223634
rect 546646 223398 546882 223634
rect 546326 187718 546562 187954
rect 546646 187718 546882 187954
rect 546326 187398 546562 187634
rect 546646 187398 546882 187634
rect 546326 151718 546562 151954
rect 546646 151718 546882 151954
rect 546326 151398 546562 151634
rect 546646 151398 546882 151634
rect 546326 115718 546562 115954
rect 546646 115718 546882 115954
rect 546326 115398 546562 115634
rect 546646 115398 546882 115634
rect 546326 79718 546562 79954
rect 546646 79718 546882 79954
rect 546326 79398 546562 79634
rect 546646 79398 546882 79634
rect 546326 43718 546562 43954
rect 546646 43718 546882 43954
rect 546326 43398 546562 43634
rect 546646 43398 546882 43634
rect 546326 7718 546562 7954
rect 546646 7718 546882 7954
rect 546326 7398 546562 7634
rect 546646 7398 546882 7634
rect 546326 -1542 546562 -1306
rect 546646 -1542 546882 -1306
rect 546326 -1862 546562 -1626
rect 546646 -1862 546882 -1626
rect 550826 706522 551062 706758
rect 551146 706522 551382 706758
rect 550826 706202 551062 706438
rect 551146 706202 551382 706438
rect 550826 696218 551062 696454
rect 551146 696218 551382 696454
rect 550826 695898 551062 696134
rect 551146 695898 551382 696134
rect 550826 660218 551062 660454
rect 551146 660218 551382 660454
rect 550826 659898 551062 660134
rect 551146 659898 551382 660134
rect 550826 624218 551062 624454
rect 551146 624218 551382 624454
rect 550826 623898 551062 624134
rect 551146 623898 551382 624134
rect 550826 588218 551062 588454
rect 551146 588218 551382 588454
rect 550826 587898 551062 588134
rect 551146 587898 551382 588134
rect 550826 552218 551062 552454
rect 551146 552218 551382 552454
rect 550826 551898 551062 552134
rect 551146 551898 551382 552134
rect 550826 516218 551062 516454
rect 551146 516218 551382 516454
rect 550826 515898 551062 516134
rect 551146 515898 551382 516134
rect 550826 480218 551062 480454
rect 551146 480218 551382 480454
rect 550826 479898 551062 480134
rect 551146 479898 551382 480134
rect 550826 444218 551062 444454
rect 551146 444218 551382 444454
rect 550826 443898 551062 444134
rect 551146 443898 551382 444134
rect 550826 408218 551062 408454
rect 551146 408218 551382 408454
rect 550826 407898 551062 408134
rect 551146 407898 551382 408134
rect 550826 372218 551062 372454
rect 551146 372218 551382 372454
rect 550826 371898 551062 372134
rect 551146 371898 551382 372134
rect 550826 336218 551062 336454
rect 551146 336218 551382 336454
rect 550826 335898 551062 336134
rect 551146 335898 551382 336134
rect 550826 300218 551062 300454
rect 551146 300218 551382 300454
rect 550826 299898 551062 300134
rect 551146 299898 551382 300134
rect 550826 264218 551062 264454
rect 551146 264218 551382 264454
rect 550826 263898 551062 264134
rect 551146 263898 551382 264134
rect 550826 228218 551062 228454
rect 551146 228218 551382 228454
rect 550826 227898 551062 228134
rect 551146 227898 551382 228134
rect 550826 192218 551062 192454
rect 551146 192218 551382 192454
rect 550826 191898 551062 192134
rect 551146 191898 551382 192134
rect 550826 156218 551062 156454
rect 551146 156218 551382 156454
rect 550826 155898 551062 156134
rect 551146 155898 551382 156134
rect 550826 120218 551062 120454
rect 551146 120218 551382 120454
rect 550826 119898 551062 120134
rect 551146 119898 551382 120134
rect 550826 84218 551062 84454
rect 551146 84218 551382 84454
rect 550826 83898 551062 84134
rect 551146 83898 551382 84134
rect 550826 48218 551062 48454
rect 551146 48218 551382 48454
rect 550826 47898 551062 48134
rect 551146 47898 551382 48134
rect 550826 12218 551062 12454
rect 551146 12218 551382 12454
rect 550826 11898 551062 12134
rect 551146 11898 551382 12134
rect 550826 -2502 551062 -2266
rect 551146 -2502 551382 -2266
rect 550826 -2822 551062 -2586
rect 551146 -2822 551382 -2586
rect 555326 707482 555562 707718
rect 555646 707482 555882 707718
rect 555326 707162 555562 707398
rect 555646 707162 555882 707398
rect 555326 700718 555562 700954
rect 555646 700718 555882 700954
rect 555326 700398 555562 700634
rect 555646 700398 555882 700634
rect 555326 664718 555562 664954
rect 555646 664718 555882 664954
rect 555326 664398 555562 664634
rect 555646 664398 555882 664634
rect 555326 628718 555562 628954
rect 555646 628718 555882 628954
rect 555326 628398 555562 628634
rect 555646 628398 555882 628634
rect 555326 592718 555562 592954
rect 555646 592718 555882 592954
rect 555326 592398 555562 592634
rect 555646 592398 555882 592634
rect 555326 556718 555562 556954
rect 555646 556718 555882 556954
rect 555326 556398 555562 556634
rect 555646 556398 555882 556634
rect 555326 520718 555562 520954
rect 555646 520718 555882 520954
rect 555326 520398 555562 520634
rect 555646 520398 555882 520634
rect 555326 484718 555562 484954
rect 555646 484718 555882 484954
rect 555326 484398 555562 484634
rect 555646 484398 555882 484634
rect 555326 448718 555562 448954
rect 555646 448718 555882 448954
rect 555326 448398 555562 448634
rect 555646 448398 555882 448634
rect 555326 412718 555562 412954
rect 555646 412718 555882 412954
rect 555326 412398 555562 412634
rect 555646 412398 555882 412634
rect 555326 376718 555562 376954
rect 555646 376718 555882 376954
rect 555326 376398 555562 376634
rect 555646 376398 555882 376634
rect 555326 340718 555562 340954
rect 555646 340718 555882 340954
rect 555326 340398 555562 340634
rect 555646 340398 555882 340634
rect 555326 304718 555562 304954
rect 555646 304718 555882 304954
rect 555326 304398 555562 304634
rect 555646 304398 555882 304634
rect 555326 268718 555562 268954
rect 555646 268718 555882 268954
rect 555326 268398 555562 268634
rect 555646 268398 555882 268634
rect 555326 232718 555562 232954
rect 555646 232718 555882 232954
rect 555326 232398 555562 232634
rect 555646 232398 555882 232634
rect 555326 196718 555562 196954
rect 555646 196718 555882 196954
rect 555326 196398 555562 196634
rect 555646 196398 555882 196634
rect 555326 160718 555562 160954
rect 555646 160718 555882 160954
rect 555326 160398 555562 160634
rect 555646 160398 555882 160634
rect 555326 124718 555562 124954
rect 555646 124718 555882 124954
rect 555326 124398 555562 124634
rect 555646 124398 555882 124634
rect 555326 88718 555562 88954
rect 555646 88718 555882 88954
rect 555326 88398 555562 88634
rect 555646 88398 555882 88634
rect 555326 52718 555562 52954
rect 555646 52718 555882 52954
rect 555326 52398 555562 52634
rect 555646 52398 555882 52634
rect 555326 16718 555562 16954
rect 555646 16718 555882 16954
rect 555326 16398 555562 16634
rect 555646 16398 555882 16634
rect 555326 -3462 555562 -3226
rect 555646 -3462 555882 -3226
rect 555326 -3782 555562 -3546
rect 555646 -3782 555882 -3546
rect 559826 708442 560062 708678
rect 560146 708442 560382 708678
rect 559826 708122 560062 708358
rect 560146 708122 560382 708358
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -4422 560062 -4186
rect 560146 -4422 560382 -4186
rect 559826 -4742 560062 -4506
rect 560146 -4742 560382 -4506
rect 564326 709402 564562 709638
rect 564646 709402 564882 709638
rect 564326 709082 564562 709318
rect 564646 709082 564882 709318
rect 564326 673718 564562 673954
rect 564646 673718 564882 673954
rect 564326 673398 564562 673634
rect 564646 673398 564882 673634
rect 564326 637718 564562 637954
rect 564646 637718 564882 637954
rect 564326 637398 564562 637634
rect 564646 637398 564882 637634
rect 564326 601718 564562 601954
rect 564646 601718 564882 601954
rect 564326 601398 564562 601634
rect 564646 601398 564882 601634
rect 564326 565718 564562 565954
rect 564646 565718 564882 565954
rect 564326 565398 564562 565634
rect 564646 565398 564882 565634
rect 564326 529718 564562 529954
rect 564646 529718 564882 529954
rect 564326 529398 564562 529634
rect 564646 529398 564882 529634
rect 564326 493718 564562 493954
rect 564646 493718 564882 493954
rect 564326 493398 564562 493634
rect 564646 493398 564882 493634
rect 564326 457718 564562 457954
rect 564646 457718 564882 457954
rect 564326 457398 564562 457634
rect 564646 457398 564882 457634
rect 564326 421718 564562 421954
rect 564646 421718 564882 421954
rect 564326 421398 564562 421634
rect 564646 421398 564882 421634
rect 564326 385718 564562 385954
rect 564646 385718 564882 385954
rect 564326 385398 564562 385634
rect 564646 385398 564882 385634
rect 564326 349718 564562 349954
rect 564646 349718 564882 349954
rect 564326 349398 564562 349634
rect 564646 349398 564882 349634
rect 564326 313718 564562 313954
rect 564646 313718 564882 313954
rect 564326 313398 564562 313634
rect 564646 313398 564882 313634
rect 564326 277718 564562 277954
rect 564646 277718 564882 277954
rect 564326 277398 564562 277634
rect 564646 277398 564882 277634
rect 564326 241718 564562 241954
rect 564646 241718 564882 241954
rect 564326 241398 564562 241634
rect 564646 241398 564882 241634
rect 564326 205718 564562 205954
rect 564646 205718 564882 205954
rect 564326 205398 564562 205634
rect 564646 205398 564882 205634
rect 564326 169718 564562 169954
rect 564646 169718 564882 169954
rect 564326 169398 564562 169634
rect 564646 169398 564882 169634
rect 564326 133718 564562 133954
rect 564646 133718 564882 133954
rect 564326 133398 564562 133634
rect 564646 133398 564882 133634
rect 564326 97718 564562 97954
rect 564646 97718 564882 97954
rect 564326 97398 564562 97634
rect 564646 97398 564882 97634
rect 564326 61718 564562 61954
rect 564646 61718 564882 61954
rect 564326 61398 564562 61634
rect 564646 61398 564882 61634
rect 564326 25718 564562 25954
rect 564646 25718 564882 25954
rect 564326 25398 564562 25634
rect 564646 25398 564882 25634
rect 564326 -5382 564562 -5146
rect 564646 -5382 564882 -5146
rect 564326 -5702 564562 -5466
rect 564646 -5702 564882 -5466
rect 568826 710362 569062 710598
rect 569146 710362 569382 710598
rect 568826 710042 569062 710278
rect 569146 710042 569382 710278
rect 568826 678218 569062 678454
rect 569146 678218 569382 678454
rect 568826 677898 569062 678134
rect 569146 677898 569382 678134
rect 568826 642218 569062 642454
rect 569146 642218 569382 642454
rect 568826 641898 569062 642134
rect 569146 641898 569382 642134
rect 568826 606218 569062 606454
rect 569146 606218 569382 606454
rect 568826 605898 569062 606134
rect 569146 605898 569382 606134
rect 568826 570218 569062 570454
rect 569146 570218 569382 570454
rect 568826 569898 569062 570134
rect 569146 569898 569382 570134
rect 568826 534218 569062 534454
rect 569146 534218 569382 534454
rect 568826 533898 569062 534134
rect 569146 533898 569382 534134
rect 568826 498218 569062 498454
rect 569146 498218 569382 498454
rect 568826 497898 569062 498134
rect 569146 497898 569382 498134
rect 568826 462218 569062 462454
rect 569146 462218 569382 462454
rect 568826 461898 569062 462134
rect 569146 461898 569382 462134
rect 568826 426218 569062 426454
rect 569146 426218 569382 426454
rect 568826 425898 569062 426134
rect 569146 425898 569382 426134
rect 568826 390218 569062 390454
rect 569146 390218 569382 390454
rect 568826 389898 569062 390134
rect 569146 389898 569382 390134
rect 568826 354218 569062 354454
rect 569146 354218 569382 354454
rect 568826 353898 569062 354134
rect 569146 353898 569382 354134
rect 568826 318218 569062 318454
rect 569146 318218 569382 318454
rect 568826 317898 569062 318134
rect 569146 317898 569382 318134
rect 568826 282218 569062 282454
rect 569146 282218 569382 282454
rect 568826 281898 569062 282134
rect 569146 281898 569382 282134
rect 568826 246218 569062 246454
rect 569146 246218 569382 246454
rect 568826 245898 569062 246134
rect 569146 245898 569382 246134
rect 568826 210218 569062 210454
rect 569146 210218 569382 210454
rect 568826 209898 569062 210134
rect 569146 209898 569382 210134
rect 568826 174218 569062 174454
rect 569146 174218 569382 174454
rect 568826 173898 569062 174134
rect 569146 173898 569382 174134
rect 568826 138218 569062 138454
rect 569146 138218 569382 138454
rect 568826 137898 569062 138134
rect 569146 137898 569382 138134
rect 568826 102218 569062 102454
rect 569146 102218 569382 102454
rect 568826 101898 569062 102134
rect 569146 101898 569382 102134
rect 568826 66218 569062 66454
rect 569146 66218 569382 66454
rect 568826 65898 569062 66134
rect 569146 65898 569382 66134
rect 568826 30218 569062 30454
rect 569146 30218 569382 30454
rect 568826 29898 569062 30134
rect 569146 29898 569382 30134
rect 568826 -6342 569062 -6106
rect 569146 -6342 569382 -6106
rect 568826 -6662 569062 -6426
rect 569146 -6662 569382 -6426
rect 573326 711322 573562 711558
rect 573646 711322 573882 711558
rect 573326 711002 573562 711238
rect 573646 711002 573882 711238
rect 573326 682718 573562 682954
rect 573646 682718 573882 682954
rect 573326 682398 573562 682634
rect 573646 682398 573882 682634
rect 573326 646718 573562 646954
rect 573646 646718 573882 646954
rect 573326 646398 573562 646634
rect 573646 646398 573882 646634
rect 573326 610718 573562 610954
rect 573646 610718 573882 610954
rect 573326 610398 573562 610634
rect 573646 610398 573882 610634
rect 573326 574718 573562 574954
rect 573646 574718 573882 574954
rect 573326 574398 573562 574634
rect 573646 574398 573882 574634
rect 573326 538718 573562 538954
rect 573646 538718 573882 538954
rect 573326 538398 573562 538634
rect 573646 538398 573882 538634
rect 573326 502718 573562 502954
rect 573646 502718 573882 502954
rect 573326 502398 573562 502634
rect 573646 502398 573882 502634
rect 573326 466718 573562 466954
rect 573646 466718 573882 466954
rect 573326 466398 573562 466634
rect 573646 466398 573882 466634
rect 573326 430718 573562 430954
rect 573646 430718 573882 430954
rect 573326 430398 573562 430634
rect 573646 430398 573882 430634
rect 573326 394718 573562 394954
rect 573646 394718 573882 394954
rect 573326 394398 573562 394634
rect 573646 394398 573882 394634
rect 573326 358718 573562 358954
rect 573646 358718 573882 358954
rect 573326 358398 573562 358634
rect 573646 358398 573882 358634
rect 573326 322718 573562 322954
rect 573646 322718 573882 322954
rect 573326 322398 573562 322634
rect 573646 322398 573882 322634
rect 573326 286718 573562 286954
rect 573646 286718 573882 286954
rect 573326 286398 573562 286634
rect 573646 286398 573882 286634
rect 573326 250718 573562 250954
rect 573646 250718 573882 250954
rect 573326 250398 573562 250634
rect 573646 250398 573882 250634
rect 573326 214718 573562 214954
rect 573646 214718 573882 214954
rect 573326 214398 573562 214634
rect 573646 214398 573882 214634
rect 573326 178718 573562 178954
rect 573646 178718 573882 178954
rect 573326 178398 573562 178634
rect 573646 178398 573882 178634
rect 573326 142718 573562 142954
rect 573646 142718 573882 142954
rect 573326 142398 573562 142634
rect 573646 142398 573882 142634
rect 573326 106718 573562 106954
rect 573646 106718 573882 106954
rect 573326 106398 573562 106634
rect 573646 106398 573882 106634
rect 573326 70718 573562 70954
rect 573646 70718 573882 70954
rect 573326 70398 573562 70634
rect 573646 70398 573882 70634
rect 573326 34718 573562 34954
rect 573646 34718 573882 34954
rect 573326 34398 573562 34634
rect 573646 34398 573882 34634
rect 573326 -7302 573562 -7066
rect 573646 -7302 573882 -7066
rect 573326 -7622 573562 -7386
rect 573646 -7622 573882 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 691718 582562 691954
rect 582646 691718 582882 691954
rect 582326 691398 582562 691634
rect 582646 691398 582882 691634
rect 582326 655718 582562 655954
rect 582646 655718 582882 655954
rect 582326 655398 582562 655634
rect 582646 655398 582882 655634
rect 582326 619718 582562 619954
rect 582646 619718 582882 619954
rect 582326 619398 582562 619634
rect 582646 619398 582882 619634
rect 582326 583718 582562 583954
rect 582646 583718 582882 583954
rect 582326 583398 582562 583634
rect 582646 583398 582882 583634
rect 582326 547718 582562 547954
rect 582646 547718 582882 547954
rect 582326 547398 582562 547634
rect 582646 547398 582882 547634
rect 582326 511718 582562 511954
rect 582646 511718 582882 511954
rect 582326 511398 582562 511634
rect 582646 511398 582882 511634
rect 582326 475718 582562 475954
rect 582646 475718 582882 475954
rect 582326 475398 582562 475634
rect 582646 475398 582882 475634
rect 582326 439718 582562 439954
rect 582646 439718 582882 439954
rect 582326 439398 582562 439634
rect 582646 439398 582882 439634
rect 582326 403718 582562 403954
rect 582646 403718 582882 403954
rect 582326 403398 582562 403634
rect 582646 403398 582882 403634
rect 582326 367718 582562 367954
rect 582646 367718 582882 367954
rect 582326 367398 582562 367634
rect 582646 367398 582882 367634
rect 582326 331718 582562 331954
rect 582646 331718 582882 331954
rect 582326 331398 582562 331634
rect 582646 331398 582882 331634
rect 582326 295718 582562 295954
rect 582646 295718 582882 295954
rect 582326 295398 582562 295634
rect 582646 295398 582882 295634
rect 582326 259718 582562 259954
rect 582646 259718 582882 259954
rect 582326 259398 582562 259634
rect 582646 259398 582882 259634
rect 582326 223718 582562 223954
rect 582646 223718 582882 223954
rect 582326 223398 582562 223634
rect 582646 223398 582882 223634
rect 582326 187718 582562 187954
rect 582646 187718 582882 187954
rect 582326 187398 582562 187634
rect 582646 187398 582882 187634
rect 582326 151718 582562 151954
rect 582646 151718 582882 151954
rect 582326 151398 582562 151634
rect 582646 151398 582882 151634
rect 582326 115718 582562 115954
rect 582646 115718 582882 115954
rect 582326 115398 582562 115634
rect 582646 115398 582882 115634
rect 582326 79718 582562 79954
rect 582646 79718 582882 79954
rect 582326 79398 582562 79634
rect 582646 79398 582882 79634
rect 582326 43718 582562 43954
rect 582646 43718 582882 43954
rect 582326 43398 582562 43634
rect 582646 43398 582882 43634
rect 582326 7718 582562 7954
rect 582646 7718 582882 7954
rect 582326 7398 582562 7634
rect 582646 7398 582882 7634
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 691718 586538 691954
rect 586622 691718 586858 691954
rect 586302 691398 586538 691634
rect 586622 691398 586858 691634
rect 586302 655718 586538 655954
rect 586622 655718 586858 655954
rect 586302 655398 586538 655634
rect 586622 655398 586858 655634
rect 586302 619718 586538 619954
rect 586622 619718 586858 619954
rect 586302 619398 586538 619634
rect 586622 619398 586858 619634
rect 586302 583718 586538 583954
rect 586622 583718 586858 583954
rect 586302 583398 586538 583634
rect 586622 583398 586858 583634
rect 586302 547718 586538 547954
rect 586622 547718 586858 547954
rect 586302 547398 586538 547634
rect 586622 547398 586858 547634
rect 586302 511718 586538 511954
rect 586622 511718 586858 511954
rect 586302 511398 586538 511634
rect 586622 511398 586858 511634
rect 586302 475718 586538 475954
rect 586622 475718 586858 475954
rect 586302 475398 586538 475634
rect 586622 475398 586858 475634
rect 586302 439718 586538 439954
rect 586622 439718 586858 439954
rect 586302 439398 586538 439634
rect 586622 439398 586858 439634
rect 586302 403718 586538 403954
rect 586622 403718 586858 403954
rect 586302 403398 586538 403634
rect 586622 403398 586858 403634
rect 586302 367718 586538 367954
rect 586622 367718 586858 367954
rect 586302 367398 586538 367634
rect 586622 367398 586858 367634
rect 586302 331718 586538 331954
rect 586622 331718 586858 331954
rect 586302 331398 586538 331634
rect 586622 331398 586858 331634
rect 586302 295718 586538 295954
rect 586622 295718 586858 295954
rect 586302 295398 586538 295634
rect 586622 295398 586858 295634
rect 586302 259718 586538 259954
rect 586622 259718 586858 259954
rect 586302 259398 586538 259634
rect 586622 259398 586858 259634
rect 586302 223718 586538 223954
rect 586622 223718 586858 223954
rect 586302 223398 586538 223634
rect 586622 223398 586858 223634
rect 586302 187718 586538 187954
rect 586622 187718 586858 187954
rect 586302 187398 586538 187634
rect 586622 187398 586858 187634
rect 586302 151718 586538 151954
rect 586622 151718 586858 151954
rect 586302 151398 586538 151634
rect 586622 151398 586858 151634
rect 586302 115718 586538 115954
rect 586622 115718 586858 115954
rect 586302 115398 586538 115634
rect 586622 115398 586858 115634
rect 586302 79718 586538 79954
rect 586622 79718 586858 79954
rect 586302 79398 586538 79634
rect 586622 79398 586858 79634
rect 586302 43718 586538 43954
rect 586622 43718 586858 43954
rect 586302 43398 586538 43634
rect 586622 43398 586858 43634
rect 586302 7718 586538 7954
rect 586622 7718 586858 7954
rect 586302 7398 586538 7634
rect 586622 7398 586858 7634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 696218 587498 696454
rect 587582 696218 587818 696454
rect 587262 695898 587498 696134
rect 587582 695898 587818 696134
rect 587262 660218 587498 660454
rect 587582 660218 587818 660454
rect 587262 659898 587498 660134
rect 587582 659898 587818 660134
rect 587262 624218 587498 624454
rect 587582 624218 587818 624454
rect 587262 623898 587498 624134
rect 587582 623898 587818 624134
rect 587262 588218 587498 588454
rect 587582 588218 587818 588454
rect 587262 587898 587498 588134
rect 587582 587898 587818 588134
rect 587262 552218 587498 552454
rect 587582 552218 587818 552454
rect 587262 551898 587498 552134
rect 587582 551898 587818 552134
rect 587262 516218 587498 516454
rect 587582 516218 587818 516454
rect 587262 515898 587498 516134
rect 587582 515898 587818 516134
rect 587262 480218 587498 480454
rect 587582 480218 587818 480454
rect 587262 479898 587498 480134
rect 587582 479898 587818 480134
rect 587262 444218 587498 444454
rect 587582 444218 587818 444454
rect 587262 443898 587498 444134
rect 587582 443898 587818 444134
rect 587262 408218 587498 408454
rect 587582 408218 587818 408454
rect 587262 407898 587498 408134
rect 587582 407898 587818 408134
rect 587262 372218 587498 372454
rect 587582 372218 587818 372454
rect 587262 371898 587498 372134
rect 587582 371898 587818 372134
rect 587262 336218 587498 336454
rect 587582 336218 587818 336454
rect 587262 335898 587498 336134
rect 587582 335898 587818 336134
rect 587262 300218 587498 300454
rect 587582 300218 587818 300454
rect 587262 299898 587498 300134
rect 587582 299898 587818 300134
rect 587262 264218 587498 264454
rect 587582 264218 587818 264454
rect 587262 263898 587498 264134
rect 587582 263898 587818 264134
rect 587262 228218 587498 228454
rect 587582 228218 587818 228454
rect 587262 227898 587498 228134
rect 587582 227898 587818 228134
rect 587262 192218 587498 192454
rect 587582 192218 587818 192454
rect 587262 191898 587498 192134
rect 587582 191898 587818 192134
rect 587262 156218 587498 156454
rect 587582 156218 587818 156454
rect 587262 155898 587498 156134
rect 587582 155898 587818 156134
rect 587262 120218 587498 120454
rect 587582 120218 587818 120454
rect 587262 119898 587498 120134
rect 587582 119898 587818 120134
rect 587262 84218 587498 84454
rect 587582 84218 587818 84454
rect 587262 83898 587498 84134
rect 587582 83898 587818 84134
rect 587262 48218 587498 48454
rect 587582 48218 587818 48454
rect 587262 47898 587498 48134
rect 587582 47898 587818 48134
rect 587262 12218 587498 12454
rect 587582 12218 587818 12454
rect 587262 11898 587498 12134
rect 587582 11898 587818 12134
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 700718 588458 700954
rect 588542 700718 588778 700954
rect 588222 700398 588458 700634
rect 588542 700398 588778 700634
rect 588222 664718 588458 664954
rect 588542 664718 588778 664954
rect 588222 664398 588458 664634
rect 588542 664398 588778 664634
rect 588222 628718 588458 628954
rect 588542 628718 588778 628954
rect 588222 628398 588458 628634
rect 588542 628398 588778 628634
rect 588222 592718 588458 592954
rect 588542 592718 588778 592954
rect 588222 592398 588458 592634
rect 588542 592398 588778 592634
rect 588222 556718 588458 556954
rect 588542 556718 588778 556954
rect 588222 556398 588458 556634
rect 588542 556398 588778 556634
rect 588222 520718 588458 520954
rect 588542 520718 588778 520954
rect 588222 520398 588458 520634
rect 588542 520398 588778 520634
rect 588222 484718 588458 484954
rect 588542 484718 588778 484954
rect 588222 484398 588458 484634
rect 588542 484398 588778 484634
rect 588222 448718 588458 448954
rect 588542 448718 588778 448954
rect 588222 448398 588458 448634
rect 588542 448398 588778 448634
rect 588222 412718 588458 412954
rect 588542 412718 588778 412954
rect 588222 412398 588458 412634
rect 588542 412398 588778 412634
rect 588222 376718 588458 376954
rect 588542 376718 588778 376954
rect 588222 376398 588458 376634
rect 588542 376398 588778 376634
rect 588222 340718 588458 340954
rect 588542 340718 588778 340954
rect 588222 340398 588458 340634
rect 588542 340398 588778 340634
rect 588222 304718 588458 304954
rect 588542 304718 588778 304954
rect 588222 304398 588458 304634
rect 588542 304398 588778 304634
rect 588222 268718 588458 268954
rect 588542 268718 588778 268954
rect 588222 268398 588458 268634
rect 588542 268398 588778 268634
rect 588222 232718 588458 232954
rect 588542 232718 588778 232954
rect 588222 232398 588458 232634
rect 588542 232398 588778 232634
rect 588222 196718 588458 196954
rect 588542 196718 588778 196954
rect 588222 196398 588458 196634
rect 588542 196398 588778 196634
rect 588222 160718 588458 160954
rect 588542 160718 588778 160954
rect 588222 160398 588458 160634
rect 588542 160398 588778 160634
rect 588222 124718 588458 124954
rect 588542 124718 588778 124954
rect 588222 124398 588458 124634
rect 588542 124398 588778 124634
rect 588222 88718 588458 88954
rect 588542 88718 588778 88954
rect 588222 88398 588458 88634
rect 588542 88398 588778 88634
rect 588222 52718 588458 52954
rect 588542 52718 588778 52954
rect 588222 52398 588458 52634
rect 588542 52398 588778 52634
rect 588222 16718 588458 16954
rect 588542 16718 588778 16954
rect 588222 16398 588458 16634
rect 588542 16398 588778 16634
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 669218 589418 669454
rect 589502 669218 589738 669454
rect 589182 668898 589418 669134
rect 589502 668898 589738 669134
rect 589182 633218 589418 633454
rect 589502 633218 589738 633454
rect 589182 632898 589418 633134
rect 589502 632898 589738 633134
rect 589182 597218 589418 597454
rect 589502 597218 589738 597454
rect 589182 596898 589418 597134
rect 589502 596898 589738 597134
rect 589182 561218 589418 561454
rect 589502 561218 589738 561454
rect 589182 560898 589418 561134
rect 589502 560898 589738 561134
rect 589182 525218 589418 525454
rect 589502 525218 589738 525454
rect 589182 524898 589418 525134
rect 589502 524898 589738 525134
rect 589182 489218 589418 489454
rect 589502 489218 589738 489454
rect 589182 488898 589418 489134
rect 589502 488898 589738 489134
rect 589182 453218 589418 453454
rect 589502 453218 589738 453454
rect 589182 452898 589418 453134
rect 589502 452898 589738 453134
rect 589182 417218 589418 417454
rect 589502 417218 589738 417454
rect 589182 416898 589418 417134
rect 589502 416898 589738 417134
rect 589182 381218 589418 381454
rect 589502 381218 589738 381454
rect 589182 380898 589418 381134
rect 589502 380898 589738 381134
rect 589182 345218 589418 345454
rect 589502 345218 589738 345454
rect 589182 344898 589418 345134
rect 589502 344898 589738 345134
rect 589182 309218 589418 309454
rect 589502 309218 589738 309454
rect 589182 308898 589418 309134
rect 589502 308898 589738 309134
rect 589182 273218 589418 273454
rect 589502 273218 589738 273454
rect 589182 272898 589418 273134
rect 589502 272898 589738 273134
rect 589182 237218 589418 237454
rect 589502 237218 589738 237454
rect 589182 236898 589418 237134
rect 589502 236898 589738 237134
rect 589182 201218 589418 201454
rect 589502 201218 589738 201454
rect 589182 200898 589418 201134
rect 589502 200898 589738 201134
rect 589182 165218 589418 165454
rect 589502 165218 589738 165454
rect 589182 164898 589418 165134
rect 589502 164898 589738 165134
rect 589182 129218 589418 129454
rect 589502 129218 589738 129454
rect 589182 128898 589418 129134
rect 589502 128898 589738 129134
rect 589182 93218 589418 93454
rect 589502 93218 589738 93454
rect 589182 92898 589418 93134
rect 589502 92898 589738 93134
rect 589182 57218 589418 57454
rect 589502 57218 589738 57454
rect 589182 56898 589418 57134
rect 589502 56898 589738 57134
rect 589182 21218 589418 21454
rect 589502 21218 589738 21454
rect 589182 20898 589418 21134
rect 589502 20898 589738 21134
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 673718 590378 673954
rect 590462 673718 590698 673954
rect 590142 673398 590378 673634
rect 590462 673398 590698 673634
rect 590142 637718 590378 637954
rect 590462 637718 590698 637954
rect 590142 637398 590378 637634
rect 590462 637398 590698 637634
rect 590142 601718 590378 601954
rect 590462 601718 590698 601954
rect 590142 601398 590378 601634
rect 590462 601398 590698 601634
rect 590142 565718 590378 565954
rect 590462 565718 590698 565954
rect 590142 565398 590378 565634
rect 590462 565398 590698 565634
rect 590142 529718 590378 529954
rect 590462 529718 590698 529954
rect 590142 529398 590378 529634
rect 590462 529398 590698 529634
rect 590142 493718 590378 493954
rect 590462 493718 590698 493954
rect 590142 493398 590378 493634
rect 590462 493398 590698 493634
rect 590142 457718 590378 457954
rect 590462 457718 590698 457954
rect 590142 457398 590378 457634
rect 590462 457398 590698 457634
rect 590142 421718 590378 421954
rect 590462 421718 590698 421954
rect 590142 421398 590378 421634
rect 590462 421398 590698 421634
rect 590142 385718 590378 385954
rect 590462 385718 590698 385954
rect 590142 385398 590378 385634
rect 590462 385398 590698 385634
rect 590142 349718 590378 349954
rect 590462 349718 590698 349954
rect 590142 349398 590378 349634
rect 590462 349398 590698 349634
rect 590142 313718 590378 313954
rect 590462 313718 590698 313954
rect 590142 313398 590378 313634
rect 590462 313398 590698 313634
rect 590142 277718 590378 277954
rect 590462 277718 590698 277954
rect 590142 277398 590378 277634
rect 590462 277398 590698 277634
rect 590142 241718 590378 241954
rect 590462 241718 590698 241954
rect 590142 241398 590378 241634
rect 590462 241398 590698 241634
rect 590142 205718 590378 205954
rect 590462 205718 590698 205954
rect 590142 205398 590378 205634
rect 590462 205398 590698 205634
rect 590142 169718 590378 169954
rect 590462 169718 590698 169954
rect 590142 169398 590378 169634
rect 590462 169398 590698 169634
rect 590142 133718 590378 133954
rect 590462 133718 590698 133954
rect 590142 133398 590378 133634
rect 590462 133398 590698 133634
rect 590142 97718 590378 97954
rect 590462 97718 590698 97954
rect 590142 97398 590378 97634
rect 590462 97398 590698 97634
rect 590142 61718 590378 61954
rect 590462 61718 590698 61954
rect 590142 61398 590378 61634
rect 590462 61398 590698 61634
rect 590142 25718 590378 25954
rect 590462 25718 590698 25954
rect 590142 25398 590378 25634
rect 590462 25398 590698 25634
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 678218 591338 678454
rect 591422 678218 591658 678454
rect 591102 677898 591338 678134
rect 591422 677898 591658 678134
rect 591102 642218 591338 642454
rect 591422 642218 591658 642454
rect 591102 641898 591338 642134
rect 591422 641898 591658 642134
rect 591102 606218 591338 606454
rect 591422 606218 591658 606454
rect 591102 605898 591338 606134
rect 591422 605898 591658 606134
rect 591102 570218 591338 570454
rect 591422 570218 591658 570454
rect 591102 569898 591338 570134
rect 591422 569898 591658 570134
rect 591102 534218 591338 534454
rect 591422 534218 591658 534454
rect 591102 533898 591338 534134
rect 591422 533898 591658 534134
rect 591102 498218 591338 498454
rect 591422 498218 591658 498454
rect 591102 497898 591338 498134
rect 591422 497898 591658 498134
rect 591102 462218 591338 462454
rect 591422 462218 591658 462454
rect 591102 461898 591338 462134
rect 591422 461898 591658 462134
rect 591102 426218 591338 426454
rect 591422 426218 591658 426454
rect 591102 425898 591338 426134
rect 591422 425898 591658 426134
rect 591102 390218 591338 390454
rect 591422 390218 591658 390454
rect 591102 389898 591338 390134
rect 591422 389898 591658 390134
rect 591102 354218 591338 354454
rect 591422 354218 591658 354454
rect 591102 353898 591338 354134
rect 591422 353898 591658 354134
rect 591102 318218 591338 318454
rect 591422 318218 591658 318454
rect 591102 317898 591338 318134
rect 591422 317898 591658 318134
rect 591102 282218 591338 282454
rect 591422 282218 591658 282454
rect 591102 281898 591338 282134
rect 591422 281898 591658 282134
rect 591102 246218 591338 246454
rect 591422 246218 591658 246454
rect 591102 245898 591338 246134
rect 591422 245898 591658 246134
rect 591102 210218 591338 210454
rect 591422 210218 591658 210454
rect 591102 209898 591338 210134
rect 591422 209898 591658 210134
rect 591102 174218 591338 174454
rect 591422 174218 591658 174454
rect 591102 173898 591338 174134
rect 591422 173898 591658 174134
rect 591102 138218 591338 138454
rect 591422 138218 591658 138454
rect 591102 137898 591338 138134
rect 591422 137898 591658 138134
rect 591102 102218 591338 102454
rect 591422 102218 591658 102454
rect 591102 101898 591338 102134
rect 591422 101898 591658 102134
rect 591102 66218 591338 66454
rect 591422 66218 591658 66454
rect 591102 65898 591338 66134
rect 591422 65898 591658 66134
rect 591102 30218 591338 30454
rect 591422 30218 591658 30454
rect 591102 29898 591338 30134
rect 591422 29898 591658 30134
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 682718 592298 682954
rect 592382 682718 592618 682954
rect 592062 682398 592298 682634
rect 592382 682398 592618 682634
rect 592062 646718 592298 646954
rect 592382 646718 592618 646954
rect 592062 646398 592298 646634
rect 592382 646398 592618 646634
rect 592062 610718 592298 610954
rect 592382 610718 592618 610954
rect 592062 610398 592298 610634
rect 592382 610398 592618 610634
rect 592062 574718 592298 574954
rect 592382 574718 592618 574954
rect 592062 574398 592298 574634
rect 592382 574398 592618 574634
rect 592062 538718 592298 538954
rect 592382 538718 592618 538954
rect 592062 538398 592298 538634
rect 592382 538398 592618 538634
rect 592062 502718 592298 502954
rect 592382 502718 592618 502954
rect 592062 502398 592298 502634
rect 592382 502398 592618 502634
rect 592062 466718 592298 466954
rect 592382 466718 592618 466954
rect 592062 466398 592298 466634
rect 592382 466398 592618 466634
rect 592062 430718 592298 430954
rect 592382 430718 592618 430954
rect 592062 430398 592298 430634
rect 592382 430398 592618 430634
rect 592062 394718 592298 394954
rect 592382 394718 592618 394954
rect 592062 394398 592298 394634
rect 592382 394398 592618 394634
rect 592062 358718 592298 358954
rect 592382 358718 592618 358954
rect 592062 358398 592298 358634
rect 592382 358398 592618 358634
rect 592062 322718 592298 322954
rect 592382 322718 592618 322954
rect 592062 322398 592298 322634
rect 592382 322398 592618 322634
rect 592062 286718 592298 286954
rect 592382 286718 592618 286954
rect 592062 286398 592298 286634
rect 592382 286398 592618 286634
rect 592062 250718 592298 250954
rect 592382 250718 592618 250954
rect 592062 250398 592298 250634
rect 592382 250398 592618 250634
rect 592062 214718 592298 214954
rect 592382 214718 592618 214954
rect 592062 214398 592298 214634
rect 592382 214398 592618 214634
rect 592062 178718 592298 178954
rect 592382 178718 592618 178954
rect 592062 178398 592298 178634
rect 592382 178398 592618 178634
rect 592062 142718 592298 142954
rect 592382 142718 592618 142954
rect 592062 142398 592298 142634
rect 592382 142398 592618 142634
rect 592062 106718 592298 106954
rect 592382 106718 592618 106954
rect 592062 106398 592298 106634
rect 592382 106398 592618 106634
rect 592062 70718 592298 70954
rect 592382 70718 592618 70954
rect 592062 70398 592298 70634
rect 592382 70398 592618 70634
rect 592062 34718 592298 34954
rect 592382 34718 592618 34954
rect 592062 34398 592298 34634
rect 592382 34398 592618 34634
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 33326 711558
rect 33562 711322 33646 711558
rect 33882 711322 69326 711558
rect 69562 711322 69646 711558
rect 69882 711322 105326 711558
rect 105562 711322 105646 711558
rect 105882 711322 141326 711558
rect 141562 711322 141646 711558
rect 141882 711322 177326 711558
rect 177562 711322 177646 711558
rect 177882 711322 213326 711558
rect 213562 711322 213646 711558
rect 213882 711322 249326 711558
rect 249562 711322 249646 711558
rect 249882 711322 285326 711558
rect 285562 711322 285646 711558
rect 285882 711322 321326 711558
rect 321562 711322 321646 711558
rect 321882 711322 357326 711558
rect 357562 711322 357646 711558
rect 357882 711322 393326 711558
rect 393562 711322 393646 711558
rect 393882 711322 429326 711558
rect 429562 711322 429646 711558
rect 429882 711322 465326 711558
rect 465562 711322 465646 711558
rect 465882 711322 501326 711558
rect 501562 711322 501646 711558
rect 501882 711322 537326 711558
rect 537562 711322 537646 711558
rect 537882 711322 573326 711558
rect 573562 711322 573646 711558
rect 573882 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 33326 711238
rect 33562 711002 33646 711238
rect 33882 711002 69326 711238
rect 69562 711002 69646 711238
rect 69882 711002 105326 711238
rect 105562 711002 105646 711238
rect 105882 711002 141326 711238
rect 141562 711002 141646 711238
rect 141882 711002 177326 711238
rect 177562 711002 177646 711238
rect 177882 711002 213326 711238
rect 213562 711002 213646 711238
rect 213882 711002 249326 711238
rect 249562 711002 249646 711238
rect 249882 711002 285326 711238
rect 285562 711002 285646 711238
rect 285882 711002 321326 711238
rect 321562 711002 321646 711238
rect 321882 711002 357326 711238
rect 357562 711002 357646 711238
rect 357882 711002 393326 711238
rect 393562 711002 393646 711238
rect 393882 711002 429326 711238
rect 429562 711002 429646 711238
rect 429882 711002 465326 711238
rect 465562 711002 465646 711238
rect 465882 711002 501326 711238
rect 501562 711002 501646 711238
rect 501882 711002 537326 711238
rect 537562 711002 537646 711238
rect 537882 711002 573326 711238
rect 573562 711002 573646 711238
rect 573882 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 28826 710598
rect 29062 710362 29146 710598
rect 29382 710362 64826 710598
rect 65062 710362 65146 710598
rect 65382 710362 100826 710598
rect 101062 710362 101146 710598
rect 101382 710362 136826 710598
rect 137062 710362 137146 710598
rect 137382 710362 172826 710598
rect 173062 710362 173146 710598
rect 173382 710362 208826 710598
rect 209062 710362 209146 710598
rect 209382 710362 244826 710598
rect 245062 710362 245146 710598
rect 245382 710362 280826 710598
rect 281062 710362 281146 710598
rect 281382 710362 316826 710598
rect 317062 710362 317146 710598
rect 317382 710362 352826 710598
rect 353062 710362 353146 710598
rect 353382 710362 388826 710598
rect 389062 710362 389146 710598
rect 389382 710362 424826 710598
rect 425062 710362 425146 710598
rect 425382 710362 460826 710598
rect 461062 710362 461146 710598
rect 461382 710362 496826 710598
rect 497062 710362 497146 710598
rect 497382 710362 532826 710598
rect 533062 710362 533146 710598
rect 533382 710362 568826 710598
rect 569062 710362 569146 710598
rect 569382 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 28826 710278
rect 29062 710042 29146 710278
rect 29382 710042 64826 710278
rect 65062 710042 65146 710278
rect 65382 710042 100826 710278
rect 101062 710042 101146 710278
rect 101382 710042 136826 710278
rect 137062 710042 137146 710278
rect 137382 710042 172826 710278
rect 173062 710042 173146 710278
rect 173382 710042 208826 710278
rect 209062 710042 209146 710278
rect 209382 710042 244826 710278
rect 245062 710042 245146 710278
rect 245382 710042 280826 710278
rect 281062 710042 281146 710278
rect 281382 710042 316826 710278
rect 317062 710042 317146 710278
rect 317382 710042 352826 710278
rect 353062 710042 353146 710278
rect 353382 710042 388826 710278
rect 389062 710042 389146 710278
rect 389382 710042 424826 710278
rect 425062 710042 425146 710278
rect 425382 710042 460826 710278
rect 461062 710042 461146 710278
rect 461382 710042 496826 710278
rect 497062 710042 497146 710278
rect 497382 710042 532826 710278
rect 533062 710042 533146 710278
rect 533382 710042 568826 710278
rect 569062 710042 569146 710278
rect 569382 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 24326 709638
rect 24562 709402 24646 709638
rect 24882 709402 60326 709638
rect 60562 709402 60646 709638
rect 60882 709402 96326 709638
rect 96562 709402 96646 709638
rect 96882 709402 132326 709638
rect 132562 709402 132646 709638
rect 132882 709402 168326 709638
rect 168562 709402 168646 709638
rect 168882 709402 204326 709638
rect 204562 709402 204646 709638
rect 204882 709402 240326 709638
rect 240562 709402 240646 709638
rect 240882 709402 276326 709638
rect 276562 709402 276646 709638
rect 276882 709402 312326 709638
rect 312562 709402 312646 709638
rect 312882 709402 348326 709638
rect 348562 709402 348646 709638
rect 348882 709402 384326 709638
rect 384562 709402 384646 709638
rect 384882 709402 420326 709638
rect 420562 709402 420646 709638
rect 420882 709402 456326 709638
rect 456562 709402 456646 709638
rect 456882 709402 492326 709638
rect 492562 709402 492646 709638
rect 492882 709402 528326 709638
rect 528562 709402 528646 709638
rect 528882 709402 564326 709638
rect 564562 709402 564646 709638
rect 564882 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 24326 709318
rect 24562 709082 24646 709318
rect 24882 709082 60326 709318
rect 60562 709082 60646 709318
rect 60882 709082 96326 709318
rect 96562 709082 96646 709318
rect 96882 709082 132326 709318
rect 132562 709082 132646 709318
rect 132882 709082 168326 709318
rect 168562 709082 168646 709318
rect 168882 709082 204326 709318
rect 204562 709082 204646 709318
rect 204882 709082 240326 709318
rect 240562 709082 240646 709318
rect 240882 709082 276326 709318
rect 276562 709082 276646 709318
rect 276882 709082 312326 709318
rect 312562 709082 312646 709318
rect 312882 709082 348326 709318
rect 348562 709082 348646 709318
rect 348882 709082 384326 709318
rect 384562 709082 384646 709318
rect 384882 709082 420326 709318
rect 420562 709082 420646 709318
rect 420882 709082 456326 709318
rect 456562 709082 456646 709318
rect 456882 709082 492326 709318
rect 492562 709082 492646 709318
rect 492882 709082 528326 709318
rect 528562 709082 528646 709318
rect 528882 709082 564326 709318
rect 564562 709082 564646 709318
rect 564882 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 19826 708678
rect 20062 708442 20146 708678
rect 20382 708442 55826 708678
rect 56062 708442 56146 708678
rect 56382 708442 91826 708678
rect 92062 708442 92146 708678
rect 92382 708442 127826 708678
rect 128062 708442 128146 708678
rect 128382 708442 163826 708678
rect 164062 708442 164146 708678
rect 164382 708442 199826 708678
rect 200062 708442 200146 708678
rect 200382 708442 235826 708678
rect 236062 708442 236146 708678
rect 236382 708442 271826 708678
rect 272062 708442 272146 708678
rect 272382 708442 307826 708678
rect 308062 708442 308146 708678
rect 308382 708442 343826 708678
rect 344062 708442 344146 708678
rect 344382 708442 379826 708678
rect 380062 708442 380146 708678
rect 380382 708442 415826 708678
rect 416062 708442 416146 708678
rect 416382 708442 451826 708678
rect 452062 708442 452146 708678
rect 452382 708442 487826 708678
rect 488062 708442 488146 708678
rect 488382 708442 523826 708678
rect 524062 708442 524146 708678
rect 524382 708442 559826 708678
rect 560062 708442 560146 708678
rect 560382 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 19826 708358
rect 20062 708122 20146 708358
rect 20382 708122 55826 708358
rect 56062 708122 56146 708358
rect 56382 708122 91826 708358
rect 92062 708122 92146 708358
rect 92382 708122 127826 708358
rect 128062 708122 128146 708358
rect 128382 708122 163826 708358
rect 164062 708122 164146 708358
rect 164382 708122 199826 708358
rect 200062 708122 200146 708358
rect 200382 708122 235826 708358
rect 236062 708122 236146 708358
rect 236382 708122 271826 708358
rect 272062 708122 272146 708358
rect 272382 708122 307826 708358
rect 308062 708122 308146 708358
rect 308382 708122 343826 708358
rect 344062 708122 344146 708358
rect 344382 708122 379826 708358
rect 380062 708122 380146 708358
rect 380382 708122 415826 708358
rect 416062 708122 416146 708358
rect 416382 708122 451826 708358
rect 452062 708122 452146 708358
rect 452382 708122 487826 708358
rect 488062 708122 488146 708358
rect 488382 708122 523826 708358
rect 524062 708122 524146 708358
rect 524382 708122 559826 708358
rect 560062 708122 560146 708358
rect 560382 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 15326 707718
rect 15562 707482 15646 707718
rect 15882 707482 51326 707718
rect 51562 707482 51646 707718
rect 51882 707482 87326 707718
rect 87562 707482 87646 707718
rect 87882 707482 123326 707718
rect 123562 707482 123646 707718
rect 123882 707482 159326 707718
rect 159562 707482 159646 707718
rect 159882 707482 195326 707718
rect 195562 707482 195646 707718
rect 195882 707482 231326 707718
rect 231562 707482 231646 707718
rect 231882 707482 267326 707718
rect 267562 707482 267646 707718
rect 267882 707482 303326 707718
rect 303562 707482 303646 707718
rect 303882 707482 339326 707718
rect 339562 707482 339646 707718
rect 339882 707482 375326 707718
rect 375562 707482 375646 707718
rect 375882 707482 411326 707718
rect 411562 707482 411646 707718
rect 411882 707482 447326 707718
rect 447562 707482 447646 707718
rect 447882 707482 483326 707718
rect 483562 707482 483646 707718
rect 483882 707482 519326 707718
rect 519562 707482 519646 707718
rect 519882 707482 555326 707718
rect 555562 707482 555646 707718
rect 555882 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 15326 707398
rect 15562 707162 15646 707398
rect 15882 707162 51326 707398
rect 51562 707162 51646 707398
rect 51882 707162 87326 707398
rect 87562 707162 87646 707398
rect 87882 707162 123326 707398
rect 123562 707162 123646 707398
rect 123882 707162 159326 707398
rect 159562 707162 159646 707398
rect 159882 707162 195326 707398
rect 195562 707162 195646 707398
rect 195882 707162 231326 707398
rect 231562 707162 231646 707398
rect 231882 707162 267326 707398
rect 267562 707162 267646 707398
rect 267882 707162 303326 707398
rect 303562 707162 303646 707398
rect 303882 707162 339326 707398
rect 339562 707162 339646 707398
rect 339882 707162 375326 707398
rect 375562 707162 375646 707398
rect 375882 707162 411326 707398
rect 411562 707162 411646 707398
rect 411882 707162 447326 707398
rect 447562 707162 447646 707398
rect 447882 707162 483326 707398
rect 483562 707162 483646 707398
rect 483882 707162 519326 707398
rect 519562 707162 519646 707398
rect 519882 707162 555326 707398
rect 555562 707162 555646 707398
rect 555882 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 10826 706758
rect 11062 706522 11146 706758
rect 11382 706522 46826 706758
rect 47062 706522 47146 706758
rect 47382 706522 82826 706758
rect 83062 706522 83146 706758
rect 83382 706522 118826 706758
rect 119062 706522 119146 706758
rect 119382 706522 154826 706758
rect 155062 706522 155146 706758
rect 155382 706522 190826 706758
rect 191062 706522 191146 706758
rect 191382 706522 226826 706758
rect 227062 706522 227146 706758
rect 227382 706522 262826 706758
rect 263062 706522 263146 706758
rect 263382 706522 298826 706758
rect 299062 706522 299146 706758
rect 299382 706522 334826 706758
rect 335062 706522 335146 706758
rect 335382 706522 370826 706758
rect 371062 706522 371146 706758
rect 371382 706522 406826 706758
rect 407062 706522 407146 706758
rect 407382 706522 442826 706758
rect 443062 706522 443146 706758
rect 443382 706522 478826 706758
rect 479062 706522 479146 706758
rect 479382 706522 514826 706758
rect 515062 706522 515146 706758
rect 515382 706522 550826 706758
rect 551062 706522 551146 706758
rect 551382 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 10826 706438
rect 11062 706202 11146 706438
rect 11382 706202 46826 706438
rect 47062 706202 47146 706438
rect 47382 706202 82826 706438
rect 83062 706202 83146 706438
rect 83382 706202 118826 706438
rect 119062 706202 119146 706438
rect 119382 706202 154826 706438
rect 155062 706202 155146 706438
rect 155382 706202 190826 706438
rect 191062 706202 191146 706438
rect 191382 706202 226826 706438
rect 227062 706202 227146 706438
rect 227382 706202 262826 706438
rect 263062 706202 263146 706438
rect 263382 706202 298826 706438
rect 299062 706202 299146 706438
rect 299382 706202 334826 706438
rect 335062 706202 335146 706438
rect 335382 706202 370826 706438
rect 371062 706202 371146 706438
rect 371382 706202 406826 706438
rect 407062 706202 407146 706438
rect 407382 706202 442826 706438
rect 443062 706202 443146 706438
rect 443382 706202 478826 706438
rect 479062 706202 479146 706438
rect 479382 706202 514826 706438
rect 515062 706202 515146 706438
rect 515382 706202 550826 706438
rect 551062 706202 551146 706438
rect 551382 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 6326 705798
rect 6562 705562 6646 705798
rect 6882 705562 42326 705798
rect 42562 705562 42646 705798
rect 42882 705562 78326 705798
rect 78562 705562 78646 705798
rect 78882 705562 114326 705798
rect 114562 705562 114646 705798
rect 114882 705562 150326 705798
rect 150562 705562 150646 705798
rect 150882 705562 186326 705798
rect 186562 705562 186646 705798
rect 186882 705562 222326 705798
rect 222562 705562 222646 705798
rect 222882 705562 258326 705798
rect 258562 705562 258646 705798
rect 258882 705562 294326 705798
rect 294562 705562 294646 705798
rect 294882 705562 330326 705798
rect 330562 705562 330646 705798
rect 330882 705562 366326 705798
rect 366562 705562 366646 705798
rect 366882 705562 402326 705798
rect 402562 705562 402646 705798
rect 402882 705562 438326 705798
rect 438562 705562 438646 705798
rect 438882 705562 474326 705798
rect 474562 705562 474646 705798
rect 474882 705562 510326 705798
rect 510562 705562 510646 705798
rect 510882 705562 546326 705798
rect 546562 705562 546646 705798
rect 546882 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 6326 705478
rect 6562 705242 6646 705478
rect 6882 705242 42326 705478
rect 42562 705242 42646 705478
rect 42882 705242 78326 705478
rect 78562 705242 78646 705478
rect 78882 705242 114326 705478
rect 114562 705242 114646 705478
rect 114882 705242 150326 705478
rect 150562 705242 150646 705478
rect 150882 705242 186326 705478
rect 186562 705242 186646 705478
rect 186882 705242 222326 705478
rect 222562 705242 222646 705478
rect 222882 705242 258326 705478
rect 258562 705242 258646 705478
rect 258882 705242 294326 705478
rect 294562 705242 294646 705478
rect 294882 705242 330326 705478
rect 330562 705242 330646 705478
rect 330882 705242 366326 705478
rect 366562 705242 366646 705478
rect 366882 705242 402326 705478
rect 402562 705242 402646 705478
rect 402882 705242 438326 705478
rect 438562 705242 438646 705478
rect 438882 705242 474326 705478
rect 474562 705242 474646 705478
rect 474882 705242 510326 705478
rect 510562 705242 510646 705478
rect 510882 705242 546326 705478
rect 546562 705242 546646 705478
rect 546882 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -4854 700954
rect -4618 700718 -4534 700954
rect -4298 700718 15326 700954
rect 15562 700718 15646 700954
rect 15882 700718 51326 700954
rect 51562 700718 51646 700954
rect 51882 700718 87326 700954
rect 87562 700718 87646 700954
rect 87882 700718 123326 700954
rect 123562 700718 123646 700954
rect 123882 700718 159326 700954
rect 159562 700718 159646 700954
rect 159882 700718 195326 700954
rect 195562 700718 195646 700954
rect 195882 700718 231326 700954
rect 231562 700718 231646 700954
rect 231882 700718 267326 700954
rect 267562 700718 267646 700954
rect 267882 700718 303326 700954
rect 303562 700718 303646 700954
rect 303882 700718 339326 700954
rect 339562 700718 339646 700954
rect 339882 700718 375326 700954
rect 375562 700718 375646 700954
rect 375882 700718 411326 700954
rect 411562 700718 411646 700954
rect 411882 700718 447326 700954
rect 447562 700718 447646 700954
rect 447882 700718 483326 700954
rect 483562 700718 483646 700954
rect 483882 700718 519326 700954
rect 519562 700718 519646 700954
rect 519882 700718 555326 700954
rect 555562 700718 555646 700954
rect 555882 700718 588222 700954
rect 588458 700718 588542 700954
rect 588778 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -4854 700634
rect -4618 700398 -4534 700634
rect -4298 700398 15326 700634
rect 15562 700398 15646 700634
rect 15882 700398 51326 700634
rect 51562 700398 51646 700634
rect 51882 700398 87326 700634
rect 87562 700398 87646 700634
rect 87882 700398 123326 700634
rect 123562 700398 123646 700634
rect 123882 700398 159326 700634
rect 159562 700398 159646 700634
rect 159882 700398 195326 700634
rect 195562 700398 195646 700634
rect 195882 700398 231326 700634
rect 231562 700398 231646 700634
rect 231882 700398 267326 700634
rect 267562 700398 267646 700634
rect 267882 700398 303326 700634
rect 303562 700398 303646 700634
rect 303882 700398 339326 700634
rect 339562 700398 339646 700634
rect 339882 700398 375326 700634
rect 375562 700398 375646 700634
rect 375882 700398 411326 700634
rect 411562 700398 411646 700634
rect 411882 700398 447326 700634
rect 447562 700398 447646 700634
rect 447882 700398 483326 700634
rect 483562 700398 483646 700634
rect 483882 700398 519326 700634
rect 519562 700398 519646 700634
rect 519882 700398 555326 700634
rect 555562 700398 555646 700634
rect 555882 700398 588222 700634
rect 588458 700398 588542 700634
rect 588778 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -3894 696454
rect -3658 696218 -3574 696454
rect -3338 696218 10826 696454
rect 11062 696218 11146 696454
rect 11382 696218 46826 696454
rect 47062 696218 47146 696454
rect 47382 696218 82826 696454
rect 83062 696218 83146 696454
rect 83382 696218 118826 696454
rect 119062 696218 119146 696454
rect 119382 696218 154826 696454
rect 155062 696218 155146 696454
rect 155382 696218 190826 696454
rect 191062 696218 191146 696454
rect 191382 696218 226826 696454
rect 227062 696218 227146 696454
rect 227382 696218 262826 696454
rect 263062 696218 263146 696454
rect 263382 696218 298826 696454
rect 299062 696218 299146 696454
rect 299382 696218 334826 696454
rect 335062 696218 335146 696454
rect 335382 696218 370826 696454
rect 371062 696218 371146 696454
rect 371382 696218 406826 696454
rect 407062 696218 407146 696454
rect 407382 696218 442826 696454
rect 443062 696218 443146 696454
rect 443382 696218 478826 696454
rect 479062 696218 479146 696454
rect 479382 696218 514826 696454
rect 515062 696218 515146 696454
rect 515382 696218 550826 696454
rect 551062 696218 551146 696454
rect 551382 696218 587262 696454
rect 587498 696218 587582 696454
rect 587818 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -3894 696134
rect -3658 695898 -3574 696134
rect -3338 695898 10826 696134
rect 11062 695898 11146 696134
rect 11382 695898 46826 696134
rect 47062 695898 47146 696134
rect 47382 695898 82826 696134
rect 83062 695898 83146 696134
rect 83382 695898 118826 696134
rect 119062 695898 119146 696134
rect 119382 695898 154826 696134
rect 155062 695898 155146 696134
rect 155382 695898 190826 696134
rect 191062 695898 191146 696134
rect 191382 695898 226826 696134
rect 227062 695898 227146 696134
rect 227382 695898 262826 696134
rect 263062 695898 263146 696134
rect 263382 695898 298826 696134
rect 299062 695898 299146 696134
rect 299382 695898 334826 696134
rect 335062 695898 335146 696134
rect 335382 695898 370826 696134
rect 371062 695898 371146 696134
rect 371382 695898 406826 696134
rect 407062 695898 407146 696134
rect 407382 695898 442826 696134
rect 443062 695898 443146 696134
rect 443382 695898 478826 696134
rect 479062 695898 479146 696134
rect 479382 695898 514826 696134
rect 515062 695898 515146 696134
rect 515382 695898 550826 696134
rect 551062 695898 551146 696134
rect 551382 695898 587262 696134
rect 587498 695898 587582 696134
rect 587818 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 691954 592650 691986
rect -8726 691718 -2934 691954
rect -2698 691718 -2614 691954
rect -2378 691718 6326 691954
rect 6562 691718 6646 691954
rect 6882 691718 42326 691954
rect 42562 691718 42646 691954
rect 42882 691718 78326 691954
rect 78562 691718 78646 691954
rect 78882 691718 114326 691954
rect 114562 691718 114646 691954
rect 114882 691718 150326 691954
rect 150562 691718 150646 691954
rect 150882 691718 186326 691954
rect 186562 691718 186646 691954
rect 186882 691718 222326 691954
rect 222562 691718 222646 691954
rect 222882 691718 258326 691954
rect 258562 691718 258646 691954
rect 258882 691718 294326 691954
rect 294562 691718 294646 691954
rect 294882 691718 330326 691954
rect 330562 691718 330646 691954
rect 330882 691718 366326 691954
rect 366562 691718 366646 691954
rect 366882 691718 402326 691954
rect 402562 691718 402646 691954
rect 402882 691718 438326 691954
rect 438562 691718 438646 691954
rect 438882 691718 474326 691954
rect 474562 691718 474646 691954
rect 474882 691718 510326 691954
rect 510562 691718 510646 691954
rect 510882 691718 546326 691954
rect 546562 691718 546646 691954
rect 546882 691718 582326 691954
rect 582562 691718 582646 691954
rect 582882 691718 586302 691954
rect 586538 691718 586622 691954
rect 586858 691718 592650 691954
rect -8726 691634 592650 691718
rect -8726 691398 -2934 691634
rect -2698 691398 -2614 691634
rect -2378 691398 6326 691634
rect 6562 691398 6646 691634
rect 6882 691398 42326 691634
rect 42562 691398 42646 691634
rect 42882 691398 78326 691634
rect 78562 691398 78646 691634
rect 78882 691398 114326 691634
rect 114562 691398 114646 691634
rect 114882 691398 150326 691634
rect 150562 691398 150646 691634
rect 150882 691398 186326 691634
rect 186562 691398 186646 691634
rect 186882 691398 222326 691634
rect 222562 691398 222646 691634
rect 222882 691398 258326 691634
rect 258562 691398 258646 691634
rect 258882 691398 294326 691634
rect 294562 691398 294646 691634
rect 294882 691398 330326 691634
rect 330562 691398 330646 691634
rect 330882 691398 366326 691634
rect 366562 691398 366646 691634
rect 366882 691398 402326 691634
rect 402562 691398 402646 691634
rect 402882 691398 438326 691634
rect 438562 691398 438646 691634
rect 438882 691398 474326 691634
rect 474562 691398 474646 691634
rect 474882 691398 510326 691634
rect 510562 691398 510646 691634
rect 510882 691398 546326 691634
rect 546562 691398 546646 691634
rect 546882 691398 582326 691634
rect 582562 691398 582646 691634
rect 582882 691398 586302 691634
rect 586538 691398 586622 691634
rect 586858 691398 592650 691634
rect -8726 691366 592650 691398
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 682954 592650 682986
rect -8726 682718 -8694 682954
rect -8458 682718 -8374 682954
rect -8138 682718 33326 682954
rect 33562 682718 33646 682954
rect 33882 682718 69326 682954
rect 69562 682718 69646 682954
rect 69882 682718 105326 682954
rect 105562 682718 105646 682954
rect 105882 682718 141326 682954
rect 141562 682718 141646 682954
rect 141882 682718 177326 682954
rect 177562 682718 177646 682954
rect 177882 682718 213326 682954
rect 213562 682718 213646 682954
rect 213882 682718 249326 682954
rect 249562 682718 249646 682954
rect 249882 682718 285326 682954
rect 285562 682718 285646 682954
rect 285882 682718 321326 682954
rect 321562 682718 321646 682954
rect 321882 682718 357326 682954
rect 357562 682718 357646 682954
rect 357882 682718 393326 682954
rect 393562 682718 393646 682954
rect 393882 682718 429326 682954
rect 429562 682718 429646 682954
rect 429882 682718 465326 682954
rect 465562 682718 465646 682954
rect 465882 682718 501326 682954
rect 501562 682718 501646 682954
rect 501882 682718 537326 682954
rect 537562 682718 537646 682954
rect 537882 682718 573326 682954
rect 573562 682718 573646 682954
rect 573882 682718 592062 682954
rect 592298 682718 592382 682954
rect 592618 682718 592650 682954
rect -8726 682634 592650 682718
rect -8726 682398 -8694 682634
rect -8458 682398 -8374 682634
rect -8138 682398 33326 682634
rect 33562 682398 33646 682634
rect 33882 682398 69326 682634
rect 69562 682398 69646 682634
rect 69882 682398 105326 682634
rect 105562 682398 105646 682634
rect 105882 682398 141326 682634
rect 141562 682398 141646 682634
rect 141882 682398 177326 682634
rect 177562 682398 177646 682634
rect 177882 682398 213326 682634
rect 213562 682398 213646 682634
rect 213882 682398 249326 682634
rect 249562 682398 249646 682634
rect 249882 682398 285326 682634
rect 285562 682398 285646 682634
rect 285882 682398 321326 682634
rect 321562 682398 321646 682634
rect 321882 682398 357326 682634
rect 357562 682398 357646 682634
rect 357882 682398 393326 682634
rect 393562 682398 393646 682634
rect 393882 682398 429326 682634
rect 429562 682398 429646 682634
rect 429882 682398 465326 682634
rect 465562 682398 465646 682634
rect 465882 682398 501326 682634
rect 501562 682398 501646 682634
rect 501882 682398 537326 682634
rect 537562 682398 537646 682634
rect 537882 682398 573326 682634
rect 573562 682398 573646 682634
rect 573882 682398 592062 682634
rect 592298 682398 592382 682634
rect 592618 682398 592650 682634
rect -8726 682366 592650 682398
rect -8726 678454 592650 678486
rect -8726 678218 -7734 678454
rect -7498 678218 -7414 678454
rect -7178 678218 28826 678454
rect 29062 678218 29146 678454
rect 29382 678218 64826 678454
rect 65062 678218 65146 678454
rect 65382 678218 100826 678454
rect 101062 678218 101146 678454
rect 101382 678218 136826 678454
rect 137062 678218 137146 678454
rect 137382 678218 172826 678454
rect 173062 678218 173146 678454
rect 173382 678218 208826 678454
rect 209062 678218 209146 678454
rect 209382 678218 244826 678454
rect 245062 678218 245146 678454
rect 245382 678218 280826 678454
rect 281062 678218 281146 678454
rect 281382 678218 316826 678454
rect 317062 678218 317146 678454
rect 317382 678218 352826 678454
rect 353062 678218 353146 678454
rect 353382 678218 388826 678454
rect 389062 678218 389146 678454
rect 389382 678218 424826 678454
rect 425062 678218 425146 678454
rect 425382 678218 460826 678454
rect 461062 678218 461146 678454
rect 461382 678218 496826 678454
rect 497062 678218 497146 678454
rect 497382 678218 532826 678454
rect 533062 678218 533146 678454
rect 533382 678218 568826 678454
rect 569062 678218 569146 678454
rect 569382 678218 591102 678454
rect 591338 678218 591422 678454
rect 591658 678218 592650 678454
rect -8726 678134 592650 678218
rect -8726 677898 -7734 678134
rect -7498 677898 -7414 678134
rect -7178 677898 28826 678134
rect 29062 677898 29146 678134
rect 29382 677898 64826 678134
rect 65062 677898 65146 678134
rect 65382 677898 100826 678134
rect 101062 677898 101146 678134
rect 101382 677898 136826 678134
rect 137062 677898 137146 678134
rect 137382 677898 172826 678134
rect 173062 677898 173146 678134
rect 173382 677898 208826 678134
rect 209062 677898 209146 678134
rect 209382 677898 244826 678134
rect 245062 677898 245146 678134
rect 245382 677898 280826 678134
rect 281062 677898 281146 678134
rect 281382 677898 316826 678134
rect 317062 677898 317146 678134
rect 317382 677898 352826 678134
rect 353062 677898 353146 678134
rect 353382 677898 388826 678134
rect 389062 677898 389146 678134
rect 389382 677898 424826 678134
rect 425062 677898 425146 678134
rect 425382 677898 460826 678134
rect 461062 677898 461146 678134
rect 461382 677898 496826 678134
rect 497062 677898 497146 678134
rect 497382 677898 532826 678134
rect 533062 677898 533146 678134
rect 533382 677898 568826 678134
rect 569062 677898 569146 678134
rect 569382 677898 591102 678134
rect 591338 677898 591422 678134
rect 591658 677898 592650 678134
rect -8726 677866 592650 677898
rect -8726 673954 592650 673986
rect -8726 673718 -6774 673954
rect -6538 673718 -6454 673954
rect -6218 673718 24326 673954
rect 24562 673718 24646 673954
rect 24882 673718 60326 673954
rect 60562 673718 60646 673954
rect 60882 673718 96326 673954
rect 96562 673718 96646 673954
rect 96882 673718 132326 673954
rect 132562 673718 132646 673954
rect 132882 673718 168326 673954
rect 168562 673718 168646 673954
rect 168882 673718 204326 673954
rect 204562 673718 204646 673954
rect 204882 673718 240326 673954
rect 240562 673718 240646 673954
rect 240882 673718 276326 673954
rect 276562 673718 276646 673954
rect 276882 673718 312326 673954
rect 312562 673718 312646 673954
rect 312882 673718 348326 673954
rect 348562 673718 348646 673954
rect 348882 673718 384326 673954
rect 384562 673718 384646 673954
rect 384882 673718 420326 673954
rect 420562 673718 420646 673954
rect 420882 673718 456326 673954
rect 456562 673718 456646 673954
rect 456882 673718 492326 673954
rect 492562 673718 492646 673954
rect 492882 673718 528326 673954
rect 528562 673718 528646 673954
rect 528882 673718 564326 673954
rect 564562 673718 564646 673954
rect 564882 673718 590142 673954
rect 590378 673718 590462 673954
rect 590698 673718 592650 673954
rect -8726 673634 592650 673718
rect -8726 673398 -6774 673634
rect -6538 673398 -6454 673634
rect -6218 673398 24326 673634
rect 24562 673398 24646 673634
rect 24882 673398 60326 673634
rect 60562 673398 60646 673634
rect 60882 673398 96326 673634
rect 96562 673398 96646 673634
rect 96882 673398 132326 673634
rect 132562 673398 132646 673634
rect 132882 673398 168326 673634
rect 168562 673398 168646 673634
rect 168882 673398 204326 673634
rect 204562 673398 204646 673634
rect 204882 673398 240326 673634
rect 240562 673398 240646 673634
rect 240882 673398 276326 673634
rect 276562 673398 276646 673634
rect 276882 673398 312326 673634
rect 312562 673398 312646 673634
rect 312882 673398 348326 673634
rect 348562 673398 348646 673634
rect 348882 673398 384326 673634
rect 384562 673398 384646 673634
rect 384882 673398 420326 673634
rect 420562 673398 420646 673634
rect 420882 673398 456326 673634
rect 456562 673398 456646 673634
rect 456882 673398 492326 673634
rect 492562 673398 492646 673634
rect 492882 673398 528326 673634
rect 528562 673398 528646 673634
rect 528882 673398 564326 673634
rect 564562 673398 564646 673634
rect 564882 673398 590142 673634
rect 590378 673398 590462 673634
rect 590698 673398 592650 673634
rect -8726 673366 592650 673398
rect -8726 669454 592650 669486
rect -8726 669218 -5814 669454
rect -5578 669218 -5494 669454
rect -5258 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 589182 669454
rect 589418 669218 589502 669454
rect 589738 669218 592650 669454
rect -8726 669134 592650 669218
rect -8726 668898 -5814 669134
rect -5578 668898 -5494 669134
rect -5258 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 589182 669134
rect 589418 668898 589502 669134
rect 589738 668898 592650 669134
rect -8726 668866 592650 668898
rect -8726 664954 592650 664986
rect -8726 664718 -4854 664954
rect -4618 664718 -4534 664954
rect -4298 664718 15326 664954
rect 15562 664718 15646 664954
rect 15882 664718 51326 664954
rect 51562 664718 51646 664954
rect 51882 664718 87326 664954
rect 87562 664718 87646 664954
rect 87882 664718 123326 664954
rect 123562 664718 123646 664954
rect 123882 664718 159326 664954
rect 159562 664718 159646 664954
rect 159882 664718 195326 664954
rect 195562 664718 195646 664954
rect 195882 664718 231326 664954
rect 231562 664718 231646 664954
rect 231882 664718 267326 664954
rect 267562 664718 267646 664954
rect 267882 664718 303326 664954
rect 303562 664718 303646 664954
rect 303882 664718 339326 664954
rect 339562 664718 339646 664954
rect 339882 664718 375326 664954
rect 375562 664718 375646 664954
rect 375882 664718 411326 664954
rect 411562 664718 411646 664954
rect 411882 664718 447326 664954
rect 447562 664718 447646 664954
rect 447882 664718 483326 664954
rect 483562 664718 483646 664954
rect 483882 664718 519326 664954
rect 519562 664718 519646 664954
rect 519882 664718 555326 664954
rect 555562 664718 555646 664954
rect 555882 664718 588222 664954
rect 588458 664718 588542 664954
rect 588778 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -4854 664634
rect -4618 664398 -4534 664634
rect -4298 664398 15326 664634
rect 15562 664398 15646 664634
rect 15882 664398 51326 664634
rect 51562 664398 51646 664634
rect 51882 664398 87326 664634
rect 87562 664398 87646 664634
rect 87882 664398 123326 664634
rect 123562 664398 123646 664634
rect 123882 664398 159326 664634
rect 159562 664398 159646 664634
rect 159882 664398 195326 664634
rect 195562 664398 195646 664634
rect 195882 664398 231326 664634
rect 231562 664398 231646 664634
rect 231882 664398 267326 664634
rect 267562 664398 267646 664634
rect 267882 664398 303326 664634
rect 303562 664398 303646 664634
rect 303882 664398 339326 664634
rect 339562 664398 339646 664634
rect 339882 664398 375326 664634
rect 375562 664398 375646 664634
rect 375882 664398 411326 664634
rect 411562 664398 411646 664634
rect 411882 664398 447326 664634
rect 447562 664398 447646 664634
rect 447882 664398 483326 664634
rect 483562 664398 483646 664634
rect 483882 664398 519326 664634
rect 519562 664398 519646 664634
rect 519882 664398 555326 664634
rect 555562 664398 555646 664634
rect 555882 664398 588222 664634
rect 588458 664398 588542 664634
rect 588778 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -3894 660454
rect -3658 660218 -3574 660454
rect -3338 660218 10826 660454
rect 11062 660218 11146 660454
rect 11382 660218 46826 660454
rect 47062 660218 47146 660454
rect 47382 660218 262826 660454
rect 263062 660218 263146 660454
rect 263382 660218 298826 660454
rect 299062 660218 299146 660454
rect 299382 660218 334826 660454
rect 335062 660218 335146 660454
rect 335382 660218 370826 660454
rect 371062 660218 371146 660454
rect 371382 660218 406826 660454
rect 407062 660218 407146 660454
rect 407382 660218 442826 660454
rect 443062 660218 443146 660454
rect 443382 660218 478826 660454
rect 479062 660218 479146 660454
rect 479382 660218 514826 660454
rect 515062 660218 515146 660454
rect 515382 660218 550826 660454
rect 551062 660218 551146 660454
rect 551382 660218 587262 660454
rect 587498 660218 587582 660454
rect 587818 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -3894 660134
rect -3658 659898 -3574 660134
rect -3338 659898 10826 660134
rect 11062 659898 11146 660134
rect 11382 659898 46826 660134
rect 47062 659898 47146 660134
rect 47382 659898 262826 660134
rect 263062 659898 263146 660134
rect 263382 659898 298826 660134
rect 299062 659898 299146 660134
rect 299382 659898 334826 660134
rect 335062 659898 335146 660134
rect 335382 659898 370826 660134
rect 371062 659898 371146 660134
rect 371382 659898 406826 660134
rect 407062 659898 407146 660134
rect 407382 659898 442826 660134
rect 443062 659898 443146 660134
rect 443382 659898 478826 660134
rect 479062 659898 479146 660134
rect 479382 659898 514826 660134
rect 515062 659898 515146 660134
rect 515382 659898 550826 660134
rect 551062 659898 551146 660134
rect 551382 659898 587262 660134
rect 587498 659898 587582 660134
rect 587818 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 655954 592650 655986
rect -8726 655718 -2934 655954
rect -2698 655718 -2614 655954
rect -2378 655718 6326 655954
rect 6562 655718 6646 655954
rect 6882 655718 42326 655954
rect 42562 655718 42646 655954
rect 42882 655718 71610 655954
rect 71846 655718 102330 655954
rect 102566 655718 133050 655954
rect 133286 655718 163770 655954
rect 164006 655718 194490 655954
rect 194726 655718 225210 655954
rect 225446 655718 258326 655954
rect 258562 655718 258646 655954
rect 258882 655718 294326 655954
rect 294562 655718 294646 655954
rect 294882 655718 330326 655954
rect 330562 655718 330646 655954
rect 330882 655718 366326 655954
rect 366562 655718 366646 655954
rect 366882 655718 402326 655954
rect 402562 655718 402646 655954
rect 402882 655718 438326 655954
rect 438562 655718 438646 655954
rect 438882 655718 474326 655954
rect 474562 655718 474646 655954
rect 474882 655718 510326 655954
rect 510562 655718 510646 655954
rect 510882 655718 546326 655954
rect 546562 655718 546646 655954
rect 546882 655718 582326 655954
rect 582562 655718 582646 655954
rect 582882 655718 586302 655954
rect 586538 655718 586622 655954
rect 586858 655718 592650 655954
rect -8726 655634 592650 655718
rect -8726 655398 -2934 655634
rect -2698 655398 -2614 655634
rect -2378 655398 6326 655634
rect 6562 655398 6646 655634
rect 6882 655398 42326 655634
rect 42562 655398 42646 655634
rect 42882 655398 71610 655634
rect 71846 655398 102330 655634
rect 102566 655398 133050 655634
rect 133286 655398 163770 655634
rect 164006 655398 194490 655634
rect 194726 655398 225210 655634
rect 225446 655398 258326 655634
rect 258562 655398 258646 655634
rect 258882 655398 294326 655634
rect 294562 655398 294646 655634
rect 294882 655398 330326 655634
rect 330562 655398 330646 655634
rect 330882 655398 366326 655634
rect 366562 655398 366646 655634
rect 366882 655398 402326 655634
rect 402562 655398 402646 655634
rect 402882 655398 438326 655634
rect 438562 655398 438646 655634
rect 438882 655398 474326 655634
rect 474562 655398 474646 655634
rect 474882 655398 510326 655634
rect 510562 655398 510646 655634
rect 510882 655398 546326 655634
rect 546562 655398 546646 655634
rect 546882 655398 582326 655634
rect 582562 655398 582646 655634
rect 582882 655398 586302 655634
rect 586538 655398 586622 655634
rect 586858 655398 592650 655634
rect -8726 655366 592650 655398
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 56250 651454
rect 56486 651218 86970 651454
rect 87206 651218 117690 651454
rect 117926 651218 148410 651454
rect 148646 651218 179130 651454
rect 179366 651218 209850 651454
rect 210086 651218 240570 651454
rect 240806 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 56250 651134
rect 56486 650898 86970 651134
rect 87206 650898 117690 651134
rect 117926 650898 148410 651134
rect 148646 650898 179130 651134
rect 179366 650898 209850 651134
rect 210086 650898 240570 651134
rect 240806 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 646954 592650 646986
rect -8726 646718 -8694 646954
rect -8458 646718 -8374 646954
rect -8138 646718 33326 646954
rect 33562 646718 33646 646954
rect 33882 646718 285326 646954
rect 285562 646718 285646 646954
rect 285882 646718 321326 646954
rect 321562 646718 321646 646954
rect 321882 646718 357326 646954
rect 357562 646718 357646 646954
rect 357882 646718 393326 646954
rect 393562 646718 393646 646954
rect 393882 646718 429326 646954
rect 429562 646718 429646 646954
rect 429882 646718 465326 646954
rect 465562 646718 465646 646954
rect 465882 646718 501326 646954
rect 501562 646718 501646 646954
rect 501882 646718 537326 646954
rect 537562 646718 537646 646954
rect 537882 646718 573326 646954
rect 573562 646718 573646 646954
rect 573882 646718 592062 646954
rect 592298 646718 592382 646954
rect 592618 646718 592650 646954
rect -8726 646634 592650 646718
rect -8726 646398 -8694 646634
rect -8458 646398 -8374 646634
rect -8138 646398 33326 646634
rect 33562 646398 33646 646634
rect 33882 646398 285326 646634
rect 285562 646398 285646 646634
rect 285882 646398 321326 646634
rect 321562 646398 321646 646634
rect 321882 646398 357326 646634
rect 357562 646398 357646 646634
rect 357882 646398 393326 646634
rect 393562 646398 393646 646634
rect 393882 646398 429326 646634
rect 429562 646398 429646 646634
rect 429882 646398 465326 646634
rect 465562 646398 465646 646634
rect 465882 646398 501326 646634
rect 501562 646398 501646 646634
rect 501882 646398 537326 646634
rect 537562 646398 537646 646634
rect 537882 646398 573326 646634
rect 573562 646398 573646 646634
rect 573882 646398 592062 646634
rect 592298 646398 592382 646634
rect 592618 646398 592650 646634
rect -8726 646366 592650 646398
rect -8726 642454 592650 642486
rect -8726 642218 -7734 642454
rect -7498 642218 -7414 642454
rect -7178 642218 28826 642454
rect 29062 642218 29146 642454
rect 29382 642361 352826 642454
rect 29382 642218 280826 642361
rect -8726 642134 280826 642218
rect -8726 641898 -7734 642134
rect -7498 641898 -7414 642134
rect -7178 641898 28826 642134
rect 29062 641898 29146 642134
rect 29382 642125 280826 642134
rect 281062 642125 281146 642361
rect 281382 642125 316826 642361
rect 317062 642125 317146 642361
rect 317382 642218 352826 642361
rect 353062 642218 353146 642454
rect 353382 642361 424826 642454
rect 353382 642218 388826 642361
rect 317382 642134 388826 642218
rect 317382 642125 352826 642134
rect 29382 641898 352826 642125
rect 353062 641898 353146 642134
rect 353382 642125 388826 642134
rect 389062 642125 389146 642361
rect 389382 642218 424826 642361
rect 425062 642218 425146 642454
rect 425382 642218 460826 642454
rect 461062 642218 461146 642454
rect 461382 642361 532826 642454
rect 461382 642218 496826 642361
rect 389382 642134 496826 642218
rect 389382 642125 424826 642134
rect 353382 641898 424826 642125
rect 425062 641898 425146 642134
rect 425382 641898 460826 642134
rect 461062 641898 461146 642134
rect 461382 642125 496826 642134
rect 497062 642125 497146 642361
rect 497382 642218 532826 642361
rect 533062 642218 533146 642454
rect 533382 642218 568826 642454
rect 569062 642218 569146 642454
rect 569382 642218 591102 642454
rect 591338 642218 591422 642454
rect 591658 642218 592650 642454
rect 497382 642134 592650 642218
rect 497382 642125 532826 642134
rect 461382 641898 532826 642125
rect 533062 641898 533146 642134
rect 533382 641898 568826 642134
rect 569062 641898 569146 642134
rect 569382 641898 591102 642134
rect 591338 641898 591422 642134
rect 591658 641898 592650 642134
rect -8726 641866 592650 641898
rect -8726 637954 592650 637986
rect -8726 637718 -6774 637954
rect -6538 637718 -6454 637954
rect -6218 637718 24326 637954
rect 24562 637718 24646 637954
rect 24882 637718 348326 637954
rect 348562 637718 348646 637954
rect 348882 637718 420326 637954
rect 420562 637718 420646 637954
rect 420882 637718 456326 637954
rect 456562 637718 456646 637954
rect 456882 637718 528326 637954
rect 528562 637718 528646 637954
rect 528882 637718 564326 637954
rect 564562 637718 564646 637954
rect 564882 637718 590142 637954
rect 590378 637718 590462 637954
rect 590698 637718 592650 637954
rect -8726 637634 592650 637718
rect -8726 637398 -6774 637634
rect -6538 637398 -6454 637634
rect -6218 637398 24326 637634
rect 24562 637398 24646 637634
rect 24882 637398 348326 637634
rect 348562 637398 348646 637634
rect 348882 637398 420326 637634
rect 420562 637398 420646 637634
rect 420882 637398 456326 637634
rect 456562 637398 456646 637634
rect 456882 637398 528326 637634
rect 528562 637398 528646 637634
rect 528882 637398 564326 637634
rect 564562 637398 564646 637634
rect 564882 637398 590142 637634
rect 590378 637398 590462 637634
rect 590698 637398 592650 637634
rect -8726 637366 592650 637398
rect -8726 633454 592650 633486
rect -8726 633218 -5814 633454
rect -5578 633218 -5494 633454
rect -5258 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 589182 633454
rect 589418 633218 589502 633454
rect 589738 633218 592650 633454
rect -8726 633134 592650 633218
rect -8726 632898 -5814 633134
rect -5578 632898 -5494 633134
rect -5258 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 589182 633134
rect 589418 632898 589502 633134
rect 589738 632898 592650 633134
rect -8726 632866 592650 632898
rect -8726 628954 592650 628986
rect -8726 628718 -4854 628954
rect -4618 628718 -4534 628954
rect -4298 628718 15326 628954
rect 15562 628718 15646 628954
rect 15882 628718 267326 628954
rect 267562 628718 267646 628954
rect 267882 628718 339326 628954
rect 339562 628718 339646 628954
rect 339882 628718 411326 628954
rect 411562 628718 411646 628954
rect 411882 628718 447326 628954
rect 447562 628718 447646 628954
rect 447882 628718 555326 628954
rect 555562 628718 555646 628954
rect 555882 628718 588222 628954
rect 588458 628718 588542 628954
rect 588778 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -4854 628634
rect -4618 628398 -4534 628634
rect -4298 628398 15326 628634
rect 15562 628398 15646 628634
rect 15882 628398 267326 628634
rect 267562 628398 267646 628634
rect 267882 628398 339326 628634
rect 339562 628398 339646 628634
rect 339882 628398 411326 628634
rect 411562 628398 411646 628634
rect 411882 628398 447326 628634
rect 447562 628398 447646 628634
rect 447882 628398 555326 628634
rect 555562 628398 555646 628634
rect 555882 628398 588222 628634
rect 588458 628398 588542 628634
rect 588778 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -3894 624454
rect -3658 624218 -3574 624454
rect -3338 624218 10826 624454
rect 11062 624218 11146 624454
rect 11382 624218 46826 624454
rect 47062 624218 47146 624454
rect 47382 624218 262826 624454
rect 263062 624218 263146 624454
rect 263382 624218 334826 624454
rect 335062 624218 335146 624454
rect 335382 624218 406826 624454
rect 407062 624218 407146 624454
rect 407382 624218 442826 624454
rect 443062 624218 443146 624454
rect 443382 624218 550826 624454
rect 551062 624218 551146 624454
rect 551382 624218 587262 624454
rect 587498 624218 587582 624454
rect 587818 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -3894 624134
rect -3658 623898 -3574 624134
rect -3338 623898 10826 624134
rect 11062 623898 11146 624134
rect 11382 623898 46826 624134
rect 47062 623898 47146 624134
rect 47382 623898 262826 624134
rect 263062 623898 263146 624134
rect 263382 623898 334826 624134
rect 335062 623898 335146 624134
rect 335382 623898 406826 624134
rect 407062 623898 407146 624134
rect 407382 623898 442826 624134
rect 443062 623898 443146 624134
rect 443382 623898 550826 624134
rect 551062 623898 551146 624134
rect 551382 623898 587262 624134
rect 587498 623898 587582 624134
rect 587818 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 619954 592650 619986
rect -8726 619718 -2934 619954
rect -2698 619718 -2614 619954
rect -2378 619718 6326 619954
rect 6562 619718 6646 619954
rect 6882 619718 42326 619954
rect 42562 619718 42646 619954
rect 42882 619718 71610 619954
rect 71846 619718 102330 619954
rect 102566 619718 133050 619954
rect 133286 619718 163770 619954
rect 164006 619718 194490 619954
rect 194726 619718 225210 619954
rect 225446 619718 258326 619954
rect 258562 619718 258646 619954
rect 258882 619718 299610 619954
rect 299846 619718 330326 619954
rect 330562 619718 330646 619954
rect 330882 619718 379610 619954
rect 379846 619718 438326 619954
rect 438562 619718 438646 619954
rect 438882 619718 474326 619954
rect 474562 619718 474646 619954
rect 474882 619718 499610 619954
rect 499846 619718 546326 619954
rect 546562 619718 546646 619954
rect 546882 619718 582326 619954
rect 582562 619718 582646 619954
rect 582882 619718 586302 619954
rect 586538 619718 586622 619954
rect 586858 619718 592650 619954
rect -8726 619634 592650 619718
rect -8726 619398 -2934 619634
rect -2698 619398 -2614 619634
rect -2378 619398 6326 619634
rect 6562 619398 6646 619634
rect 6882 619398 42326 619634
rect 42562 619398 42646 619634
rect 42882 619398 71610 619634
rect 71846 619398 102330 619634
rect 102566 619398 133050 619634
rect 133286 619398 163770 619634
rect 164006 619398 194490 619634
rect 194726 619398 225210 619634
rect 225446 619398 258326 619634
rect 258562 619398 258646 619634
rect 258882 619398 299610 619634
rect 299846 619398 330326 619634
rect 330562 619398 330646 619634
rect 330882 619398 379610 619634
rect 379846 619398 438326 619634
rect 438562 619398 438646 619634
rect 438882 619398 474326 619634
rect 474562 619398 474646 619634
rect 474882 619398 499610 619634
rect 499846 619398 546326 619634
rect 546562 619398 546646 619634
rect 546882 619398 582326 619634
rect 582562 619398 582646 619634
rect 582882 619398 586302 619634
rect 586538 619398 586622 619634
rect 586858 619398 592650 619634
rect -8726 619366 592650 619398
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 56250 615454
rect 56486 615218 86970 615454
rect 87206 615218 117690 615454
rect 117926 615218 148410 615454
rect 148646 615218 179130 615454
rect 179366 615218 209850 615454
rect 210086 615218 240570 615454
rect 240806 615218 284250 615454
rect 284486 615218 314970 615454
rect 315206 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 364250 615454
rect 364486 615218 394970 615454
rect 395206 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 484250 615454
rect 484486 615218 514970 615454
rect 515206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 56250 615134
rect 56486 614898 86970 615134
rect 87206 614898 117690 615134
rect 117926 614898 148410 615134
rect 148646 614898 179130 615134
rect 179366 614898 209850 615134
rect 210086 614898 240570 615134
rect 240806 614898 284250 615134
rect 284486 614898 314970 615134
rect 315206 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 364250 615134
rect 364486 614898 394970 615134
rect 395206 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 484250 615134
rect 484486 614898 514970 615134
rect 515206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 610954 592650 610986
rect -8726 610718 -8694 610954
rect -8458 610718 -8374 610954
rect -8138 610718 33326 610954
rect 33562 610718 33646 610954
rect 33882 610718 429326 610954
rect 429562 610718 429646 610954
rect 429882 610718 465326 610954
rect 465562 610718 465646 610954
rect 465882 610718 537326 610954
rect 537562 610718 537646 610954
rect 537882 610718 573326 610954
rect 573562 610718 573646 610954
rect 573882 610718 592062 610954
rect 592298 610718 592382 610954
rect 592618 610718 592650 610954
rect -8726 610634 592650 610718
rect -8726 610398 -8694 610634
rect -8458 610398 -8374 610634
rect -8138 610398 33326 610634
rect 33562 610398 33646 610634
rect 33882 610398 429326 610634
rect 429562 610398 429646 610634
rect 429882 610398 465326 610634
rect 465562 610398 465646 610634
rect 465882 610398 537326 610634
rect 537562 610398 537646 610634
rect 537882 610398 573326 610634
rect 573562 610398 573646 610634
rect 573882 610398 592062 610634
rect 592298 610398 592382 610634
rect 592618 610398 592650 610634
rect -8726 610366 592650 610398
rect -8726 606454 592650 606486
rect -8726 606218 -7734 606454
rect -7498 606218 -7414 606454
rect -7178 606218 28826 606454
rect 29062 606218 29146 606454
rect 29382 606218 352826 606454
rect 353062 606218 353146 606454
rect 353382 606218 424826 606454
rect 425062 606218 425146 606454
rect 425382 606218 460826 606454
rect 461062 606218 461146 606454
rect 461382 606218 532826 606454
rect 533062 606218 533146 606454
rect 533382 606218 568826 606454
rect 569062 606218 569146 606454
rect 569382 606218 591102 606454
rect 591338 606218 591422 606454
rect 591658 606218 592650 606454
rect -8726 606134 592650 606218
rect -8726 605898 -7734 606134
rect -7498 605898 -7414 606134
rect -7178 605898 28826 606134
rect 29062 605898 29146 606134
rect 29382 605898 352826 606134
rect 353062 605898 353146 606134
rect 353382 605898 424826 606134
rect 425062 605898 425146 606134
rect 425382 605898 460826 606134
rect 461062 605898 461146 606134
rect 461382 605898 532826 606134
rect 533062 605898 533146 606134
rect 533382 605898 568826 606134
rect 569062 605898 569146 606134
rect 569382 605898 591102 606134
rect 591338 605898 591422 606134
rect 591658 605898 592650 606134
rect -8726 605866 592650 605898
rect -8726 601954 592650 601986
rect -8726 601718 -6774 601954
rect -6538 601718 -6454 601954
rect -6218 601718 24326 601954
rect 24562 601718 24646 601954
rect 24882 601718 348326 601954
rect 348562 601718 348646 601954
rect 348882 601718 420326 601954
rect 420562 601718 420646 601954
rect 420882 601718 456326 601954
rect 456562 601718 456646 601954
rect 456882 601718 528326 601954
rect 528562 601718 528646 601954
rect 528882 601718 564326 601954
rect 564562 601718 564646 601954
rect 564882 601718 590142 601954
rect 590378 601718 590462 601954
rect 590698 601718 592650 601954
rect -8726 601634 592650 601718
rect -8726 601398 -6774 601634
rect -6538 601398 -6454 601634
rect -6218 601398 24326 601634
rect 24562 601398 24646 601634
rect 24882 601398 348326 601634
rect 348562 601398 348646 601634
rect 348882 601398 420326 601634
rect 420562 601398 420646 601634
rect 420882 601398 456326 601634
rect 456562 601398 456646 601634
rect 456882 601398 528326 601634
rect 528562 601398 528646 601634
rect 528882 601398 564326 601634
rect 564562 601398 564646 601634
rect 564882 601398 590142 601634
rect 590378 601398 590462 601634
rect 590698 601398 592650 601634
rect -8726 601366 592650 601398
rect -8726 597454 592650 597486
rect -8726 597218 -5814 597454
rect -5578 597218 -5494 597454
rect -5258 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 589182 597454
rect 589418 597218 589502 597454
rect 589738 597218 592650 597454
rect -8726 597134 592650 597218
rect -8726 596898 -5814 597134
rect -5578 596898 -5494 597134
rect -5258 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 589182 597134
rect 589418 596898 589502 597134
rect 589738 596898 592650 597134
rect -8726 596866 592650 596898
rect -8726 592954 592650 592986
rect -8726 592718 -4854 592954
rect -4618 592718 -4534 592954
rect -4298 592718 15326 592954
rect 15562 592718 15646 592954
rect 15882 592718 267326 592954
rect 267562 592718 267646 592954
rect 267882 592718 303326 592954
rect 303562 592718 303646 592954
rect 303882 592718 339326 592954
rect 339562 592718 339646 592954
rect 339882 592718 375326 592954
rect 375562 592718 375646 592954
rect 375882 592718 411326 592954
rect 411562 592718 411646 592954
rect 411882 592718 447326 592954
rect 447562 592718 447646 592954
rect 447882 592718 483326 592954
rect 483562 592718 483646 592954
rect 483882 592718 519326 592954
rect 519562 592718 519646 592954
rect 519882 592718 555326 592954
rect 555562 592718 555646 592954
rect 555882 592718 588222 592954
rect 588458 592718 588542 592954
rect 588778 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -4854 592634
rect -4618 592398 -4534 592634
rect -4298 592398 15326 592634
rect 15562 592398 15646 592634
rect 15882 592398 267326 592634
rect 267562 592398 267646 592634
rect 267882 592398 303326 592634
rect 303562 592398 303646 592634
rect 303882 592398 339326 592634
rect 339562 592398 339646 592634
rect 339882 592398 375326 592634
rect 375562 592398 375646 592634
rect 375882 592398 411326 592634
rect 411562 592398 411646 592634
rect 411882 592398 447326 592634
rect 447562 592398 447646 592634
rect 447882 592398 483326 592634
rect 483562 592398 483646 592634
rect 483882 592398 519326 592634
rect 519562 592398 519646 592634
rect 519882 592398 555326 592634
rect 555562 592398 555646 592634
rect 555882 592398 588222 592634
rect 588458 592398 588542 592634
rect 588778 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -3894 588454
rect -3658 588218 -3574 588454
rect -3338 588218 10826 588454
rect 11062 588218 11146 588454
rect 11382 588218 46826 588454
rect 47062 588218 47146 588454
rect 47382 588218 262826 588454
rect 263062 588218 263146 588454
rect 263382 588218 298826 588454
rect 299062 588218 299146 588454
rect 299382 588218 334826 588454
rect 335062 588218 335146 588454
rect 335382 588218 370826 588454
rect 371062 588218 371146 588454
rect 371382 588218 406826 588454
rect 407062 588218 407146 588454
rect 407382 588218 442826 588454
rect 443062 588218 443146 588454
rect 443382 588218 478826 588454
rect 479062 588218 479146 588454
rect 479382 588218 514826 588454
rect 515062 588218 515146 588454
rect 515382 588218 550826 588454
rect 551062 588218 551146 588454
rect 551382 588218 587262 588454
rect 587498 588218 587582 588454
rect 587818 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -3894 588134
rect -3658 587898 -3574 588134
rect -3338 587898 10826 588134
rect 11062 587898 11146 588134
rect 11382 587898 46826 588134
rect 47062 587898 47146 588134
rect 47382 587898 262826 588134
rect 263062 587898 263146 588134
rect 263382 587898 298826 588134
rect 299062 587898 299146 588134
rect 299382 587898 334826 588134
rect 335062 587898 335146 588134
rect 335382 587898 370826 588134
rect 371062 587898 371146 588134
rect 371382 587898 406826 588134
rect 407062 587898 407146 588134
rect 407382 587898 442826 588134
rect 443062 587898 443146 588134
rect 443382 587898 478826 588134
rect 479062 587898 479146 588134
rect 479382 587898 514826 588134
rect 515062 587898 515146 588134
rect 515382 587898 550826 588134
rect 551062 587898 551146 588134
rect 551382 587898 587262 588134
rect 587498 587898 587582 588134
rect 587818 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 583954 592650 583986
rect -8726 583718 -2934 583954
rect -2698 583718 -2614 583954
rect -2378 583718 6326 583954
rect 6562 583718 6646 583954
rect 6882 583718 42326 583954
rect 42562 583718 42646 583954
rect 42882 583718 71610 583954
rect 71846 583718 102330 583954
rect 102566 583718 133050 583954
rect 133286 583718 163770 583954
rect 164006 583718 194490 583954
rect 194726 583718 225210 583954
rect 225446 583718 258326 583954
rect 258562 583718 258646 583954
rect 258882 583718 294326 583954
rect 294562 583718 294646 583954
rect 294882 583718 330326 583954
rect 330562 583718 330646 583954
rect 330882 583718 438326 583954
rect 438562 583718 438646 583954
rect 438882 583718 474326 583954
rect 474562 583718 474646 583954
rect 474882 583718 510326 583954
rect 510562 583718 510646 583954
rect 510882 583718 546326 583954
rect 546562 583718 546646 583954
rect 546882 583718 582326 583954
rect 582562 583718 582646 583954
rect 582882 583718 586302 583954
rect 586538 583718 586622 583954
rect 586858 583718 592650 583954
rect -8726 583634 592650 583718
rect -8726 583398 -2934 583634
rect -2698 583398 -2614 583634
rect -2378 583398 6326 583634
rect 6562 583398 6646 583634
rect 6882 583398 42326 583634
rect 42562 583398 42646 583634
rect 42882 583398 71610 583634
rect 71846 583398 102330 583634
rect 102566 583398 133050 583634
rect 133286 583398 163770 583634
rect 164006 583398 194490 583634
rect 194726 583398 225210 583634
rect 225446 583398 258326 583634
rect 258562 583398 258646 583634
rect 258882 583398 294326 583634
rect 294562 583398 294646 583634
rect 294882 583398 330326 583634
rect 330562 583398 330646 583634
rect 330882 583398 438326 583634
rect 438562 583398 438646 583634
rect 438882 583398 474326 583634
rect 474562 583398 474646 583634
rect 474882 583398 510326 583634
rect 510562 583398 510646 583634
rect 510882 583398 546326 583634
rect 546562 583398 546646 583634
rect 546882 583398 582326 583634
rect 582562 583398 582646 583634
rect 582882 583398 586302 583634
rect 586538 583398 586622 583634
rect 586858 583398 592650 583634
rect -8726 583366 592650 583398
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 56250 579454
rect 56486 579218 86970 579454
rect 87206 579218 117690 579454
rect 117926 579218 148410 579454
rect 148646 579218 179130 579454
rect 179366 579218 209850 579454
rect 210086 579218 240570 579454
rect 240806 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 56250 579134
rect 56486 578898 86970 579134
rect 87206 578898 117690 579134
rect 117926 578898 148410 579134
rect 148646 578898 179130 579134
rect 179366 578898 209850 579134
rect 210086 578898 240570 579134
rect 240806 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 574954 592650 574986
rect -8726 574718 -8694 574954
rect -8458 574718 -8374 574954
rect -8138 574718 33326 574954
rect 33562 574718 33646 574954
rect 33882 574718 429326 574954
rect 429562 574718 429646 574954
rect 429882 574718 465326 574954
rect 465562 574718 465646 574954
rect 465882 574718 537326 574954
rect 537562 574718 537646 574954
rect 537882 574718 573326 574954
rect 573562 574718 573646 574954
rect 573882 574718 592062 574954
rect 592298 574718 592382 574954
rect 592618 574718 592650 574954
rect -8726 574634 592650 574718
rect -8726 574398 -8694 574634
rect -8458 574398 -8374 574634
rect -8138 574398 33326 574634
rect 33562 574398 33646 574634
rect 33882 574398 429326 574634
rect 429562 574398 429646 574634
rect 429882 574398 465326 574634
rect 465562 574398 465646 574634
rect 465882 574398 537326 574634
rect 537562 574398 537646 574634
rect 537882 574398 573326 574634
rect 573562 574398 573646 574634
rect 573882 574398 592062 574634
rect 592298 574398 592382 574634
rect 592618 574398 592650 574634
rect -8726 574366 592650 574398
rect -8726 570454 592650 570486
rect -8726 570218 -7734 570454
rect -7498 570218 -7414 570454
rect -7178 570218 28826 570454
rect 29062 570218 29146 570454
rect 29382 570218 352826 570454
rect 353062 570218 353146 570454
rect 353382 570218 424826 570454
rect 425062 570218 425146 570454
rect 425382 570218 460826 570454
rect 461062 570218 461146 570454
rect 461382 570218 532826 570454
rect 533062 570218 533146 570454
rect 533382 570218 568826 570454
rect 569062 570218 569146 570454
rect 569382 570218 591102 570454
rect 591338 570218 591422 570454
rect 591658 570218 592650 570454
rect -8726 570134 592650 570218
rect -8726 569898 -7734 570134
rect -7498 569898 -7414 570134
rect -7178 569898 28826 570134
rect 29062 569898 29146 570134
rect 29382 569898 352826 570134
rect 353062 569898 353146 570134
rect 353382 569898 424826 570134
rect 425062 569898 425146 570134
rect 425382 569898 460826 570134
rect 461062 569898 461146 570134
rect 461382 569898 532826 570134
rect 533062 569898 533146 570134
rect 533382 569898 568826 570134
rect 569062 569898 569146 570134
rect 569382 569898 591102 570134
rect 591338 569898 591422 570134
rect 591658 569898 592650 570134
rect -8726 569866 592650 569898
rect -8726 565954 592650 565986
rect -8726 565718 -6774 565954
rect -6538 565718 -6454 565954
rect -6218 565718 24326 565954
rect 24562 565718 24646 565954
rect 24882 565718 348326 565954
rect 348562 565718 348646 565954
rect 348882 565718 420326 565954
rect 420562 565718 420646 565954
rect 420882 565718 456326 565954
rect 456562 565718 456646 565954
rect 456882 565718 528326 565954
rect 528562 565718 528646 565954
rect 528882 565718 564326 565954
rect 564562 565718 564646 565954
rect 564882 565718 590142 565954
rect 590378 565718 590462 565954
rect 590698 565718 592650 565954
rect -8726 565634 592650 565718
rect -8726 565398 -6774 565634
rect -6538 565398 -6454 565634
rect -6218 565398 24326 565634
rect 24562 565398 24646 565634
rect 24882 565398 348326 565634
rect 348562 565398 348646 565634
rect 348882 565398 420326 565634
rect 420562 565398 420646 565634
rect 420882 565398 456326 565634
rect 456562 565398 456646 565634
rect 456882 565398 528326 565634
rect 528562 565398 528646 565634
rect 528882 565398 564326 565634
rect 564562 565398 564646 565634
rect 564882 565398 590142 565634
rect 590378 565398 590462 565634
rect 590698 565398 592650 565634
rect -8726 565366 592650 565398
rect -8726 561454 592650 561486
rect -8726 561218 -5814 561454
rect -5578 561218 -5494 561454
rect -5258 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 589182 561454
rect 589418 561218 589502 561454
rect 589738 561218 592650 561454
rect -8726 561134 592650 561218
rect -8726 560898 -5814 561134
rect -5578 560898 -5494 561134
rect -5258 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 589182 561134
rect 589418 560898 589502 561134
rect 589738 560898 592650 561134
rect -8726 560866 592650 560898
rect -8726 556954 592650 556986
rect -8726 556718 -4854 556954
rect -4618 556718 -4534 556954
rect -4298 556718 15326 556954
rect 15562 556718 15646 556954
rect 15882 556718 267326 556954
rect 267562 556718 267646 556954
rect 267882 556718 303326 556954
rect 303562 556718 303646 556954
rect 303882 556718 339326 556954
rect 339562 556718 339646 556954
rect 339882 556718 375326 556954
rect 375562 556718 375646 556954
rect 375882 556718 411326 556954
rect 411562 556718 411646 556954
rect 411882 556718 447326 556954
rect 447562 556718 447646 556954
rect 447882 556718 483326 556954
rect 483562 556718 483646 556954
rect 483882 556718 519326 556954
rect 519562 556718 519646 556954
rect 519882 556718 555326 556954
rect 555562 556718 555646 556954
rect 555882 556718 588222 556954
rect 588458 556718 588542 556954
rect 588778 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -4854 556634
rect -4618 556398 -4534 556634
rect -4298 556398 15326 556634
rect 15562 556398 15646 556634
rect 15882 556398 267326 556634
rect 267562 556398 267646 556634
rect 267882 556398 303326 556634
rect 303562 556398 303646 556634
rect 303882 556398 339326 556634
rect 339562 556398 339646 556634
rect 339882 556398 375326 556634
rect 375562 556398 375646 556634
rect 375882 556398 411326 556634
rect 411562 556398 411646 556634
rect 411882 556398 447326 556634
rect 447562 556398 447646 556634
rect 447882 556398 483326 556634
rect 483562 556398 483646 556634
rect 483882 556398 519326 556634
rect 519562 556398 519646 556634
rect 519882 556398 555326 556634
rect 555562 556398 555646 556634
rect 555882 556398 588222 556634
rect 588458 556398 588542 556634
rect 588778 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -3894 552454
rect -3658 552218 -3574 552454
rect -3338 552218 10826 552454
rect 11062 552218 11146 552454
rect 11382 552218 46826 552454
rect 47062 552218 47146 552454
rect 47382 552218 262826 552454
rect 263062 552218 263146 552454
rect 263382 552218 298826 552454
rect 299062 552218 299146 552454
rect 299382 552218 334826 552454
rect 335062 552218 335146 552454
rect 335382 552361 406826 552454
rect 335382 552218 370826 552361
rect -8726 552134 370826 552218
rect -8726 551898 -3894 552134
rect -3658 551898 -3574 552134
rect -3338 551898 10826 552134
rect 11062 551898 11146 552134
rect 11382 551898 46826 552134
rect 47062 551898 47146 552134
rect 47382 551898 262826 552134
rect 263062 551898 263146 552134
rect 263382 551898 298826 552134
rect 299062 551898 299146 552134
rect 299382 551898 334826 552134
rect 335062 551898 335146 552134
rect 335382 552125 370826 552134
rect 371062 552125 371146 552361
rect 371382 552218 406826 552361
rect 407062 552218 407146 552454
rect 407382 552218 442826 552454
rect 443062 552218 443146 552454
rect 443382 552218 478826 552454
rect 479062 552218 479146 552454
rect 479382 552218 514826 552454
rect 515062 552218 515146 552454
rect 515382 552218 550826 552454
rect 551062 552218 551146 552454
rect 551382 552218 587262 552454
rect 587498 552218 587582 552454
rect 587818 552218 592650 552454
rect 371382 552134 592650 552218
rect 371382 552125 406826 552134
rect 335382 551898 406826 552125
rect 407062 551898 407146 552134
rect 407382 551898 442826 552134
rect 443062 551898 443146 552134
rect 443382 551898 478826 552134
rect 479062 551898 479146 552134
rect 479382 551898 514826 552134
rect 515062 551898 515146 552134
rect 515382 551898 550826 552134
rect 551062 551898 551146 552134
rect 551382 551898 587262 552134
rect 587498 551898 587582 552134
rect 587818 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 547954 592650 547986
rect -8726 547718 -2934 547954
rect -2698 547718 -2614 547954
rect -2378 547718 6326 547954
rect 6562 547718 6646 547954
rect 6882 547718 42326 547954
rect 42562 547718 42646 547954
rect 42882 547718 71610 547954
rect 71846 547718 102330 547954
rect 102566 547718 133050 547954
rect 133286 547718 163770 547954
rect 164006 547718 194490 547954
rect 194726 547718 225210 547954
rect 225446 547718 258326 547954
rect 258562 547718 258646 547954
rect 258882 547718 294326 547954
rect 294562 547718 294646 547954
rect 294882 547718 330326 547954
rect 330562 547718 330646 547954
rect 330882 547718 438326 547954
rect 438562 547718 438646 547954
rect 438882 547718 474326 547954
rect 474562 547718 474646 547954
rect 474882 547718 510326 547954
rect 510562 547718 510646 547954
rect 510882 547718 546326 547954
rect 546562 547718 546646 547954
rect 546882 547718 582326 547954
rect 582562 547718 582646 547954
rect 582882 547718 586302 547954
rect 586538 547718 586622 547954
rect 586858 547718 592650 547954
rect -8726 547634 592650 547718
rect -8726 547398 -2934 547634
rect -2698 547398 -2614 547634
rect -2378 547398 6326 547634
rect 6562 547398 6646 547634
rect 6882 547398 42326 547634
rect 42562 547398 42646 547634
rect 42882 547398 71610 547634
rect 71846 547398 102330 547634
rect 102566 547398 133050 547634
rect 133286 547398 163770 547634
rect 164006 547398 194490 547634
rect 194726 547398 225210 547634
rect 225446 547398 258326 547634
rect 258562 547398 258646 547634
rect 258882 547398 294326 547634
rect 294562 547398 294646 547634
rect 294882 547398 330326 547634
rect 330562 547398 330646 547634
rect 330882 547398 438326 547634
rect 438562 547398 438646 547634
rect 438882 547398 474326 547634
rect 474562 547398 474646 547634
rect 474882 547398 510326 547634
rect 510562 547398 510646 547634
rect 510882 547398 546326 547634
rect 546562 547398 546646 547634
rect 546882 547398 582326 547634
rect 582562 547398 582646 547634
rect 582882 547398 586302 547634
rect 586538 547398 586622 547634
rect 586858 547398 592650 547634
rect -8726 547366 592650 547398
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 56250 543454
rect 56486 543218 86970 543454
rect 87206 543218 117690 543454
rect 117926 543218 148410 543454
rect 148646 543218 179130 543454
rect 179366 543218 209850 543454
rect 210086 543218 240570 543454
rect 240806 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 364250 543454
rect 364486 543218 394970 543454
rect 395206 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 56250 543134
rect 56486 542898 86970 543134
rect 87206 542898 117690 543134
rect 117926 542898 148410 543134
rect 148646 542898 179130 543134
rect 179366 542898 209850 543134
rect 210086 542898 240570 543134
rect 240806 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 364250 543134
rect 364486 542898 394970 543134
rect 395206 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 538954 592650 538986
rect -8726 538718 -8694 538954
rect -8458 538718 -8374 538954
rect -8138 538718 33326 538954
rect 33562 538718 33646 538954
rect 33882 538718 429326 538954
rect 429562 538718 429646 538954
rect 429882 538718 465326 538954
rect 465562 538718 465646 538954
rect 465882 538718 537326 538954
rect 537562 538718 537646 538954
rect 537882 538718 573326 538954
rect 573562 538718 573646 538954
rect 573882 538718 592062 538954
rect 592298 538718 592382 538954
rect 592618 538718 592650 538954
rect -8726 538634 592650 538718
rect -8726 538398 -8694 538634
rect -8458 538398 -8374 538634
rect -8138 538398 33326 538634
rect 33562 538398 33646 538634
rect 33882 538398 429326 538634
rect 429562 538398 429646 538634
rect 429882 538398 465326 538634
rect 465562 538398 465646 538634
rect 465882 538398 537326 538634
rect 537562 538398 537646 538634
rect 537882 538398 573326 538634
rect 573562 538398 573646 538634
rect 573882 538398 592062 538634
rect 592298 538398 592382 538634
rect 592618 538398 592650 538634
rect -8726 538366 592650 538398
rect -8726 534454 592650 534486
rect -8726 534218 -7734 534454
rect -7498 534218 -7414 534454
rect -7178 534218 28826 534454
rect 29062 534218 29146 534454
rect 29382 534218 352826 534454
rect 353062 534218 353146 534454
rect 353382 534218 424826 534454
rect 425062 534218 425146 534454
rect 425382 534218 460826 534454
rect 461062 534218 461146 534454
rect 461382 534218 532826 534454
rect 533062 534218 533146 534454
rect 533382 534218 568826 534454
rect 569062 534218 569146 534454
rect 569382 534218 591102 534454
rect 591338 534218 591422 534454
rect 591658 534218 592650 534454
rect -8726 534134 592650 534218
rect -8726 533898 -7734 534134
rect -7498 533898 -7414 534134
rect -7178 533898 28826 534134
rect 29062 533898 29146 534134
rect 29382 533898 352826 534134
rect 353062 533898 353146 534134
rect 353382 533898 424826 534134
rect 425062 533898 425146 534134
rect 425382 533898 460826 534134
rect 461062 533898 461146 534134
rect 461382 533898 532826 534134
rect 533062 533898 533146 534134
rect 533382 533898 568826 534134
rect 569062 533898 569146 534134
rect 569382 533898 591102 534134
rect 591338 533898 591422 534134
rect 591658 533898 592650 534134
rect -8726 533866 592650 533898
rect -8726 529954 592650 529986
rect -8726 529718 -6774 529954
rect -6538 529718 -6454 529954
rect -6218 529718 24326 529954
rect 24562 529718 24646 529954
rect 24882 529718 348326 529954
rect 348562 529718 348646 529954
rect 348882 529718 420326 529954
rect 420562 529718 420646 529954
rect 420882 529718 456326 529954
rect 456562 529718 456646 529954
rect 456882 529718 528326 529954
rect 528562 529718 528646 529954
rect 528882 529718 564326 529954
rect 564562 529718 564646 529954
rect 564882 529718 590142 529954
rect 590378 529718 590462 529954
rect 590698 529718 592650 529954
rect -8726 529634 592650 529718
rect -8726 529398 -6774 529634
rect -6538 529398 -6454 529634
rect -6218 529398 24326 529634
rect 24562 529398 24646 529634
rect 24882 529398 348326 529634
rect 348562 529398 348646 529634
rect 348882 529398 420326 529634
rect 420562 529398 420646 529634
rect 420882 529398 456326 529634
rect 456562 529398 456646 529634
rect 456882 529398 528326 529634
rect 528562 529398 528646 529634
rect 528882 529398 564326 529634
rect 564562 529398 564646 529634
rect 564882 529398 590142 529634
rect 590378 529398 590462 529634
rect 590698 529398 592650 529634
rect -8726 529366 592650 529398
rect -8726 525454 592650 525486
rect -8726 525218 -5814 525454
rect -5578 525218 -5494 525454
rect -5258 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 589182 525454
rect 589418 525218 589502 525454
rect 589738 525218 592650 525454
rect -8726 525134 592650 525218
rect -8726 524898 -5814 525134
rect -5578 524898 -5494 525134
rect -5258 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 589182 525134
rect 589418 524898 589502 525134
rect 589738 524898 592650 525134
rect -8726 524866 592650 524898
rect -8726 520954 592650 520986
rect -8726 520718 -4854 520954
rect -4618 520718 -4534 520954
rect -4298 520718 15326 520954
rect 15562 520718 15646 520954
rect 15882 520718 267326 520954
rect 267562 520718 267646 520954
rect 267882 520718 339326 520954
rect 339562 520718 339646 520954
rect 339882 520718 411326 520954
rect 411562 520718 411646 520954
rect 411882 520718 447326 520954
rect 447562 520718 447646 520954
rect 447882 520718 555326 520954
rect 555562 520718 555646 520954
rect 555882 520718 588222 520954
rect 588458 520718 588542 520954
rect 588778 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -4854 520634
rect -4618 520398 -4534 520634
rect -4298 520398 15326 520634
rect 15562 520398 15646 520634
rect 15882 520398 267326 520634
rect 267562 520398 267646 520634
rect 267882 520398 339326 520634
rect 339562 520398 339646 520634
rect 339882 520398 411326 520634
rect 411562 520398 411646 520634
rect 411882 520398 447326 520634
rect 447562 520398 447646 520634
rect 447882 520398 555326 520634
rect 555562 520398 555646 520634
rect 555882 520398 588222 520634
rect 588458 520398 588542 520634
rect 588778 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -3894 516454
rect -3658 516218 -3574 516454
rect -3338 516218 10826 516454
rect 11062 516218 11146 516454
rect 11382 516218 46826 516454
rect 47062 516218 47146 516454
rect 47382 516218 262826 516454
rect 263062 516218 263146 516454
rect 263382 516218 334826 516454
rect 335062 516218 335146 516454
rect 335382 516218 406826 516454
rect 407062 516218 407146 516454
rect 407382 516218 442826 516454
rect 443062 516218 443146 516454
rect 443382 516218 550826 516454
rect 551062 516218 551146 516454
rect 551382 516218 587262 516454
rect 587498 516218 587582 516454
rect 587818 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -3894 516134
rect -3658 515898 -3574 516134
rect -3338 515898 10826 516134
rect 11062 515898 11146 516134
rect 11382 515898 46826 516134
rect 47062 515898 47146 516134
rect 47382 515898 262826 516134
rect 263062 515898 263146 516134
rect 263382 515898 334826 516134
rect 335062 515898 335146 516134
rect 335382 515898 406826 516134
rect 407062 515898 407146 516134
rect 407382 515898 442826 516134
rect 443062 515898 443146 516134
rect 443382 515898 550826 516134
rect 551062 515898 551146 516134
rect 551382 515898 587262 516134
rect 587498 515898 587582 516134
rect 587818 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 511954 592650 511986
rect -8726 511718 -2934 511954
rect -2698 511718 -2614 511954
rect -2378 511718 6326 511954
rect 6562 511718 6646 511954
rect 6882 511718 42326 511954
rect 42562 511718 42646 511954
rect 42882 511718 71610 511954
rect 71846 511718 102330 511954
rect 102566 511718 133050 511954
rect 133286 511718 163770 511954
rect 164006 511718 194490 511954
rect 194726 511718 225210 511954
rect 225446 511718 258326 511954
rect 258562 511718 258646 511954
rect 258882 511718 299610 511954
rect 299846 511718 330326 511954
rect 330562 511718 330646 511954
rect 330882 511718 379610 511954
rect 379846 511718 438326 511954
rect 438562 511718 438646 511954
rect 438882 511718 474326 511954
rect 474562 511718 474646 511954
rect 474882 511718 499610 511954
rect 499846 511718 546326 511954
rect 546562 511718 546646 511954
rect 546882 511718 582326 511954
rect 582562 511718 582646 511954
rect 582882 511718 586302 511954
rect 586538 511718 586622 511954
rect 586858 511718 592650 511954
rect -8726 511634 592650 511718
rect -8726 511398 -2934 511634
rect -2698 511398 -2614 511634
rect -2378 511398 6326 511634
rect 6562 511398 6646 511634
rect 6882 511398 42326 511634
rect 42562 511398 42646 511634
rect 42882 511398 71610 511634
rect 71846 511398 102330 511634
rect 102566 511398 133050 511634
rect 133286 511398 163770 511634
rect 164006 511398 194490 511634
rect 194726 511398 225210 511634
rect 225446 511398 258326 511634
rect 258562 511398 258646 511634
rect 258882 511398 299610 511634
rect 299846 511398 330326 511634
rect 330562 511398 330646 511634
rect 330882 511398 379610 511634
rect 379846 511398 438326 511634
rect 438562 511398 438646 511634
rect 438882 511398 474326 511634
rect 474562 511398 474646 511634
rect 474882 511398 499610 511634
rect 499846 511398 546326 511634
rect 546562 511398 546646 511634
rect 546882 511398 582326 511634
rect 582562 511398 582646 511634
rect 582882 511398 586302 511634
rect 586538 511398 586622 511634
rect 586858 511398 592650 511634
rect -8726 511366 592650 511398
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 56250 507454
rect 56486 507218 86970 507454
rect 87206 507218 117690 507454
rect 117926 507218 148410 507454
rect 148646 507218 179130 507454
rect 179366 507218 209850 507454
rect 210086 507218 240570 507454
rect 240806 507218 284250 507454
rect 284486 507218 314970 507454
rect 315206 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 364250 507454
rect 364486 507218 394970 507454
rect 395206 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 484250 507454
rect 484486 507218 514970 507454
rect 515206 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 56250 507134
rect 56486 506898 86970 507134
rect 87206 506898 117690 507134
rect 117926 506898 148410 507134
rect 148646 506898 179130 507134
rect 179366 506898 209850 507134
rect 210086 506898 240570 507134
rect 240806 506898 284250 507134
rect 284486 506898 314970 507134
rect 315206 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 364250 507134
rect 364486 506898 394970 507134
rect 395206 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 484250 507134
rect 484486 506898 514970 507134
rect 515206 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 502954 592650 502986
rect -8726 502718 -8694 502954
rect -8458 502718 -8374 502954
rect -8138 502718 33326 502954
rect 33562 502718 33646 502954
rect 33882 502718 429326 502954
rect 429562 502718 429646 502954
rect 429882 502718 465326 502954
rect 465562 502718 465646 502954
rect 465882 502718 537326 502954
rect 537562 502718 537646 502954
rect 537882 502718 573326 502954
rect 573562 502718 573646 502954
rect 573882 502718 592062 502954
rect 592298 502718 592382 502954
rect 592618 502718 592650 502954
rect -8726 502634 592650 502718
rect -8726 502398 -8694 502634
rect -8458 502398 -8374 502634
rect -8138 502398 33326 502634
rect 33562 502398 33646 502634
rect 33882 502398 429326 502634
rect 429562 502398 429646 502634
rect 429882 502398 465326 502634
rect 465562 502398 465646 502634
rect 465882 502398 537326 502634
rect 537562 502398 537646 502634
rect 537882 502398 573326 502634
rect 573562 502398 573646 502634
rect 573882 502398 592062 502634
rect 592298 502398 592382 502634
rect 592618 502398 592650 502634
rect -8726 502366 592650 502398
rect -8726 498454 592650 498486
rect -8726 498218 -7734 498454
rect -7498 498218 -7414 498454
rect -7178 498218 28826 498454
rect 29062 498218 29146 498454
rect 29382 498218 352826 498454
rect 353062 498218 353146 498454
rect 353382 498218 424826 498454
rect 425062 498218 425146 498454
rect 425382 498218 460826 498454
rect 461062 498218 461146 498454
rect 461382 498218 532826 498454
rect 533062 498218 533146 498454
rect 533382 498218 568826 498454
rect 569062 498218 569146 498454
rect 569382 498218 591102 498454
rect 591338 498218 591422 498454
rect 591658 498218 592650 498454
rect -8726 498134 592650 498218
rect -8726 497898 -7734 498134
rect -7498 497898 -7414 498134
rect -7178 497898 28826 498134
rect 29062 497898 29146 498134
rect 29382 497898 352826 498134
rect 353062 497898 353146 498134
rect 353382 497898 424826 498134
rect 425062 497898 425146 498134
rect 425382 497898 460826 498134
rect 461062 497898 461146 498134
rect 461382 497898 532826 498134
rect 533062 497898 533146 498134
rect 533382 497898 568826 498134
rect 569062 497898 569146 498134
rect 569382 497898 591102 498134
rect 591338 497898 591422 498134
rect 591658 497898 592650 498134
rect -8726 497866 592650 497898
rect -8726 493954 592650 493986
rect -8726 493718 -6774 493954
rect -6538 493718 -6454 493954
rect -6218 493718 24326 493954
rect 24562 493718 24646 493954
rect 24882 493718 276326 493954
rect 276562 493718 276646 493954
rect 276882 493718 312326 493954
rect 312562 493718 312646 493954
rect 312882 493718 348326 493954
rect 348562 493718 348646 493954
rect 348882 493718 384326 493954
rect 384562 493718 384646 493954
rect 384882 493718 420326 493954
rect 420562 493718 420646 493954
rect 420882 493718 456326 493954
rect 456562 493718 456646 493954
rect 456882 493718 492326 493954
rect 492562 493718 492646 493954
rect 492882 493718 528326 493954
rect 528562 493718 528646 493954
rect 528882 493718 564326 493954
rect 564562 493718 564646 493954
rect 564882 493718 590142 493954
rect 590378 493718 590462 493954
rect 590698 493718 592650 493954
rect -8726 493634 592650 493718
rect -8726 493398 -6774 493634
rect -6538 493398 -6454 493634
rect -6218 493398 24326 493634
rect 24562 493398 24646 493634
rect 24882 493398 276326 493634
rect 276562 493398 276646 493634
rect 276882 493398 312326 493634
rect 312562 493398 312646 493634
rect 312882 493398 348326 493634
rect 348562 493398 348646 493634
rect 348882 493398 384326 493634
rect 384562 493398 384646 493634
rect 384882 493398 420326 493634
rect 420562 493398 420646 493634
rect 420882 493398 456326 493634
rect 456562 493398 456646 493634
rect 456882 493398 492326 493634
rect 492562 493398 492646 493634
rect 492882 493398 528326 493634
rect 528562 493398 528646 493634
rect 528882 493398 564326 493634
rect 564562 493398 564646 493634
rect 564882 493398 590142 493634
rect 590378 493398 590462 493634
rect 590698 493398 592650 493634
rect -8726 493366 592650 493398
rect -8726 489454 592650 489486
rect -8726 489218 -5814 489454
rect -5578 489218 -5494 489454
rect -5258 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 589182 489454
rect 589418 489218 589502 489454
rect 589738 489218 592650 489454
rect -8726 489134 592650 489218
rect -8726 488898 -5814 489134
rect -5578 488898 -5494 489134
rect -5258 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 589182 489134
rect 589418 488898 589502 489134
rect 589738 488898 592650 489134
rect -8726 488866 592650 488898
rect -8726 484954 592650 484986
rect -8726 484718 -4854 484954
rect -4618 484718 -4534 484954
rect -4298 484718 15326 484954
rect 15562 484718 15646 484954
rect 15882 484718 267326 484954
rect 267562 484718 267646 484954
rect 267882 484718 303326 484954
rect 303562 484718 303646 484954
rect 303882 484718 339326 484954
rect 339562 484718 339646 484954
rect 339882 484718 375326 484954
rect 375562 484718 375646 484954
rect 375882 484718 411326 484954
rect 411562 484718 411646 484954
rect 411882 484718 447326 484954
rect 447562 484718 447646 484954
rect 447882 484718 483326 484954
rect 483562 484718 483646 484954
rect 483882 484718 519326 484954
rect 519562 484718 519646 484954
rect 519882 484718 555326 484954
rect 555562 484718 555646 484954
rect 555882 484718 588222 484954
rect 588458 484718 588542 484954
rect 588778 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -4854 484634
rect -4618 484398 -4534 484634
rect -4298 484398 15326 484634
rect 15562 484398 15646 484634
rect 15882 484398 267326 484634
rect 267562 484398 267646 484634
rect 267882 484398 303326 484634
rect 303562 484398 303646 484634
rect 303882 484398 339326 484634
rect 339562 484398 339646 484634
rect 339882 484398 375326 484634
rect 375562 484398 375646 484634
rect 375882 484398 411326 484634
rect 411562 484398 411646 484634
rect 411882 484398 447326 484634
rect 447562 484398 447646 484634
rect 447882 484398 483326 484634
rect 483562 484398 483646 484634
rect 483882 484398 519326 484634
rect 519562 484398 519646 484634
rect 519882 484398 555326 484634
rect 555562 484398 555646 484634
rect 555882 484398 588222 484634
rect 588458 484398 588542 484634
rect 588778 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -3894 480454
rect -3658 480218 -3574 480454
rect -3338 480218 10826 480454
rect 11062 480218 11146 480454
rect 11382 480218 46826 480454
rect 47062 480218 47146 480454
rect 47382 480218 262826 480454
rect 263062 480218 263146 480454
rect 263382 480218 298826 480454
rect 299062 480218 299146 480454
rect 299382 480218 334826 480454
rect 335062 480218 335146 480454
rect 335382 480218 370826 480454
rect 371062 480218 371146 480454
rect 371382 480218 406826 480454
rect 407062 480218 407146 480454
rect 407382 480218 442826 480454
rect 443062 480218 443146 480454
rect 443382 480218 478826 480454
rect 479062 480218 479146 480454
rect 479382 480218 514826 480454
rect 515062 480218 515146 480454
rect 515382 480218 550826 480454
rect 551062 480218 551146 480454
rect 551382 480218 587262 480454
rect 587498 480218 587582 480454
rect 587818 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -3894 480134
rect -3658 479898 -3574 480134
rect -3338 479898 10826 480134
rect 11062 479898 11146 480134
rect 11382 479898 46826 480134
rect 47062 479898 47146 480134
rect 47382 479898 262826 480134
rect 263062 479898 263146 480134
rect 263382 479898 298826 480134
rect 299062 479898 299146 480134
rect 299382 479898 334826 480134
rect 335062 479898 335146 480134
rect 335382 479898 370826 480134
rect 371062 479898 371146 480134
rect 371382 479898 406826 480134
rect 407062 479898 407146 480134
rect 407382 479898 442826 480134
rect 443062 479898 443146 480134
rect 443382 479898 478826 480134
rect 479062 479898 479146 480134
rect 479382 479898 514826 480134
rect 515062 479898 515146 480134
rect 515382 479898 550826 480134
rect 551062 479898 551146 480134
rect 551382 479898 587262 480134
rect 587498 479898 587582 480134
rect 587818 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 475954 592650 475986
rect -8726 475718 -2934 475954
rect -2698 475718 -2614 475954
rect -2378 475718 6326 475954
rect 6562 475718 6646 475954
rect 6882 475718 42326 475954
rect 42562 475718 42646 475954
rect 42882 475718 71610 475954
rect 71846 475718 102330 475954
rect 102566 475718 133050 475954
rect 133286 475718 163770 475954
rect 164006 475718 194490 475954
rect 194726 475718 225210 475954
rect 225446 475718 258326 475954
rect 258562 475718 258646 475954
rect 258882 475718 294326 475954
rect 294562 475718 294646 475954
rect 294882 475718 330326 475954
rect 330562 475718 330646 475954
rect 330882 475718 366326 475954
rect 366562 475718 366646 475954
rect 366882 475718 402326 475954
rect 402562 475718 402646 475954
rect 402882 475718 438326 475954
rect 438562 475718 438646 475954
rect 438882 475718 474326 475954
rect 474562 475718 474646 475954
rect 474882 475718 510326 475954
rect 510562 475718 510646 475954
rect 510882 475718 546326 475954
rect 546562 475718 546646 475954
rect 546882 475718 582326 475954
rect 582562 475718 582646 475954
rect 582882 475718 586302 475954
rect 586538 475718 586622 475954
rect 586858 475718 592650 475954
rect -8726 475634 592650 475718
rect -8726 475398 -2934 475634
rect -2698 475398 -2614 475634
rect -2378 475398 6326 475634
rect 6562 475398 6646 475634
rect 6882 475398 42326 475634
rect 42562 475398 42646 475634
rect 42882 475398 71610 475634
rect 71846 475398 102330 475634
rect 102566 475398 133050 475634
rect 133286 475398 163770 475634
rect 164006 475398 194490 475634
rect 194726 475398 225210 475634
rect 225446 475398 258326 475634
rect 258562 475398 258646 475634
rect 258882 475398 294326 475634
rect 294562 475398 294646 475634
rect 294882 475398 330326 475634
rect 330562 475398 330646 475634
rect 330882 475398 366326 475634
rect 366562 475398 366646 475634
rect 366882 475398 402326 475634
rect 402562 475398 402646 475634
rect 402882 475398 438326 475634
rect 438562 475398 438646 475634
rect 438882 475398 474326 475634
rect 474562 475398 474646 475634
rect 474882 475398 510326 475634
rect 510562 475398 510646 475634
rect 510882 475398 546326 475634
rect 546562 475398 546646 475634
rect 546882 475398 582326 475634
rect 582562 475398 582646 475634
rect 582882 475398 586302 475634
rect 586538 475398 586622 475634
rect 586858 475398 592650 475634
rect -8726 475366 592650 475398
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 56250 471454
rect 56486 471218 86970 471454
rect 87206 471218 117690 471454
rect 117926 471218 148410 471454
rect 148646 471218 179130 471454
rect 179366 471218 209850 471454
rect 210086 471218 240570 471454
rect 240806 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 56250 471134
rect 56486 470898 86970 471134
rect 87206 470898 117690 471134
rect 117926 470898 148410 471134
rect 148646 470898 179130 471134
rect 179366 470898 209850 471134
rect 210086 470898 240570 471134
rect 240806 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 466954 592650 466986
rect -8726 466718 -8694 466954
rect -8458 466718 -8374 466954
rect -8138 466718 33326 466954
rect 33562 466718 33646 466954
rect 33882 466718 285326 466954
rect 285562 466718 285646 466954
rect 285882 466718 321326 466954
rect 321562 466718 321646 466954
rect 321882 466718 357326 466954
rect 357562 466718 357646 466954
rect 357882 466718 393326 466954
rect 393562 466718 393646 466954
rect 393882 466718 429326 466954
rect 429562 466718 429646 466954
rect 429882 466718 465326 466954
rect 465562 466718 465646 466954
rect 465882 466718 501326 466954
rect 501562 466718 501646 466954
rect 501882 466718 537326 466954
rect 537562 466718 537646 466954
rect 537882 466718 573326 466954
rect 573562 466718 573646 466954
rect 573882 466718 592062 466954
rect 592298 466718 592382 466954
rect 592618 466718 592650 466954
rect -8726 466634 592650 466718
rect -8726 466398 -8694 466634
rect -8458 466398 -8374 466634
rect -8138 466398 33326 466634
rect 33562 466398 33646 466634
rect 33882 466398 285326 466634
rect 285562 466398 285646 466634
rect 285882 466398 321326 466634
rect 321562 466398 321646 466634
rect 321882 466398 357326 466634
rect 357562 466398 357646 466634
rect 357882 466398 393326 466634
rect 393562 466398 393646 466634
rect 393882 466398 429326 466634
rect 429562 466398 429646 466634
rect 429882 466398 465326 466634
rect 465562 466398 465646 466634
rect 465882 466398 501326 466634
rect 501562 466398 501646 466634
rect 501882 466398 537326 466634
rect 537562 466398 537646 466634
rect 537882 466398 573326 466634
rect 573562 466398 573646 466634
rect 573882 466398 592062 466634
rect 592298 466398 592382 466634
rect 592618 466398 592650 466634
rect -8726 466366 592650 466398
rect -8726 462454 592650 462486
rect -8726 462218 -7734 462454
rect -7498 462218 -7414 462454
rect -7178 462218 28826 462454
rect 29062 462218 29146 462454
rect 29382 462218 280826 462454
rect 281062 462218 281146 462454
rect 281382 462218 316826 462454
rect 317062 462218 317146 462454
rect 317382 462218 352826 462454
rect 353062 462218 353146 462454
rect 353382 462218 388826 462454
rect 389062 462218 389146 462454
rect 389382 462218 424826 462454
rect 425062 462218 425146 462454
rect 425382 462218 460826 462454
rect 461062 462218 461146 462454
rect 461382 462218 496826 462454
rect 497062 462218 497146 462454
rect 497382 462218 532826 462454
rect 533062 462218 533146 462454
rect 533382 462218 568826 462454
rect 569062 462218 569146 462454
rect 569382 462218 591102 462454
rect 591338 462218 591422 462454
rect 591658 462218 592650 462454
rect -8726 462134 592650 462218
rect -8726 461898 -7734 462134
rect -7498 461898 -7414 462134
rect -7178 461898 28826 462134
rect 29062 461898 29146 462134
rect 29382 461898 280826 462134
rect 281062 461898 281146 462134
rect 281382 461898 316826 462134
rect 317062 461898 317146 462134
rect 317382 461898 352826 462134
rect 353062 461898 353146 462134
rect 353382 461898 388826 462134
rect 389062 461898 389146 462134
rect 389382 461898 424826 462134
rect 425062 461898 425146 462134
rect 425382 461898 460826 462134
rect 461062 461898 461146 462134
rect 461382 461898 496826 462134
rect 497062 461898 497146 462134
rect 497382 461898 532826 462134
rect 533062 461898 533146 462134
rect 533382 461898 568826 462134
rect 569062 461898 569146 462134
rect 569382 461898 591102 462134
rect 591338 461898 591422 462134
rect 591658 461898 592650 462134
rect -8726 461866 592650 461898
rect -8726 457954 592650 457986
rect -8726 457718 -6774 457954
rect -6538 457718 -6454 457954
rect -6218 457718 24326 457954
rect 24562 457718 24646 457954
rect 24882 457718 276326 457954
rect 276562 457718 276646 457954
rect 276882 457718 312326 457954
rect 312562 457718 312646 457954
rect 312882 457718 348326 457954
rect 348562 457718 348646 457954
rect 348882 457718 384326 457954
rect 384562 457718 384646 457954
rect 384882 457718 420326 457954
rect 420562 457718 420646 457954
rect 420882 457718 456326 457954
rect 456562 457718 456646 457954
rect 456882 457718 492326 457954
rect 492562 457718 492646 457954
rect 492882 457718 528326 457954
rect 528562 457718 528646 457954
rect 528882 457718 564326 457954
rect 564562 457718 564646 457954
rect 564882 457718 590142 457954
rect 590378 457718 590462 457954
rect 590698 457718 592650 457954
rect -8726 457634 592650 457718
rect -8726 457398 -6774 457634
rect -6538 457398 -6454 457634
rect -6218 457398 24326 457634
rect 24562 457398 24646 457634
rect 24882 457398 276326 457634
rect 276562 457398 276646 457634
rect 276882 457398 312326 457634
rect 312562 457398 312646 457634
rect 312882 457398 348326 457634
rect 348562 457398 348646 457634
rect 348882 457398 384326 457634
rect 384562 457398 384646 457634
rect 384882 457398 420326 457634
rect 420562 457398 420646 457634
rect 420882 457398 456326 457634
rect 456562 457398 456646 457634
rect 456882 457398 492326 457634
rect 492562 457398 492646 457634
rect 492882 457398 528326 457634
rect 528562 457398 528646 457634
rect 528882 457398 564326 457634
rect 564562 457398 564646 457634
rect 564882 457398 590142 457634
rect 590378 457398 590462 457634
rect 590698 457398 592650 457634
rect -8726 457366 592650 457398
rect -8726 453454 592650 453486
rect -8726 453218 -5814 453454
rect -5578 453218 -5494 453454
rect -5258 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 589182 453454
rect 589418 453218 589502 453454
rect 589738 453218 592650 453454
rect -8726 453134 592650 453218
rect -8726 452898 -5814 453134
rect -5578 452898 -5494 453134
rect -5258 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 589182 453134
rect 589418 452898 589502 453134
rect 589738 452898 592650 453134
rect -8726 452866 592650 452898
rect -8726 448954 592650 448986
rect -8726 448718 -4854 448954
rect -4618 448718 -4534 448954
rect -4298 448718 15326 448954
rect 15562 448718 15646 448954
rect 15882 448718 267326 448954
rect 267562 448718 267646 448954
rect 267882 448718 303326 448954
rect 303562 448718 303646 448954
rect 303882 448718 339326 448954
rect 339562 448718 339646 448954
rect 339882 448718 375326 448954
rect 375562 448718 375646 448954
rect 375882 448718 411326 448954
rect 411562 448718 411646 448954
rect 411882 448718 447326 448954
rect 447562 448718 447646 448954
rect 447882 448718 483326 448954
rect 483562 448718 483646 448954
rect 483882 448718 519326 448954
rect 519562 448718 519646 448954
rect 519882 448718 555326 448954
rect 555562 448718 555646 448954
rect 555882 448718 588222 448954
rect 588458 448718 588542 448954
rect 588778 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -4854 448634
rect -4618 448398 -4534 448634
rect -4298 448398 15326 448634
rect 15562 448398 15646 448634
rect 15882 448398 267326 448634
rect 267562 448398 267646 448634
rect 267882 448398 303326 448634
rect 303562 448398 303646 448634
rect 303882 448398 339326 448634
rect 339562 448398 339646 448634
rect 339882 448398 375326 448634
rect 375562 448398 375646 448634
rect 375882 448398 411326 448634
rect 411562 448398 411646 448634
rect 411882 448398 447326 448634
rect 447562 448398 447646 448634
rect 447882 448398 483326 448634
rect 483562 448398 483646 448634
rect 483882 448398 519326 448634
rect 519562 448398 519646 448634
rect 519882 448398 555326 448634
rect 555562 448398 555646 448634
rect 555882 448398 588222 448634
rect 588458 448398 588542 448634
rect 588778 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -3894 444454
rect -3658 444218 -3574 444454
rect -3338 444218 10826 444454
rect 11062 444218 11146 444454
rect 11382 444218 46826 444454
rect 47062 444218 47146 444454
rect 47382 444218 262826 444454
rect 263062 444218 263146 444454
rect 263382 444218 298826 444454
rect 299062 444218 299146 444454
rect 299382 444218 334826 444454
rect 335062 444218 335146 444454
rect 335382 444218 370826 444454
rect 371062 444218 371146 444454
rect 371382 444218 406826 444454
rect 407062 444218 407146 444454
rect 407382 444218 442826 444454
rect 443062 444218 443146 444454
rect 443382 444218 478826 444454
rect 479062 444218 479146 444454
rect 479382 444218 514826 444454
rect 515062 444218 515146 444454
rect 515382 444218 550826 444454
rect 551062 444218 551146 444454
rect 551382 444218 587262 444454
rect 587498 444218 587582 444454
rect 587818 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -3894 444134
rect -3658 443898 -3574 444134
rect -3338 443898 10826 444134
rect 11062 443898 11146 444134
rect 11382 443898 46826 444134
rect 47062 443898 47146 444134
rect 47382 443898 262826 444134
rect 263062 443898 263146 444134
rect 263382 443898 298826 444134
rect 299062 443898 299146 444134
rect 299382 443898 334826 444134
rect 335062 443898 335146 444134
rect 335382 443898 370826 444134
rect 371062 443898 371146 444134
rect 371382 443898 406826 444134
rect 407062 443898 407146 444134
rect 407382 443898 442826 444134
rect 443062 443898 443146 444134
rect 443382 443898 478826 444134
rect 479062 443898 479146 444134
rect 479382 443898 514826 444134
rect 515062 443898 515146 444134
rect 515382 443898 550826 444134
rect 551062 443898 551146 444134
rect 551382 443898 587262 444134
rect 587498 443898 587582 444134
rect 587818 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 439954 592650 439986
rect -8726 439718 -2934 439954
rect -2698 439718 -2614 439954
rect -2378 439718 6326 439954
rect 6562 439718 6646 439954
rect 6882 439718 42326 439954
rect 42562 439718 42646 439954
rect 42882 439718 71610 439954
rect 71846 439718 102330 439954
rect 102566 439718 133050 439954
rect 133286 439718 163770 439954
rect 164006 439718 194490 439954
rect 194726 439718 225210 439954
rect 225446 439718 258326 439954
rect 258562 439718 258646 439954
rect 258882 439718 294326 439954
rect 294562 439718 294646 439954
rect 294882 439718 330326 439954
rect 330562 439718 330646 439954
rect 330882 439718 366326 439954
rect 366562 439718 366646 439954
rect 366882 439718 402326 439954
rect 402562 439718 402646 439954
rect 402882 439718 438326 439954
rect 438562 439718 438646 439954
rect 438882 439718 474326 439954
rect 474562 439718 474646 439954
rect 474882 439718 510326 439954
rect 510562 439718 510646 439954
rect 510882 439718 546326 439954
rect 546562 439718 546646 439954
rect 546882 439718 582326 439954
rect 582562 439718 582646 439954
rect 582882 439718 586302 439954
rect 586538 439718 586622 439954
rect 586858 439718 592650 439954
rect -8726 439634 592650 439718
rect -8726 439398 -2934 439634
rect -2698 439398 -2614 439634
rect -2378 439398 6326 439634
rect 6562 439398 6646 439634
rect 6882 439398 42326 439634
rect 42562 439398 42646 439634
rect 42882 439398 71610 439634
rect 71846 439398 102330 439634
rect 102566 439398 133050 439634
rect 133286 439398 163770 439634
rect 164006 439398 194490 439634
rect 194726 439398 225210 439634
rect 225446 439398 258326 439634
rect 258562 439398 258646 439634
rect 258882 439398 294326 439634
rect 294562 439398 294646 439634
rect 294882 439398 330326 439634
rect 330562 439398 330646 439634
rect 330882 439398 366326 439634
rect 366562 439398 366646 439634
rect 366882 439398 402326 439634
rect 402562 439398 402646 439634
rect 402882 439398 438326 439634
rect 438562 439398 438646 439634
rect 438882 439398 474326 439634
rect 474562 439398 474646 439634
rect 474882 439398 510326 439634
rect 510562 439398 510646 439634
rect 510882 439398 546326 439634
rect 546562 439398 546646 439634
rect 546882 439398 582326 439634
rect 582562 439398 582646 439634
rect 582882 439398 586302 439634
rect 586538 439398 586622 439634
rect 586858 439398 592650 439634
rect -8726 439366 592650 439398
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 56250 435454
rect 56486 435218 86970 435454
rect 87206 435218 117690 435454
rect 117926 435218 148410 435454
rect 148646 435218 179130 435454
rect 179366 435218 209850 435454
rect 210086 435218 240570 435454
rect 240806 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 56250 435134
rect 56486 434898 86970 435134
rect 87206 434898 117690 435134
rect 117926 434898 148410 435134
rect 148646 434898 179130 435134
rect 179366 434898 209850 435134
rect 210086 434898 240570 435134
rect 240806 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 430954 592650 430986
rect -8726 430718 -8694 430954
rect -8458 430718 -8374 430954
rect -8138 430718 33326 430954
rect 33562 430718 33646 430954
rect 33882 430718 285326 430954
rect 285562 430718 285646 430954
rect 285882 430718 321326 430954
rect 321562 430718 321646 430954
rect 321882 430718 357326 430954
rect 357562 430718 357646 430954
rect 357882 430718 393326 430954
rect 393562 430718 393646 430954
rect 393882 430718 429326 430954
rect 429562 430718 429646 430954
rect 429882 430718 465326 430954
rect 465562 430718 465646 430954
rect 465882 430718 501326 430954
rect 501562 430718 501646 430954
rect 501882 430718 537326 430954
rect 537562 430718 537646 430954
rect 537882 430718 573326 430954
rect 573562 430718 573646 430954
rect 573882 430718 592062 430954
rect 592298 430718 592382 430954
rect 592618 430718 592650 430954
rect -8726 430634 592650 430718
rect -8726 430398 -8694 430634
rect -8458 430398 -8374 430634
rect -8138 430398 33326 430634
rect 33562 430398 33646 430634
rect 33882 430398 285326 430634
rect 285562 430398 285646 430634
rect 285882 430398 321326 430634
rect 321562 430398 321646 430634
rect 321882 430398 357326 430634
rect 357562 430398 357646 430634
rect 357882 430398 393326 430634
rect 393562 430398 393646 430634
rect 393882 430398 429326 430634
rect 429562 430398 429646 430634
rect 429882 430398 465326 430634
rect 465562 430398 465646 430634
rect 465882 430398 501326 430634
rect 501562 430398 501646 430634
rect 501882 430398 537326 430634
rect 537562 430398 537646 430634
rect 537882 430398 573326 430634
rect 573562 430398 573646 430634
rect 573882 430398 592062 430634
rect 592298 430398 592382 430634
rect 592618 430398 592650 430634
rect -8726 430366 592650 430398
rect -8726 426454 592650 426486
rect -8726 426218 -7734 426454
rect -7498 426218 -7414 426454
rect -7178 426218 28826 426454
rect 29062 426218 29146 426454
rect 29382 426218 280826 426454
rect 281062 426218 281146 426454
rect 281382 426218 316826 426454
rect 317062 426218 317146 426454
rect 317382 426218 352826 426454
rect 353062 426218 353146 426454
rect 353382 426218 388826 426454
rect 389062 426218 389146 426454
rect 389382 426218 424826 426454
rect 425062 426218 425146 426454
rect 425382 426218 460826 426454
rect 461062 426218 461146 426454
rect 461382 426218 496826 426454
rect 497062 426218 497146 426454
rect 497382 426218 532826 426454
rect 533062 426218 533146 426454
rect 533382 426218 568826 426454
rect 569062 426218 569146 426454
rect 569382 426218 591102 426454
rect 591338 426218 591422 426454
rect 591658 426218 592650 426454
rect -8726 426134 592650 426218
rect -8726 425898 -7734 426134
rect -7498 425898 -7414 426134
rect -7178 425898 28826 426134
rect 29062 425898 29146 426134
rect 29382 425898 280826 426134
rect 281062 425898 281146 426134
rect 281382 425898 316826 426134
rect 317062 425898 317146 426134
rect 317382 425898 352826 426134
rect 353062 425898 353146 426134
rect 353382 425898 388826 426134
rect 389062 425898 389146 426134
rect 389382 425898 424826 426134
rect 425062 425898 425146 426134
rect 425382 425898 460826 426134
rect 461062 425898 461146 426134
rect 461382 425898 496826 426134
rect 497062 425898 497146 426134
rect 497382 425898 532826 426134
rect 533062 425898 533146 426134
rect 533382 425898 568826 426134
rect 569062 425898 569146 426134
rect 569382 425898 591102 426134
rect 591338 425898 591422 426134
rect 591658 425898 592650 426134
rect -8726 425866 592650 425898
rect -8726 421954 592650 421986
rect -8726 421718 -6774 421954
rect -6538 421718 -6454 421954
rect -6218 421718 24326 421954
rect 24562 421718 24646 421954
rect 24882 421718 276326 421954
rect 276562 421718 276646 421954
rect 276882 421718 312326 421954
rect 312562 421718 312646 421954
rect 312882 421718 348326 421954
rect 348562 421718 348646 421954
rect 348882 421718 384326 421954
rect 384562 421718 384646 421954
rect 384882 421718 420326 421954
rect 420562 421718 420646 421954
rect 420882 421718 456326 421954
rect 456562 421718 456646 421954
rect 456882 421718 492326 421954
rect 492562 421718 492646 421954
rect 492882 421718 528326 421954
rect 528562 421718 528646 421954
rect 528882 421718 564326 421954
rect 564562 421718 564646 421954
rect 564882 421718 590142 421954
rect 590378 421718 590462 421954
rect 590698 421718 592650 421954
rect -8726 421634 592650 421718
rect -8726 421398 -6774 421634
rect -6538 421398 -6454 421634
rect -6218 421398 24326 421634
rect 24562 421398 24646 421634
rect 24882 421398 276326 421634
rect 276562 421398 276646 421634
rect 276882 421398 312326 421634
rect 312562 421398 312646 421634
rect 312882 421398 348326 421634
rect 348562 421398 348646 421634
rect 348882 421398 384326 421634
rect 384562 421398 384646 421634
rect 384882 421398 420326 421634
rect 420562 421398 420646 421634
rect 420882 421398 456326 421634
rect 456562 421398 456646 421634
rect 456882 421398 492326 421634
rect 492562 421398 492646 421634
rect 492882 421398 528326 421634
rect 528562 421398 528646 421634
rect 528882 421398 564326 421634
rect 564562 421398 564646 421634
rect 564882 421398 590142 421634
rect 590378 421398 590462 421634
rect 590698 421398 592650 421634
rect -8726 421366 592650 421398
rect -8726 417454 592650 417486
rect -8726 417218 -5814 417454
rect -5578 417218 -5494 417454
rect -5258 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 589182 417454
rect 589418 417218 589502 417454
rect 589738 417218 592650 417454
rect -8726 417134 592650 417218
rect -8726 416898 -5814 417134
rect -5578 416898 -5494 417134
rect -5258 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 589182 417134
rect 589418 416898 589502 417134
rect 589738 416898 592650 417134
rect -8726 416866 592650 416898
rect -8726 412954 592650 412986
rect -8726 412718 -4854 412954
rect -4618 412718 -4534 412954
rect -4298 412718 15326 412954
rect 15562 412718 15646 412954
rect 15882 412718 267326 412954
rect 267562 412718 267646 412954
rect 267882 412718 303326 412954
rect 303562 412718 303646 412954
rect 303882 412718 339326 412954
rect 339562 412718 339646 412954
rect 339882 412718 375326 412954
rect 375562 412718 375646 412954
rect 375882 412718 411326 412954
rect 411562 412718 411646 412954
rect 411882 412718 447326 412954
rect 447562 412718 447646 412954
rect 447882 412718 483326 412954
rect 483562 412718 483646 412954
rect 483882 412718 519326 412954
rect 519562 412718 519646 412954
rect 519882 412718 555326 412954
rect 555562 412718 555646 412954
rect 555882 412718 588222 412954
rect 588458 412718 588542 412954
rect 588778 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -4854 412634
rect -4618 412398 -4534 412634
rect -4298 412398 15326 412634
rect 15562 412398 15646 412634
rect 15882 412398 267326 412634
rect 267562 412398 267646 412634
rect 267882 412398 303326 412634
rect 303562 412398 303646 412634
rect 303882 412398 339326 412634
rect 339562 412398 339646 412634
rect 339882 412398 375326 412634
rect 375562 412398 375646 412634
rect 375882 412398 411326 412634
rect 411562 412398 411646 412634
rect 411882 412398 447326 412634
rect 447562 412398 447646 412634
rect 447882 412398 483326 412634
rect 483562 412398 483646 412634
rect 483882 412398 519326 412634
rect 519562 412398 519646 412634
rect 519882 412398 555326 412634
rect 555562 412398 555646 412634
rect 555882 412398 588222 412634
rect 588458 412398 588542 412634
rect 588778 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -3894 408454
rect -3658 408218 -3574 408454
rect -3338 408218 10826 408454
rect 11062 408218 11146 408454
rect 11382 408218 46826 408454
rect 47062 408218 47146 408454
rect 47382 408218 262826 408454
rect 263062 408218 263146 408454
rect 263382 408218 298826 408454
rect 299062 408218 299146 408454
rect 299382 408218 334826 408454
rect 335062 408218 335146 408454
rect 335382 408218 370826 408454
rect 371062 408218 371146 408454
rect 371382 408218 406826 408454
rect 407062 408218 407146 408454
rect 407382 408218 442826 408454
rect 443062 408218 443146 408454
rect 443382 408218 478826 408454
rect 479062 408218 479146 408454
rect 479382 408218 514826 408454
rect 515062 408218 515146 408454
rect 515382 408218 550826 408454
rect 551062 408218 551146 408454
rect 551382 408218 587262 408454
rect 587498 408218 587582 408454
rect 587818 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -3894 408134
rect -3658 407898 -3574 408134
rect -3338 407898 10826 408134
rect 11062 407898 11146 408134
rect 11382 407898 46826 408134
rect 47062 407898 47146 408134
rect 47382 407898 262826 408134
rect 263062 407898 263146 408134
rect 263382 407898 298826 408134
rect 299062 407898 299146 408134
rect 299382 407898 334826 408134
rect 335062 407898 335146 408134
rect 335382 407898 370826 408134
rect 371062 407898 371146 408134
rect 371382 407898 406826 408134
rect 407062 407898 407146 408134
rect 407382 407898 442826 408134
rect 443062 407898 443146 408134
rect 443382 407898 478826 408134
rect 479062 407898 479146 408134
rect 479382 407898 514826 408134
rect 515062 407898 515146 408134
rect 515382 407898 550826 408134
rect 551062 407898 551146 408134
rect 551382 407898 587262 408134
rect 587498 407898 587582 408134
rect 587818 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 403954 592650 403986
rect -8726 403718 -2934 403954
rect -2698 403718 -2614 403954
rect -2378 403718 6326 403954
rect 6562 403718 6646 403954
rect 6882 403718 42326 403954
rect 42562 403718 42646 403954
rect 42882 403718 71610 403954
rect 71846 403718 102330 403954
rect 102566 403718 133050 403954
rect 133286 403718 163770 403954
rect 164006 403718 194490 403954
rect 194726 403718 225210 403954
rect 225446 403718 258326 403954
rect 258562 403718 258646 403954
rect 258882 403718 294326 403954
rect 294562 403718 294646 403954
rect 294882 403718 330326 403954
rect 330562 403718 330646 403954
rect 330882 403718 366326 403954
rect 366562 403718 366646 403954
rect 366882 403718 402326 403954
rect 402562 403718 402646 403954
rect 402882 403718 438326 403954
rect 438562 403718 438646 403954
rect 438882 403718 474326 403954
rect 474562 403718 474646 403954
rect 474882 403718 510326 403954
rect 510562 403718 510646 403954
rect 510882 403718 546326 403954
rect 546562 403718 546646 403954
rect 546882 403718 582326 403954
rect 582562 403718 582646 403954
rect 582882 403718 586302 403954
rect 586538 403718 586622 403954
rect 586858 403718 592650 403954
rect -8726 403634 592650 403718
rect -8726 403398 -2934 403634
rect -2698 403398 -2614 403634
rect -2378 403398 6326 403634
rect 6562 403398 6646 403634
rect 6882 403398 42326 403634
rect 42562 403398 42646 403634
rect 42882 403398 71610 403634
rect 71846 403398 102330 403634
rect 102566 403398 133050 403634
rect 133286 403398 163770 403634
rect 164006 403398 194490 403634
rect 194726 403398 225210 403634
rect 225446 403398 258326 403634
rect 258562 403398 258646 403634
rect 258882 403398 294326 403634
rect 294562 403398 294646 403634
rect 294882 403398 330326 403634
rect 330562 403398 330646 403634
rect 330882 403398 366326 403634
rect 366562 403398 366646 403634
rect 366882 403398 402326 403634
rect 402562 403398 402646 403634
rect 402882 403398 438326 403634
rect 438562 403398 438646 403634
rect 438882 403398 474326 403634
rect 474562 403398 474646 403634
rect 474882 403398 510326 403634
rect 510562 403398 510646 403634
rect 510882 403398 546326 403634
rect 546562 403398 546646 403634
rect 546882 403398 582326 403634
rect 582562 403398 582646 403634
rect 582882 403398 586302 403634
rect 586538 403398 586622 403634
rect 586858 403398 592650 403634
rect -8726 403366 592650 403398
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 56250 399454
rect 56486 399218 86970 399454
rect 87206 399218 117690 399454
rect 117926 399218 148410 399454
rect 148646 399218 179130 399454
rect 179366 399218 209850 399454
rect 210086 399218 240570 399454
rect 240806 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 56250 399134
rect 56486 398898 86970 399134
rect 87206 398898 117690 399134
rect 117926 398898 148410 399134
rect 148646 398898 179130 399134
rect 179366 398898 209850 399134
rect 210086 398898 240570 399134
rect 240806 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 394954 592650 394986
rect -8726 394718 -8694 394954
rect -8458 394718 -8374 394954
rect -8138 394718 33326 394954
rect 33562 394718 33646 394954
rect 33882 394718 285326 394954
rect 285562 394718 285646 394954
rect 285882 394718 321326 394954
rect 321562 394718 321646 394954
rect 321882 394718 357326 394954
rect 357562 394718 357646 394954
rect 357882 394718 393326 394954
rect 393562 394718 393646 394954
rect 393882 394718 429326 394954
rect 429562 394718 429646 394954
rect 429882 394718 465326 394954
rect 465562 394718 465646 394954
rect 465882 394718 501326 394954
rect 501562 394718 501646 394954
rect 501882 394718 537326 394954
rect 537562 394718 537646 394954
rect 537882 394718 573326 394954
rect 573562 394718 573646 394954
rect 573882 394718 592062 394954
rect 592298 394718 592382 394954
rect 592618 394718 592650 394954
rect -8726 394634 592650 394718
rect -8726 394398 -8694 394634
rect -8458 394398 -8374 394634
rect -8138 394398 33326 394634
rect 33562 394398 33646 394634
rect 33882 394398 285326 394634
rect 285562 394398 285646 394634
rect 285882 394398 321326 394634
rect 321562 394398 321646 394634
rect 321882 394398 357326 394634
rect 357562 394398 357646 394634
rect 357882 394398 393326 394634
rect 393562 394398 393646 394634
rect 393882 394398 429326 394634
rect 429562 394398 429646 394634
rect 429882 394398 465326 394634
rect 465562 394398 465646 394634
rect 465882 394398 501326 394634
rect 501562 394398 501646 394634
rect 501882 394398 537326 394634
rect 537562 394398 537646 394634
rect 537882 394398 573326 394634
rect 573562 394398 573646 394634
rect 573882 394398 592062 394634
rect 592298 394398 592382 394634
rect 592618 394398 592650 394634
rect -8726 394366 592650 394398
rect -8726 390454 592650 390486
rect -8726 390218 -7734 390454
rect -7498 390218 -7414 390454
rect -7178 390218 28826 390454
rect 29062 390218 29146 390454
rect 29382 390218 280826 390454
rect 281062 390218 281146 390454
rect 281382 390218 316826 390454
rect 317062 390218 317146 390454
rect 317382 390218 352826 390454
rect 353062 390218 353146 390454
rect 353382 390218 388826 390454
rect 389062 390218 389146 390454
rect 389382 390218 424826 390454
rect 425062 390218 425146 390454
rect 425382 390218 460826 390454
rect 461062 390218 461146 390454
rect 461382 390218 496826 390454
rect 497062 390218 497146 390454
rect 497382 390218 532826 390454
rect 533062 390218 533146 390454
rect 533382 390218 568826 390454
rect 569062 390218 569146 390454
rect 569382 390218 591102 390454
rect 591338 390218 591422 390454
rect 591658 390218 592650 390454
rect -8726 390134 592650 390218
rect -8726 389898 -7734 390134
rect -7498 389898 -7414 390134
rect -7178 389898 28826 390134
rect 29062 389898 29146 390134
rect 29382 389898 280826 390134
rect 281062 389898 281146 390134
rect 281382 389898 316826 390134
rect 317062 389898 317146 390134
rect 317382 389898 352826 390134
rect 353062 389898 353146 390134
rect 353382 389898 388826 390134
rect 389062 389898 389146 390134
rect 389382 389898 424826 390134
rect 425062 389898 425146 390134
rect 425382 389898 460826 390134
rect 461062 389898 461146 390134
rect 461382 389898 496826 390134
rect 497062 389898 497146 390134
rect 497382 389898 532826 390134
rect 533062 389898 533146 390134
rect 533382 389898 568826 390134
rect 569062 389898 569146 390134
rect 569382 389898 591102 390134
rect 591338 389898 591422 390134
rect 591658 389898 592650 390134
rect -8726 389866 592650 389898
rect -8726 385954 592650 385986
rect -8726 385718 -6774 385954
rect -6538 385718 -6454 385954
rect -6218 385718 24326 385954
rect 24562 385718 24646 385954
rect 24882 385718 276326 385954
rect 276562 385718 276646 385954
rect 276882 385718 312326 385954
rect 312562 385718 312646 385954
rect 312882 385718 348326 385954
rect 348562 385718 348646 385954
rect 348882 385718 384326 385954
rect 384562 385718 384646 385954
rect 384882 385718 420326 385954
rect 420562 385718 420646 385954
rect 420882 385718 456326 385954
rect 456562 385718 456646 385954
rect 456882 385718 492326 385954
rect 492562 385718 492646 385954
rect 492882 385718 528326 385954
rect 528562 385718 528646 385954
rect 528882 385718 564326 385954
rect 564562 385718 564646 385954
rect 564882 385718 590142 385954
rect 590378 385718 590462 385954
rect 590698 385718 592650 385954
rect -8726 385634 592650 385718
rect -8726 385398 -6774 385634
rect -6538 385398 -6454 385634
rect -6218 385398 24326 385634
rect 24562 385398 24646 385634
rect 24882 385398 276326 385634
rect 276562 385398 276646 385634
rect 276882 385398 312326 385634
rect 312562 385398 312646 385634
rect 312882 385398 348326 385634
rect 348562 385398 348646 385634
rect 348882 385398 384326 385634
rect 384562 385398 384646 385634
rect 384882 385398 420326 385634
rect 420562 385398 420646 385634
rect 420882 385398 456326 385634
rect 456562 385398 456646 385634
rect 456882 385398 492326 385634
rect 492562 385398 492646 385634
rect 492882 385398 528326 385634
rect 528562 385398 528646 385634
rect 528882 385398 564326 385634
rect 564562 385398 564646 385634
rect 564882 385398 590142 385634
rect 590378 385398 590462 385634
rect 590698 385398 592650 385634
rect -8726 385366 592650 385398
rect -8726 381454 592650 381486
rect -8726 381218 -5814 381454
rect -5578 381218 -5494 381454
rect -5258 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 589182 381454
rect 589418 381218 589502 381454
rect 589738 381218 592650 381454
rect -8726 381134 592650 381218
rect -8726 380898 -5814 381134
rect -5578 380898 -5494 381134
rect -5258 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 589182 381134
rect 589418 380898 589502 381134
rect 589738 380898 592650 381134
rect -8726 380866 592650 380898
rect -8726 376954 592650 376986
rect -8726 376718 -4854 376954
rect -4618 376718 -4534 376954
rect -4298 376718 15326 376954
rect 15562 376718 15646 376954
rect 15882 376718 267326 376954
rect 267562 376718 267646 376954
rect 267882 376718 303326 376954
rect 303562 376718 303646 376954
rect 303882 376718 339326 376954
rect 339562 376718 339646 376954
rect 339882 376718 375326 376954
rect 375562 376718 375646 376954
rect 375882 376718 411326 376954
rect 411562 376718 411646 376954
rect 411882 376718 447326 376954
rect 447562 376718 447646 376954
rect 447882 376718 483326 376954
rect 483562 376718 483646 376954
rect 483882 376718 519326 376954
rect 519562 376718 519646 376954
rect 519882 376718 555326 376954
rect 555562 376718 555646 376954
rect 555882 376718 588222 376954
rect 588458 376718 588542 376954
rect 588778 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -4854 376634
rect -4618 376398 -4534 376634
rect -4298 376398 15326 376634
rect 15562 376398 15646 376634
rect 15882 376398 267326 376634
rect 267562 376398 267646 376634
rect 267882 376398 303326 376634
rect 303562 376398 303646 376634
rect 303882 376398 339326 376634
rect 339562 376398 339646 376634
rect 339882 376398 375326 376634
rect 375562 376398 375646 376634
rect 375882 376398 411326 376634
rect 411562 376398 411646 376634
rect 411882 376398 447326 376634
rect 447562 376398 447646 376634
rect 447882 376398 483326 376634
rect 483562 376398 483646 376634
rect 483882 376398 519326 376634
rect 519562 376398 519646 376634
rect 519882 376398 555326 376634
rect 555562 376398 555646 376634
rect 555882 376398 588222 376634
rect 588458 376398 588542 376634
rect 588778 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -3894 372454
rect -3658 372218 -3574 372454
rect -3338 372218 10826 372454
rect 11062 372218 11146 372454
rect 11382 372218 46826 372454
rect 47062 372218 47146 372454
rect 47382 372218 262826 372454
rect 263062 372218 263146 372454
rect 263382 372218 298826 372454
rect 299062 372218 299146 372454
rect 299382 372218 334826 372454
rect 335062 372218 335146 372454
rect 335382 372218 370826 372454
rect 371062 372218 371146 372454
rect 371382 372218 406826 372454
rect 407062 372218 407146 372454
rect 407382 372218 442826 372454
rect 443062 372218 443146 372454
rect 443382 372218 478826 372454
rect 479062 372218 479146 372454
rect 479382 372218 514826 372454
rect 515062 372218 515146 372454
rect 515382 372218 550826 372454
rect 551062 372218 551146 372454
rect 551382 372218 587262 372454
rect 587498 372218 587582 372454
rect 587818 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -3894 372134
rect -3658 371898 -3574 372134
rect -3338 371898 10826 372134
rect 11062 371898 11146 372134
rect 11382 371898 46826 372134
rect 47062 371898 47146 372134
rect 47382 371898 262826 372134
rect 263062 371898 263146 372134
rect 263382 371898 298826 372134
rect 299062 371898 299146 372134
rect 299382 371898 334826 372134
rect 335062 371898 335146 372134
rect 335382 371898 370826 372134
rect 371062 371898 371146 372134
rect 371382 371898 406826 372134
rect 407062 371898 407146 372134
rect 407382 371898 442826 372134
rect 443062 371898 443146 372134
rect 443382 371898 478826 372134
rect 479062 371898 479146 372134
rect 479382 371898 514826 372134
rect 515062 371898 515146 372134
rect 515382 371898 550826 372134
rect 551062 371898 551146 372134
rect 551382 371898 587262 372134
rect 587498 371898 587582 372134
rect 587818 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 367954 592650 367986
rect -8726 367718 -2934 367954
rect -2698 367718 -2614 367954
rect -2378 367718 6326 367954
rect 6562 367718 6646 367954
rect 6882 367718 42326 367954
rect 42562 367718 42646 367954
rect 42882 367718 71610 367954
rect 71846 367718 102330 367954
rect 102566 367718 133050 367954
rect 133286 367718 163770 367954
rect 164006 367718 194490 367954
rect 194726 367718 225210 367954
rect 225446 367718 258326 367954
rect 258562 367718 258646 367954
rect 258882 367718 294326 367954
rect 294562 367718 294646 367954
rect 294882 367718 330326 367954
rect 330562 367718 330646 367954
rect 330882 367718 366326 367954
rect 366562 367718 366646 367954
rect 366882 367718 402326 367954
rect 402562 367718 402646 367954
rect 402882 367718 438326 367954
rect 438562 367718 438646 367954
rect 438882 367718 474326 367954
rect 474562 367718 474646 367954
rect 474882 367718 510326 367954
rect 510562 367718 510646 367954
rect 510882 367718 546326 367954
rect 546562 367718 546646 367954
rect 546882 367718 582326 367954
rect 582562 367718 582646 367954
rect 582882 367718 586302 367954
rect 586538 367718 586622 367954
rect 586858 367718 592650 367954
rect -8726 367634 592650 367718
rect -8726 367398 -2934 367634
rect -2698 367398 -2614 367634
rect -2378 367398 6326 367634
rect 6562 367398 6646 367634
rect 6882 367398 42326 367634
rect 42562 367398 42646 367634
rect 42882 367398 71610 367634
rect 71846 367398 102330 367634
rect 102566 367398 133050 367634
rect 133286 367398 163770 367634
rect 164006 367398 194490 367634
rect 194726 367398 225210 367634
rect 225446 367398 258326 367634
rect 258562 367398 258646 367634
rect 258882 367398 294326 367634
rect 294562 367398 294646 367634
rect 294882 367398 330326 367634
rect 330562 367398 330646 367634
rect 330882 367398 366326 367634
rect 366562 367398 366646 367634
rect 366882 367398 402326 367634
rect 402562 367398 402646 367634
rect 402882 367398 438326 367634
rect 438562 367398 438646 367634
rect 438882 367398 474326 367634
rect 474562 367398 474646 367634
rect 474882 367398 510326 367634
rect 510562 367398 510646 367634
rect 510882 367398 546326 367634
rect 546562 367398 546646 367634
rect 546882 367398 582326 367634
rect 582562 367398 582646 367634
rect 582882 367398 586302 367634
rect 586538 367398 586622 367634
rect 586858 367398 592650 367634
rect -8726 367366 592650 367398
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 56250 363454
rect 56486 363218 86970 363454
rect 87206 363218 117690 363454
rect 117926 363218 148410 363454
rect 148646 363218 179130 363454
rect 179366 363218 209850 363454
rect 210086 363218 240570 363454
rect 240806 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 56250 363134
rect 56486 362898 86970 363134
rect 87206 362898 117690 363134
rect 117926 362898 148410 363134
rect 148646 362898 179130 363134
rect 179366 362898 209850 363134
rect 210086 362898 240570 363134
rect 240806 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 358954 592650 358986
rect -8726 358718 -8694 358954
rect -8458 358718 -8374 358954
rect -8138 358718 33326 358954
rect 33562 358718 33646 358954
rect 33882 358718 285326 358954
rect 285562 358718 285646 358954
rect 285882 358718 321326 358954
rect 321562 358718 321646 358954
rect 321882 358718 357326 358954
rect 357562 358718 357646 358954
rect 357882 358718 393326 358954
rect 393562 358718 393646 358954
rect 393882 358718 429326 358954
rect 429562 358718 429646 358954
rect 429882 358718 465326 358954
rect 465562 358718 465646 358954
rect 465882 358718 501326 358954
rect 501562 358718 501646 358954
rect 501882 358718 537326 358954
rect 537562 358718 537646 358954
rect 537882 358718 573326 358954
rect 573562 358718 573646 358954
rect 573882 358718 592062 358954
rect 592298 358718 592382 358954
rect 592618 358718 592650 358954
rect -8726 358634 592650 358718
rect -8726 358398 -8694 358634
rect -8458 358398 -8374 358634
rect -8138 358398 33326 358634
rect 33562 358398 33646 358634
rect 33882 358398 285326 358634
rect 285562 358398 285646 358634
rect 285882 358398 321326 358634
rect 321562 358398 321646 358634
rect 321882 358398 357326 358634
rect 357562 358398 357646 358634
rect 357882 358398 393326 358634
rect 393562 358398 393646 358634
rect 393882 358398 429326 358634
rect 429562 358398 429646 358634
rect 429882 358398 465326 358634
rect 465562 358398 465646 358634
rect 465882 358398 501326 358634
rect 501562 358398 501646 358634
rect 501882 358398 537326 358634
rect 537562 358398 537646 358634
rect 537882 358398 573326 358634
rect 573562 358398 573646 358634
rect 573882 358398 592062 358634
rect 592298 358398 592382 358634
rect 592618 358398 592650 358634
rect -8726 358366 592650 358398
rect -8726 354454 592650 354486
rect -8726 354218 -7734 354454
rect -7498 354218 -7414 354454
rect -7178 354218 28826 354454
rect 29062 354218 29146 354454
rect 29382 354218 280826 354454
rect 281062 354218 281146 354454
rect 281382 354218 316826 354454
rect 317062 354218 317146 354454
rect 317382 354218 352826 354454
rect 353062 354218 353146 354454
rect 353382 354218 388826 354454
rect 389062 354218 389146 354454
rect 389382 354218 424826 354454
rect 425062 354218 425146 354454
rect 425382 354218 460826 354454
rect 461062 354218 461146 354454
rect 461382 354218 496826 354454
rect 497062 354218 497146 354454
rect 497382 354218 532826 354454
rect 533062 354218 533146 354454
rect 533382 354218 568826 354454
rect 569062 354218 569146 354454
rect 569382 354218 591102 354454
rect 591338 354218 591422 354454
rect 591658 354218 592650 354454
rect -8726 354134 592650 354218
rect -8726 353898 -7734 354134
rect -7498 353898 -7414 354134
rect -7178 353898 28826 354134
rect 29062 353898 29146 354134
rect 29382 353898 280826 354134
rect 281062 353898 281146 354134
rect 281382 353898 316826 354134
rect 317062 353898 317146 354134
rect 317382 353898 352826 354134
rect 353062 353898 353146 354134
rect 353382 353898 388826 354134
rect 389062 353898 389146 354134
rect 389382 353898 424826 354134
rect 425062 353898 425146 354134
rect 425382 353898 460826 354134
rect 461062 353898 461146 354134
rect 461382 353898 496826 354134
rect 497062 353898 497146 354134
rect 497382 353898 532826 354134
rect 533062 353898 533146 354134
rect 533382 353898 568826 354134
rect 569062 353898 569146 354134
rect 569382 353898 591102 354134
rect 591338 353898 591422 354134
rect 591658 353898 592650 354134
rect -8726 353866 592650 353898
rect -8726 349954 592650 349986
rect -8726 349718 -6774 349954
rect -6538 349718 -6454 349954
rect -6218 349718 24326 349954
rect 24562 349718 24646 349954
rect 24882 349718 276326 349954
rect 276562 349718 276646 349954
rect 276882 349718 312326 349954
rect 312562 349718 312646 349954
rect 312882 349718 348326 349954
rect 348562 349718 348646 349954
rect 348882 349718 384326 349954
rect 384562 349718 384646 349954
rect 384882 349718 420326 349954
rect 420562 349718 420646 349954
rect 420882 349718 456326 349954
rect 456562 349718 456646 349954
rect 456882 349718 492326 349954
rect 492562 349718 492646 349954
rect 492882 349718 528326 349954
rect 528562 349718 528646 349954
rect 528882 349718 564326 349954
rect 564562 349718 564646 349954
rect 564882 349718 590142 349954
rect 590378 349718 590462 349954
rect 590698 349718 592650 349954
rect -8726 349634 592650 349718
rect -8726 349398 -6774 349634
rect -6538 349398 -6454 349634
rect -6218 349398 24326 349634
rect 24562 349398 24646 349634
rect 24882 349398 276326 349634
rect 276562 349398 276646 349634
rect 276882 349398 312326 349634
rect 312562 349398 312646 349634
rect 312882 349398 348326 349634
rect 348562 349398 348646 349634
rect 348882 349398 384326 349634
rect 384562 349398 384646 349634
rect 384882 349398 420326 349634
rect 420562 349398 420646 349634
rect 420882 349398 456326 349634
rect 456562 349398 456646 349634
rect 456882 349398 492326 349634
rect 492562 349398 492646 349634
rect 492882 349398 528326 349634
rect 528562 349398 528646 349634
rect 528882 349398 564326 349634
rect 564562 349398 564646 349634
rect 564882 349398 590142 349634
rect 590378 349398 590462 349634
rect 590698 349398 592650 349634
rect -8726 349366 592650 349398
rect -8726 345454 592650 345486
rect -8726 345218 -5814 345454
rect -5578 345218 -5494 345454
rect -5258 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 589182 345454
rect 589418 345218 589502 345454
rect 589738 345218 592650 345454
rect -8726 345134 592650 345218
rect -8726 344898 -5814 345134
rect -5578 344898 -5494 345134
rect -5258 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 589182 345134
rect 589418 344898 589502 345134
rect 589738 344898 592650 345134
rect -8726 344866 592650 344898
rect -8726 340954 592650 340986
rect -8726 340718 -4854 340954
rect -4618 340718 -4534 340954
rect -4298 340718 15326 340954
rect 15562 340718 15646 340954
rect 15882 340718 267326 340954
rect 267562 340718 267646 340954
rect 267882 340718 303326 340954
rect 303562 340718 303646 340954
rect 303882 340718 339326 340954
rect 339562 340718 339646 340954
rect 339882 340718 375326 340954
rect 375562 340718 375646 340954
rect 375882 340718 411326 340954
rect 411562 340718 411646 340954
rect 411882 340718 447326 340954
rect 447562 340718 447646 340954
rect 447882 340718 483326 340954
rect 483562 340718 483646 340954
rect 483882 340718 519326 340954
rect 519562 340718 519646 340954
rect 519882 340718 555326 340954
rect 555562 340718 555646 340954
rect 555882 340718 588222 340954
rect 588458 340718 588542 340954
rect 588778 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -4854 340634
rect -4618 340398 -4534 340634
rect -4298 340398 15326 340634
rect 15562 340398 15646 340634
rect 15882 340398 267326 340634
rect 267562 340398 267646 340634
rect 267882 340398 303326 340634
rect 303562 340398 303646 340634
rect 303882 340398 339326 340634
rect 339562 340398 339646 340634
rect 339882 340398 375326 340634
rect 375562 340398 375646 340634
rect 375882 340398 411326 340634
rect 411562 340398 411646 340634
rect 411882 340398 447326 340634
rect 447562 340398 447646 340634
rect 447882 340398 483326 340634
rect 483562 340398 483646 340634
rect 483882 340398 519326 340634
rect 519562 340398 519646 340634
rect 519882 340398 555326 340634
rect 555562 340398 555646 340634
rect 555882 340398 588222 340634
rect 588458 340398 588542 340634
rect 588778 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -3894 336454
rect -3658 336218 -3574 336454
rect -3338 336218 10826 336454
rect 11062 336218 11146 336454
rect 11382 336218 46826 336454
rect 47062 336218 47146 336454
rect 47382 336218 262826 336454
rect 263062 336218 263146 336454
rect 263382 336218 298826 336454
rect 299062 336218 299146 336454
rect 299382 336218 334826 336454
rect 335062 336218 335146 336454
rect 335382 336218 370826 336454
rect 371062 336218 371146 336454
rect 371382 336218 406826 336454
rect 407062 336218 407146 336454
rect 407382 336218 442826 336454
rect 443062 336218 443146 336454
rect 443382 336218 478826 336454
rect 479062 336218 479146 336454
rect 479382 336218 514826 336454
rect 515062 336218 515146 336454
rect 515382 336218 550826 336454
rect 551062 336218 551146 336454
rect 551382 336218 587262 336454
rect 587498 336218 587582 336454
rect 587818 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -3894 336134
rect -3658 335898 -3574 336134
rect -3338 335898 10826 336134
rect 11062 335898 11146 336134
rect 11382 335898 46826 336134
rect 47062 335898 47146 336134
rect 47382 335898 262826 336134
rect 263062 335898 263146 336134
rect 263382 335898 298826 336134
rect 299062 335898 299146 336134
rect 299382 335898 334826 336134
rect 335062 335898 335146 336134
rect 335382 335898 370826 336134
rect 371062 335898 371146 336134
rect 371382 335898 406826 336134
rect 407062 335898 407146 336134
rect 407382 335898 442826 336134
rect 443062 335898 443146 336134
rect 443382 335898 478826 336134
rect 479062 335898 479146 336134
rect 479382 335898 514826 336134
rect 515062 335898 515146 336134
rect 515382 335898 550826 336134
rect 551062 335898 551146 336134
rect 551382 335898 587262 336134
rect 587498 335898 587582 336134
rect 587818 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 331954 592650 331986
rect -8726 331718 -2934 331954
rect -2698 331718 -2614 331954
rect -2378 331718 6326 331954
rect 6562 331718 6646 331954
rect 6882 331718 42326 331954
rect 42562 331718 42646 331954
rect 42882 331718 71610 331954
rect 71846 331718 102330 331954
rect 102566 331718 133050 331954
rect 133286 331718 163770 331954
rect 164006 331718 194490 331954
rect 194726 331718 225210 331954
rect 225446 331718 258326 331954
rect 258562 331718 258646 331954
rect 258882 331718 294326 331954
rect 294562 331718 294646 331954
rect 294882 331718 366326 331954
rect 366562 331718 366646 331954
rect 366882 331718 402326 331954
rect 402562 331718 402646 331954
rect 402882 331718 438326 331954
rect 438562 331718 438646 331954
rect 438882 331718 474326 331954
rect 474562 331718 474646 331954
rect 474882 331718 510326 331954
rect 510562 331718 510646 331954
rect 510882 331718 546326 331954
rect 546562 331718 546646 331954
rect 546882 331718 582326 331954
rect 582562 331718 582646 331954
rect 582882 331718 586302 331954
rect 586538 331718 586622 331954
rect 586858 331718 592650 331954
rect -8726 331634 592650 331718
rect -8726 331398 -2934 331634
rect -2698 331398 -2614 331634
rect -2378 331398 6326 331634
rect 6562 331398 6646 331634
rect 6882 331398 42326 331634
rect 42562 331398 42646 331634
rect 42882 331398 71610 331634
rect 71846 331398 102330 331634
rect 102566 331398 133050 331634
rect 133286 331398 163770 331634
rect 164006 331398 194490 331634
rect 194726 331398 225210 331634
rect 225446 331398 258326 331634
rect 258562 331398 258646 331634
rect 258882 331398 294326 331634
rect 294562 331398 294646 331634
rect 294882 331398 366326 331634
rect 366562 331398 366646 331634
rect 366882 331398 402326 331634
rect 402562 331398 402646 331634
rect 402882 331398 438326 331634
rect 438562 331398 438646 331634
rect 438882 331398 474326 331634
rect 474562 331398 474646 331634
rect 474882 331398 510326 331634
rect 510562 331398 510646 331634
rect 510882 331398 546326 331634
rect 546562 331398 546646 331634
rect 546882 331398 582326 331634
rect 582562 331398 582646 331634
rect 582882 331398 586302 331634
rect 586538 331398 586622 331634
rect 586858 331398 592650 331634
rect -8726 331366 592650 331398
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 56250 327454
rect 56486 327218 86970 327454
rect 87206 327218 117690 327454
rect 117926 327218 148410 327454
rect 148646 327218 179130 327454
rect 179366 327218 209850 327454
rect 210086 327218 240570 327454
rect 240806 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327239 361826 327454
rect 290382 327218 304250 327239
rect -8726 327134 304250 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 56250 327134
rect 56486 326898 86970 327134
rect 87206 326898 117690 327134
rect 117926 326898 148410 327134
rect 148646 326898 179130 327134
rect 179366 326898 209850 327134
rect 210086 326898 240570 327134
rect 240806 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 327003 304250 327134
rect 304486 327003 334970 327239
rect 335206 327218 361826 327239
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect 335206 327134 592650 327218
rect 335206 327003 361826 327134
rect 290382 326898 361826 327003
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 322954 592650 322986
rect -8726 322718 -8694 322954
rect -8458 322718 -8374 322954
rect -8138 322718 33326 322954
rect 33562 322718 33646 322954
rect 33882 322718 285326 322954
rect 285562 322718 285646 322954
rect 285882 322718 357326 322954
rect 357562 322718 357646 322954
rect 357882 322718 393326 322954
rect 393562 322718 393646 322954
rect 393882 322718 429326 322954
rect 429562 322718 429646 322954
rect 429882 322718 465326 322954
rect 465562 322718 465646 322954
rect 465882 322718 501326 322954
rect 501562 322718 501646 322954
rect 501882 322718 537326 322954
rect 537562 322718 537646 322954
rect 537882 322718 573326 322954
rect 573562 322718 573646 322954
rect 573882 322718 592062 322954
rect 592298 322718 592382 322954
rect 592618 322718 592650 322954
rect -8726 322634 592650 322718
rect -8726 322398 -8694 322634
rect -8458 322398 -8374 322634
rect -8138 322398 33326 322634
rect 33562 322398 33646 322634
rect 33882 322398 285326 322634
rect 285562 322398 285646 322634
rect 285882 322398 357326 322634
rect 357562 322398 357646 322634
rect 357882 322398 393326 322634
rect 393562 322398 393646 322634
rect 393882 322398 429326 322634
rect 429562 322398 429646 322634
rect 429882 322398 465326 322634
rect 465562 322398 465646 322634
rect 465882 322398 501326 322634
rect 501562 322398 501646 322634
rect 501882 322398 537326 322634
rect 537562 322398 537646 322634
rect 537882 322398 573326 322634
rect 573562 322398 573646 322634
rect 573882 322398 592062 322634
rect 592298 322398 592382 322634
rect 592618 322398 592650 322634
rect -8726 322366 592650 322398
rect -8726 318454 592650 318486
rect -8726 318218 -7734 318454
rect -7498 318218 -7414 318454
rect -7178 318218 28826 318454
rect 29062 318218 29146 318454
rect 29382 318218 280826 318454
rect 281062 318218 281146 318454
rect 281382 318218 388826 318454
rect 389062 318218 389146 318454
rect 389382 318218 424826 318454
rect 425062 318218 425146 318454
rect 425382 318218 460826 318454
rect 461062 318218 461146 318454
rect 461382 318218 496826 318454
rect 497062 318218 497146 318454
rect 497382 318218 532826 318454
rect 533062 318218 533146 318454
rect 533382 318218 568826 318454
rect 569062 318218 569146 318454
rect 569382 318218 591102 318454
rect 591338 318218 591422 318454
rect 591658 318218 592650 318454
rect -8726 318134 592650 318218
rect -8726 317898 -7734 318134
rect -7498 317898 -7414 318134
rect -7178 317898 28826 318134
rect 29062 317898 29146 318134
rect 29382 317898 280826 318134
rect 281062 317898 281146 318134
rect 281382 317898 388826 318134
rect 389062 317898 389146 318134
rect 389382 317898 424826 318134
rect 425062 317898 425146 318134
rect 425382 317898 460826 318134
rect 461062 317898 461146 318134
rect 461382 317898 496826 318134
rect 497062 317898 497146 318134
rect 497382 317898 532826 318134
rect 533062 317898 533146 318134
rect 533382 317898 568826 318134
rect 569062 317898 569146 318134
rect 569382 317898 591102 318134
rect 591338 317898 591422 318134
rect 591658 317898 592650 318134
rect -8726 317866 592650 317898
rect -8726 313954 592650 313986
rect -8726 313718 -6774 313954
rect -6538 313718 -6454 313954
rect -6218 313718 24326 313954
rect 24562 313718 24646 313954
rect 24882 313718 276326 313954
rect 276562 313718 276646 313954
rect 276882 313718 384326 313954
rect 384562 313718 384646 313954
rect 384882 313718 420326 313954
rect 420562 313718 420646 313954
rect 420882 313718 456326 313954
rect 456562 313718 456646 313954
rect 456882 313718 492326 313954
rect 492562 313718 492646 313954
rect 492882 313718 528326 313954
rect 528562 313718 528646 313954
rect 528882 313718 564326 313954
rect 564562 313718 564646 313954
rect 564882 313718 590142 313954
rect 590378 313718 590462 313954
rect 590698 313718 592650 313954
rect -8726 313634 592650 313718
rect -8726 313398 -6774 313634
rect -6538 313398 -6454 313634
rect -6218 313398 24326 313634
rect 24562 313398 24646 313634
rect 24882 313398 276326 313634
rect 276562 313398 276646 313634
rect 276882 313398 384326 313634
rect 384562 313398 384646 313634
rect 384882 313398 420326 313634
rect 420562 313398 420646 313634
rect 420882 313398 456326 313634
rect 456562 313398 456646 313634
rect 456882 313398 492326 313634
rect 492562 313398 492646 313634
rect 492882 313398 528326 313634
rect 528562 313398 528646 313634
rect 528882 313398 564326 313634
rect 564562 313398 564646 313634
rect 564882 313398 590142 313634
rect 590378 313398 590462 313634
rect 590698 313398 592650 313634
rect -8726 313366 592650 313398
rect -8726 309454 592650 309486
rect -8726 309218 -5814 309454
rect -5578 309218 -5494 309454
rect -5258 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 589182 309454
rect 589418 309218 589502 309454
rect 589738 309218 592650 309454
rect -8726 309134 592650 309218
rect -8726 308898 -5814 309134
rect -5578 308898 -5494 309134
rect -5258 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 589182 309134
rect 589418 308898 589502 309134
rect 589738 308898 592650 309134
rect -8726 308866 592650 308898
rect -8726 304954 592650 304986
rect -8726 304718 -4854 304954
rect -4618 304718 -4534 304954
rect -4298 304718 15326 304954
rect 15562 304718 15646 304954
rect 15882 304718 267326 304954
rect 267562 304718 267646 304954
rect 267882 304718 375326 304954
rect 375562 304718 375646 304954
rect 375882 304718 411326 304954
rect 411562 304718 411646 304954
rect 411882 304718 447326 304954
rect 447562 304718 447646 304954
rect 447882 304718 483326 304954
rect 483562 304718 483646 304954
rect 483882 304718 519326 304954
rect 519562 304718 519646 304954
rect 519882 304718 555326 304954
rect 555562 304718 555646 304954
rect 555882 304718 588222 304954
rect 588458 304718 588542 304954
rect 588778 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -4854 304634
rect -4618 304398 -4534 304634
rect -4298 304398 15326 304634
rect 15562 304398 15646 304634
rect 15882 304398 267326 304634
rect 267562 304398 267646 304634
rect 267882 304398 375326 304634
rect 375562 304398 375646 304634
rect 375882 304398 411326 304634
rect 411562 304398 411646 304634
rect 411882 304398 447326 304634
rect 447562 304398 447646 304634
rect 447882 304398 483326 304634
rect 483562 304398 483646 304634
rect 483882 304398 519326 304634
rect 519562 304398 519646 304634
rect 519882 304398 555326 304634
rect 555562 304398 555646 304634
rect 555882 304398 588222 304634
rect 588458 304398 588542 304634
rect 588778 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -3894 300454
rect -3658 300218 -3574 300454
rect -3338 300218 10826 300454
rect 11062 300218 11146 300454
rect 11382 300218 46826 300454
rect 47062 300218 47146 300454
rect 47382 300218 262826 300454
rect 263062 300218 263146 300454
rect 263382 300218 370826 300454
rect 371062 300218 371146 300454
rect 371382 300218 406826 300454
rect 407062 300218 407146 300454
rect 407382 300218 442826 300454
rect 443062 300218 443146 300454
rect 443382 300218 478826 300454
rect 479062 300218 479146 300454
rect 479382 300218 514826 300454
rect 515062 300218 515146 300454
rect 515382 300218 550826 300454
rect 551062 300218 551146 300454
rect 551382 300218 587262 300454
rect 587498 300218 587582 300454
rect 587818 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -3894 300134
rect -3658 299898 -3574 300134
rect -3338 299898 10826 300134
rect 11062 299898 11146 300134
rect 11382 299898 46826 300134
rect 47062 299898 47146 300134
rect 47382 299898 262826 300134
rect 263062 299898 263146 300134
rect 263382 299898 370826 300134
rect 371062 299898 371146 300134
rect 371382 299898 406826 300134
rect 407062 299898 407146 300134
rect 407382 299898 442826 300134
rect 443062 299898 443146 300134
rect 443382 299898 478826 300134
rect 479062 299898 479146 300134
rect 479382 299898 514826 300134
rect 515062 299898 515146 300134
rect 515382 299898 550826 300134
rect 551062 299898 551146 300134
rect 551382 299898 587262 300134
rect 587498 299898 587582 300134
rect 587818 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 295954 592650 295986
rect -8726 295718 -2934 295954
rect -2698 295718 -2614 295954
rect -2378 295718 6326 295954
rect 6562 295718 6646 295954
rect 6882 295718 42326 295954
rect 42562 295718 42646 295954
rect 42882 295718 71610 295954
rect 71846 295718 102330 295954
rect 102566 295718 133050 295954
rect 133286 295718 163770 295954
rect 164006 295718 194490 295954
rect 194726 295718 225210 295954
rect 225446 295718 258326 295954
rect 258562 295718 258646 295954
rect 258882 295718 294326 295954
rect 294562 295718 294646 295954
rect 294882 295718 319610 295954
rect 319846 295718 366326 295954
rect 366562 295718 366646 295954
rect 366882 295718 402326 295954
rect 402562 295718 402646 295954
rect 402882 295718 438326 295954
rect 438562 295718 438646 295954
rect 438882 295718 474326 295954
rect 474562 295718 474646 295954
rect 474882 295718 510326 295954
rect 510562 295718 510646 295954
rect 510882 295718 546326 295954
rect 546562 295718 546646 295954
rect 546882 295718 582326 295954
rect 582562 295718 582646 295954
rect 582882 295718 586302 295954
rect 586538 295718 586622 295954
rect 586858 295718 592650 295954
rect -8726 295634 592650 295718
rect -8726 295398 -2934 295634
rect -2698 295398 -2614 295634
rect -2378 295398 6326 295634
rect 6562 295398 6646 295634
rect 6882 295398 42326 295634
rect 42562 295398 42646 295634
rect 42882 295398 71610 295634
rect 71846 295398 102330 295634
rect 102566 295398 133050 295634
rect 133286 295398 163770 295634
rect 164006 295398 194490 295634
rect 194726 295398 225210 295634
rect 225446 295398 258326 295634
rect 258562 295398 258646 295634
rect 258882 295398 294326 295634
rect 294562 295398 294646 295634
rect 294882 295398 319610 295634
rect 319846 295398 366326 295634
rect 366562 295398 366646 295634
rect 366882 295398 402326 295634
rect 402562 295398 402646 295634
rect 402882 295398 438326 295634
rect 438562 295398 438646 295634
rect 438882 295398 474326 295634
rect 474562 295398 474646 295634
rect 474882 295398 510326 295634
rect 510562 295398 510646 295634
rect 510882 295398 546326 295634
rect 546562 295398 546646 295634
rect 546882 295398 582326 295634
rect 582562 295398 582646 295634
rect 582882 295398 586302 295634
rect 586538 295398 586622 295634
rect 586858 295398 592650 295634
rect -8726 295366 592650 295398
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 56250 291454
rect 56486 291218 86970 291454
rect 87206 291218 117690 291454
rect 117926 291218 148410 291454
rect 148646 291218 179130 291454
rect 179366 291218 209850 291454
rect 210086 291218 240570 291454
rect 240806 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 304250 291454
rect 304486 291218 334970 291454
rect 335206 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 56250 291134
rect 56486 290898 86970 291134
rect 87206 290898 117690 291134
rect 117926 290898 148410 291134
rect 148646 290898 179130 291134
rect 179366 290898 209850 291134
rect 210086 290898 240570 291134
rect 240806 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 304250 291134
rect 304486 290898 334970 291134
rect 335206 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 286954 592650 286986
rect -8726 286718 -8694 286954
rect -8458 286718 -8374 286954
rect -8138 286718 33326 286954
rect 33562 286718 33646 286954
rect 33882 286718 285326 286954
rect 285562 286718 285646 286954
rect 285882 286718 357326 286954
rect 357562 286718 357646 286954
rect 357882 286718 393326 286954
rect 393562 286718 393646 286954
rect 393882 286718 429326 286954
rect 429562 286718 429646 286954
rect 429882 286718 465326 286954
rect 465562 286718 465646 286954
rect 465882 286718 501326 286954
rect 501562 286718 501646 286954
rect 501882 286718 537326 286954
rect 537562 286718 537646 286954
rect 537882 286718 573326 286954
rect 573562 286718 573646 286954
rect 573882 286718 592062 286954
rect 592298 286718 592382 286954
rect 592618 286718 592650 286954
rect -8726 286634 592650 286718
rect -8726 286398 -8694 286634
rect -8458 286398 -8374 286634
rect -8138 286398 33326 286634
rect 33562 286398 33646 286634
rect 33882 286398 285326 286634
rect 285562 286398 285646 286634
rect 285882 286398 357326 286634
rect 357562 286398 357646 286634
rect 357882 286398 393326 286634
rect 393562 286398 393646 286634
rect 393882 286398 429326 286634
rect 429562 286398 429646 286634
rect 429882 286398 465326 286634
rect 465562 286398 465646 286634
rect 465882 286398 501326 286634
rect 501562 286398 501646 286634
rect 501882 286398 537326 286634
rect 537562 286398 537646 286634
rect 537882 286398 573326 286634
rect 573562 286398 573646 286634
rect 573882 286398 592062 286634
rect 592298 286398 592382 286634
rect 592618 286398 592650 286634
rect -8726 286366 592650 286398
rect -8726 282454 592650 282486
rect -8726 282218 -7734 282454
rect -7498 282218 -7414 282454
rect -7178 282218 28826 282454
rect 29062 282218 29146 282454
rect 29382 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 388826 282454
rect 389062 282218 389146 282454
rect 389382 282218 424826 282454
rect 425062 282218 425146 282454
rect 425382 282218 460826 282454
rect 461062 282218 461146 282454
rect 461382 282218 496826 282454
rect 497062 282218 497146 282454
rect 497382 282218 532826 282454
rect 533062 282218 533146 282454
rect 533382 282218 568826 282454
rect 569062 282218 569146 282454
rect 569382 282218 591102 282454
rect 591338 282218 591422 282454
rect 591658 282218 592650 282454
rect -8726 282134 592650 282218
rect -8726 281898 -7734 282134
rect -7498 281898 -7414 282134
rect -7178 281898 28826 282134
rect 29062 281898 29146 282134
rect 29382 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 388826 282134
rect 389062 281898 389146 282134
rect 389382 281898 424826 282134
rect 425062 281898 425146 282134
rect 425382 281898 460826 282134
rect 461062 281898 461146 282134
rect 461382 281898 496826 282134
rect 497062 281898 497146 282134
rect 497382 281898 532826 282134
rect 533062 281898 533146 282134
rect 533382 281898 568826 282134
rect 569062 281898 569146 282134
rect 569382 281898 591102 282134
rect 591338 281898 591422 282134
rect 591658 281898 592650 282134
rect -8726 281866 592650 281898
rect -8726 277954 592650 277986
rect -8726 277718 -6774 277954
rect -6538 277718 -6454 277954
rect -6218 277718 24326 277954
rect 24562 277718 24646 277954
rect 24882 277718 60326 277954
rect 60562 277718 60646 277954
rect 60882 277718 96326 277954
rect 96562 277718 96646 277954
rect 96882 277718 132326 277954
rect 132562 277718 132646 277954
rect 132882 277718 168326 277954
rect 168562 277718 168646 277954
rect 168882 277718 204326 277954
rect 204562 277718 204646 277954
rect 204882 277718 240326 277954
rect 240562 277718 240646 277954
rect 240882 277718 276326 277954
rect 276562 277718 276646 277954
rect 276882 277718 312326 277954
rect 312562 277718 312646 277954
rect 312882 277718 348326 277954
rect 348562 277718 348646 277954
rect 348882 277718 384326 277954
rect 384562 277718 384646 277954
rect 384882 277718 420326 277954
rect 420562 277718 420646 277954
rect 420882 277718 456326 277954
rect 456562 277718 456646 277954
rect 456882 277718 492326 277954
rect 492562 277718 492646 277954
rect 492882 277718 528326 277954
rect 528562 277718 528646 277954
rect 528882 277718 564326 277954
rect 564562 277718 564646 277954
rect 564882 277718 590142 277954
rect 590378 277718 590462 277954
rect 590698 277718 592650 277954
rect -8726 277634 592650 277718
rect -8726 277398 -6774 277634
rect -6538 277398 -6454 277634
rect -6218 277398 24326 277634
rect 24562 277398 24646 277634
rect 24882 277398 60326 277634
rect 60562 277398 60646 277634
rect 60882 277398 96326 277634
rect 96562 277398 96646 277634
rect 96882 277398 132326 277634
rect 132562 277398 132646 277634
rect 132882 277398 168326 277634
rect 168562 277398 168646 277634
rect 168882 277398 204326 277634
rect 204562 277398 204646 277634
rect 204882 277398 240326 277634
rect 240562 277398 240646 277634
rect 240882 277398 276326 277634
rect 276562 277398 276646 277634
rect 276882 277398 312326 277634
rect 312562 277398 312646 277634
rect 312882 277398 348326 277634
rect 348562 277398 348646 277634
rect 348882 277398 384326 277634
rect 384562 277398 384646 277634
rect 384882 277398 420326 277634
rect 420562 277398 420646 277634
rect 420882 277398 456326 277634
rect 456562 277398 456646 277634
rect 456882 277398 492326 277634
rect 492562 277398 492646 277634
rect 492882 277398 528326 277634
rect 528562 277398 528646 277634
rect 528882 277398 564326 277634
rect 564562 277398 564646 277634
rect 564882 277398 590142 277634
rect 590378 277398 590462 277634
rect 590698 277398 592650 277634
rect -8726 277366 592650 277398
rect -8726 273454 592650 273486
rect -8726 273218 -5814 273454
rect -5578 273218 -5494 273454
rect -5258 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 589182 273454
rect 589418 273218 589502 273454
rect 589738 273218 592650 273454
rect -8726 273134 592650 273218
rect -8726 272898 -5814 273134
rect -5578 272898 -5494 273134
rect -5258 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 589182 273134
rect 589418 272898 589502 273134
rect 589738 272898 592650 273134
rect -8726 272866 592650 272898
rect -8726 268954 592650 268986
rect -8726 268718 -4854 268954
rect -4618 268718 -4534 268954
rect -4298 268718 15326 268954
rect 15562 268718 15646 268954
rect 15882 268718 51326 268954
rect 51562 268718 51646 268954
rect 51882 268718 87326 268954
rect 87562 268718 87646 268954
rect 87882 268718 123326 268954
rect 123562 268718 123646 268954
rect 123882 268718 159326 268954
rect 159562 268718 159646 268954
rect 159882 268718 195326 268954
rect 195562 268718 195646 268954
rect 195882 268718 231326 268954
rect 231562 268718 231646 268954
rect 231882 268718 267326 268954
rect 267562 268718 267646 268954
rect 267882 268718 303326 268954
rect 303562 268718 303646 268954
rect 303882 268718 339326 268954
rect 339562 268718 339646 268954
rect 339882 268718 375326 268954
rect 375562 268718 375646 268954
rect 375882 268718 411326 268954
rect 411562 268718 411646 268954
rect 411882 268718 447326 268954
rect 447562 268718 447646 268954
rect 447882 268718 483326 268954
rect 483562 268718 483646 268954
rect 483882 268718 519326 268954
rect 519562 268718 519646 268954
rect 519882 268718 555326 268954
rect 555562 268718 555646 268954
rect 555882 268718 588222 268954
rect 588458 268718 588542 268954
rect 588778 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -4854 268634
rect -4618 268398 -4534 268634
rect -4298 268398 15326 268634
rect 15562 268398 15646 268634
rect 15882 268398 51326 268634
rect 51562 268398 51646 268634
rect 51882 268398 87326 268634
rect 87562 268398 87646 268634
rect 87882 268398 123326 268634
rect 123562 268398 123646 268634
rect 123882 268398 159326 268634
rect 159562 268398 159646 268634
rect 159882 268398 195326 268634
rect 195562 268398 195646 268634
rect 195882 268398 231326 268634
rect 231562 268398 231646 268634
rect 231882 268398 267326 268634
rect 267562 268398 267646 268634
rect 267882 268398 303326 268634
rect 303562 268398 303646 268634
rect 303882 268398 339326 268634
rect 339562 268398 339646 268634
rect 339882 268398 375326 268634
rect 375562 268398 375646 268634
rect 375882 268398 411326 268634
rect 411562 268398 411646 268634
rect 411882 268398 447326 268634
rect 447562 268398 447646 268634
rect 447882 268398 483326 268634
rect 483562 268398 483646 268634
rect 483882 268398 519326 268634
rect 519562 268398 519646 268634
rect 519882 268398 555326 268634
rect 555562 268398 555646 268634
rect 555882 268398 588222 268634
rect 588458 268398 588542 268634
rect 588778 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -3894 264454
rect -3658 264218 -3574 264454
rect -3338 264218 10826 264454
rect 11062 264218 11146 264454
rect 11382 264218 46826 264454
rect 47062 264218 47146 264454
rect 47382 264218 82826 264454
rect 83062 264218 83146 264454
rect 83382 264218 118826 264454
rect 119062 264218 119146 264454
rect 119382 264218 154826 264454
rect 155062 264218 155146 264454
rect 155382 264218 190826 264454
rect 191062 264218 191146 264454
rect 191382 264218 226826 264454
rect 227062 264218 227146 264454
rect 227382 264218 262826 264454
rect 263062 264218 263146 264454
rect 263382 264218 298826 264454
rect 299062 264218 299146 264454
rect 299382 264218 334826 264454
rect 335062 264218 335146 264454
rect 335382 264218 370826 264454
rect 371062 264218 371146 264454
rect 371382 264218 406826 264454
rect 407062 264218 407146 264454
rect 407382 264218 442826 264454
rect 443062 264218 443146 264454
rect 443382 264218 478826 264454
rect 479062 264218 479146 264454
rect 479382 264218 514826 264454
rect 515062 264218 515146 264454
rect 515382 264218 550826 264454
rect 551062 264218 551146 264454
rect 551382 264218 587262 264454
rect 587498 264218 587582 264454
rect 587818 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -3894 264134
rect -3658 263898 -3574 264134
rect -3338 263898 10826 264134
rect 11062 263898 11146 264134
rect 11382 263898 46826 264134
rect 47062 263898 47146 264134
rect 47382 263898 82826 264134
rect 83062 263898 83146 264134
rect 83382 263898 118826 264134
rect 119062 263898 119146 264134
rect 119382 263898 154826 264134
rect 155062 263898 155146 264134
rect 155382 263898 190826 264134
rect 191062 263898 191146 264134
rect 191382 263898 226826 264134
rect 227062 263898 227146 264134
rect 227382 263898 262826 264134
rect 263062 263898 263146 264134
rect 263382 263898 298826 264134
rect 299062 263898 299146 264134
rect 299382 263898 334826 264134
rect 335062 263898 335146 264134
rect 335382 263898 370826 264134
rect 371062 263898 371146 264134
rect 371382 263898 406826 264134
rect 407062 263898 407146 264134
rect 407382 263898 442826 264134
rect 443062 263898 443146 264134
rect 443382 263898 478826 264134
rect 479062 263898 479146 264134
rect 479382 263898 514826 264134
rect 515062 263898 515146 264134
rect 515382 263898 550826 264134
rect 551062 263898 551146 264134
rect 551382 263898 587262 264134
rect 587498 263898 587582 264134
rect 587818 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 259954 592650 259986
rect -8726 259718 -2934 259954
rect -2698 259718 -2614 259954
rect -2378 259718 6326 259954
rect 6562 259718 6646 259954
rect 6882 259718 42326 259954
rect 42562 259718 42646 259954
rect 42882 259718 78326 259954
rect 78562 259718 78646 259954
rect 78882 259718 114326 259954
rect 114562 259718 114646 259954
rect 114882 259718 150326 259954
rect 150562 259718 150646 259954
rect 150882 259718 186326 259954
rect 186562 259718 186646 259954
rect 186882 259718 222326 259954
rect 222562 259718 222646 259954
rect 222882 259718 258326 259954
rect 258562 259718 258646 259954
rect 258882 259718 294326 259954
rect 294562 259718 294646 259954
rect 294882 259718 330326 259954
rect 330562 259718 330646 259954
rect 330882 259718 366326 259954
rect 366562 259718 366646 259954
rect 366882 259718 402326 259954
rect 402562 259718 402646 259954
rect 402882 259718 438326 259954
rect 438562 259718 438646 259954
rect 438882 259718 474326 259954
rect 474562 259718 474646 259954
rect 474882 259718 510326 259954
rect 510562 259718 510646 259954
rect 510882 259718 546326 259954
rect 546562 259718 546646 259954
rect 546882 259718 582326 259954
rect 582562 259718 582646 259954
rect 582882 259718 586302 259954
rect 586538 259718 586622 259954
rect 586858 259718 592650 259954
rect -8726 259634 592650 259718
rect -8726 259398 -2934 259634
rect -2698 259398 -2614 259634
rect -2378 259398 6326 259634
rect 6562 259398 6646 259634
rect 6882 259398 42326 259634
rect 42562 259398 42646 259634
rect 42882 259398 78326 259634
rect 78562 259398 78646 259634
rect 78882 259398 114326 259634
rect 114562 259398 114646 259634
rect 114882 259398 150326 259634
rect 150562 259398 150646 259634
rect 150882 259398 186326 259634
rect 186562 259398 186646 259634
rect 186882 259398 222326 259634
rect 222562 259398 222646 259634
rect 222882 259398 258326 259634
rect 258562 259398 258646 259634
rect 258882 259398 294326 259634
rect 294562 259398 294646 259634
rect 294882 259398 330326 259634
rect 330562 259398 330646 259634
rect 330882 259398 366326 259634
rect 366562 259398 366646 259634
rect 366882 259398 402326 259634
rect 402562 259398 402646 259634
rect 402882 259398 438326 259634
rect 438562 259398 438646 259634
rect 438882 259398 474326 259634
rect 474562 259398 474646 259634
rect 474882 259398 510326 259634
rect 510562 259398 510646 259634
rect 510882 259398 546326 259634
rect 546562 259398 546646 259634
rect 546882 259398 582326 259634
rect 582562 259398 582646 259634
rect 582882 259398 586302 259634
rect 586538 259398 586622 259634
rect 586858 259398 592650 259634
rect -8726 259366 592650 259398
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 250954 592650 250986
rect -8726 250718 -8694 250954
rect -8458 250718 -8374 250954
rect -8138 250718 33326 250954
rect 33562 250718 33646 250954
rect 33882 250718 249326 250954
rect 249562 250718 249646 250954
rect 249882 250718 285326 250954
rect 285562 250718 285646 250954
rect 285882 250718 357326 250954
rect 357562 250718 357646 250954
rect 357882 250718 393326 250954
rect 393562 250718 393646 250954
rect 393882 250718 429326 250954
rect 429562 250718 429646 250954
rect 429882 250718 465326 250954
rect 465562 250718 465646 250954
rect 465882 250718 501326 250954
rect 501562 250718 501646 250954
rect 501882 250718 537326 250954
rect 537562 250718 537646 250954
rect 537882 250718 573326 250954
rect 573562 250718 573646 250954
rect 573882 250718 592062 250954
rect 592298 250718 592382 250954
rect 592618 250718 592650 250954
rect -8726 250634 592650 250718
rect -8726 250398 -8694 250634
rect -8458 250398 -8374 250634
rect -8138 250398 33326 250634
rect 33562 250398 33646 250634
rect 33882 250398 249326 250634
rect 249562 250398 249646 250634
rect 249882 250398 285326 250634
rect 285562 250398 285646 250634
rect 285882 250398 357326 250634
rect 357562 250398 357646 250634
rect 357882 250398 393326 250634
rect 393562 250398 393646 250634
rect 393882 250398 429326 250634
rect 429562 250398 429646 250634
rect 429882 250398 465326 250634
rect 465562 250398 465646 250634
rect 465882 250398 501326 250634
rect 501562 250398 501646 250634
rect 501882 250398 537326 250634
rect 537562 250398 537646 250634
rect 537882 250398 573326 250634
rect 573562 250398 573646 250634
rect 573882 250398 592062 250634
rect 592298 250398 592382 250634
rect 592618 250398 592650 250634
rect -8726 250366 592650 250398
rect -8726 246454 592650 246486
rect -8726 246218 -7734 246454
rect -7498 246218 -7414 246454
rect -7178 246218 28826 246454
rect 29062 246218 29146 246454
rect 29382 246218 244826 246454
rect 245062 246218 245146 246454
rect 245382 246218 280826 246454
rect 281062 246218 281146 246454
rect 281382 246218 352826 246454
rect 353062 246218 353146 246454
rect 353382 246218 388826 246454
rect 389062 246218 389146 246454
rect 389382 246218 424826 246454
rect 425062 246218 425146 246454
rect 425382 246218 460826 246454
rect 461062 246218 461146 246454
rect 461382 246218 496826 246454
rect 497062 246218 497146 246454
rect 497382 246218 532826 246454
rect 533062 246218 533146 246454
rect 533382 246218 568826 246454
rect 569062 246218 569146 246454
rect 569382 246218 591102 246454
rect 591338 246218 591422 246454
rect 591658 246218 592650 246454
rect -8726 246134 592650 246218
rect -8726 245898 -7734 246134
rect -7498 245898 -7414 246134
rect -7178 245898 28826 246134
rect 29062 245898 29146 246134
rect 29382 245898 244826 246134
rect 245062 245898 245146 246134
rect 245382 245898 280826 246134
rect 281062 245898 281146 246134
rect 281382 245898 352826 246134
rect 353062 245898 353146 246134
rect 353382 245898 388826 246134
rect 389062 245898 389146 246134
rect 389382 245898 424826 246134
rect 425062 245898 425146 246134
rect 425382 245898 460826 246134
rect 461062 245898 461146 246134
rect 461382 245898 496826 246134
rect 497062 245898 497146 246134
rect 497382 245898 532826 246134
rect 533062 245898 533146 246134
rect 533382 245898 568826 246134
rect 569062 245898 569146 246134
rect 569382 245898 591102 246134
rect 591338 245898 591422 246134
rect 591658 245898 592650 246134
rect -8726 245866 592650 245898
rect -8726 241954 592650 241986
rect -8726 241718 -6774 241954
rect -6538 241718 -6454 241954
rect -6218 241718 24326 241954
rect 24562 241718 24646 241954
rect 24882 241718 60326 241954
rect 60562 241718 60646 241954
rect 60882 241718 96326 241954
rect 96562 241718 96646 241954
rect 96882 241718 132326 241954
rect 132562 241718 132646 241954
rect 132882 241718 168326 241954
rect 168562 241718 168646 241954
rect 168882 241718 204326 241954
rect 204562 241718 204646 241954
rect 204882 241718 240326 241954
rect 240562 241718 240646 241954
rect 240882 241718 276326 241954
rect 276562 241718 276646 241954
rect 276882 241718 312326 241954
rect 312562 241718 312646 241954
rect 312882 241718 348326 241954
rect 348562 241718 348646 241954
rect 348882 241718 384326 241954
rect 384562 241718 384646 241954
rect 384882 241718 420326 241954
rect 420562 241718 420646 241954
rect 420882 241718 456326 241954
rect 456562 241718 456646 241954
rect 456882 241718 492326 241954
rect 492562 241718 492646 241954
rect 492882 241718 528326 241954
rect 528562 241718 528646 241954
rect 528882 241718 564326 241954
rect 564562 241718 564646 241954
rect 564882 241718 590142 241954
rect 590378 241718 590462 241954
rect 590698 241718 592650 241954
rect -8726 241634 592650 241718
rect -8726 241398 -6774 241634
rect -6538 241398 -6454 241634
rect -6218 241398 24326 241634
rect 24562 241398 24646 241634
rect 24882 241398 60326 241634
rect 60562 241398 60646 241634
rect 60882 241398 96326 241634
rect 96562 241398 96646 241634
rect 96882 241398 132326 241634
rect 132562 241398 132646 241634
rect 132882 241398 168326 241634
rect 168562 241398 168646 241634
rect 168882 241398 204326 241634
rect 204562 241398 204646 241634
rect 204882 241398 240326 241634
rect 240562 241398 240646 241634
rect 240882 241398 276326 241634
rect 276562 241398 276646 241634
rect 276882 241398 312326 241634
rect 312562 241398 312646 241634
rect 312882 241398 348326 241634
rect 348562 241398 348646 241634
rect 348882 241398 384326 241634
rect 384562 241398 384646 241634
rect 384882 241398 420326 241634
rect 420562 241398 420646 241634
rect 420882 241398 456326 241634
rect 456562 241398 456646 241634
rect 456882 241398 492326 241634
rect 492562 241398 492646 241634
rect 492882 241398 528326 241634
rect 528562 241398 528646 241634
rect 528882 241398 564326 241634
rect 564562 241398 564646 241634
rect 564882 241398 590142 241634
rect 590378 241398 590462 241634
rect 590698 241398 592650 241634
rect -8726 241366 592650 241398
rect -8726 237454 592650 237486
rect -8726 237218 -5814 237454
rect -5578 237218 -5494 237454
rect -5258 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 589182 237454
rect 589418 237218 589502 237454
rect 589738 237218 592650 237454
rect -8726 237134 592650 237218
rect -8726 236898 -5814 237134
rect -5578 236898 -5494 237134
rect -5258 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 589182 237134
rect 589418 236898 589502 237134
rect 589738 236898 592650 237134
rect -8726 236866 592650 236898
rect -8726 232954 592650 232986
rect -8726 232718 -4854 232954
rect -4618 232718 -4534 232954
rect -4298 232718 15326 232954
rect 15562 232718 15646 232954
rect 15882 232718 51326 232954
rect 51562 232718 51646 232954
rect 51882 232718 87326 232954
rect 87562 232718 87646 232954
rect 87882 232718 123326 232954
rect 123562 232718 123646 232954
rect 123882 232718 159326 232954
rect 159562 232718 159646 232954
rect 159882 232718 195326 232954
rect 195562 232718 195646 232954
rect 195882 232718 231326 232954
rect 231562 232718 231646 232954
rect 231882 232718 267326 232954
rect 267562 232718 267646 232954
rect 267882 232718 303326 232954
rect 303562 232718 303646 232954
rect 303882 232718 339326 232954
rect 339562 232718 339646 232954
rect 339882 232718 375326 232954
rect 375562 232718 375646 232954
rect 375882 232718 411326 232954
rect 411562 232718 411646 232954
rect 411882 232718 447326 232954
rect 447562 232718 447646 232954
rect 447882 232718 483326 232954
rect 483562 232718 483646 232954
rect 483882 232718 519326 232954
rect 519562 232718 519646 232954
rect 519882 232718 555326 232954
rect 555562 232718 555646 232954
rect 555882 232718 588222 232954
rect 588458 232718 588542 232954
rect 588778 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -4854 232634
rect -4618 232398 -4534 232634
rect -4298 232398 15326 232634
rect 15562 232398 15646 232634
rect 15882 232398 51326 232634
rect 51562 232398 51646 232634
rect 51882 232398 87326 232634
rect 87562 232398 87646 232634
rect 87882 232398 123326 232634
rect 123562 232398 123646 232634
rect 123882 232398 159326 232634
rect 159562 232398 159646 232634
rect 159882 232398 195326 232634
rect 195562 232398 195646 232634
rect 195882 232398 231326 232634
rect 231562 232398 231646 232634
rect 231882 232398 267326 232634
rect 267562 232398 267646 232634
rect 267882 232398 303326 232634
rect 303562 232398 303646 232634
rect 303882 232398 339326 232634
rect 339562 232398 339646 232634
rect 339882 232398 375326 232634
rect 375562 232398 375646 232634
rect 375882 232398 411326 232634
rect 411562 232398 411646 232634
rect 411882 232398 447326 232634
rect 447562 232398 447646 232634
rect 447882 232398 483326 232634
rect 483562 232398 483646 232634
rect 483882 232398 519326 232634
rect 519562 232398 519646 232634
rect 519882 232398 555326 232634
rect 555562 232398 555646 232634
rect 555882 232398 588222 232634
rect 588458 232398 588542 232634
rect 588778 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -3894 228454
rect -3658 228218 -3574 228454
rect -3338 228218 10826 228454
rect 11062 228218 11146 228454
rect 11382 228218 46826 228454
rect 47062 228218 47146 228454
rect 47382 228218 82826 228454
rect 83062 228218 83146 228454
rect 83382 228218 118826 228454
rect 119062 228218 119146 228454
rect 119382 228218 154826 228454
rect 155062 228218 155146 228454
rect 155382 228218 190826 228454
rect 191062 228218 191146 228454
rect 191382 228218 226826 228454
rect 227062 228218 227146 228454
rect 227382 228218 262826 228454
rect 263062 228218 263146 228454
rect 263382 228218 298826 228454
rect 299062 228218 299146 228454
rect 299382 228218 334826 228454
rect 335062 228218 335146 228454
rect 335382 228218 370826 228454
rect 371062 228218 371146 228454
rect 371382 228218 406826 228454
rect 407062 228218 407146 228454
rect 407382 228218 442826 228454
rect 443062 228218 443146 228454
rect 443382 228218 478826 228454
rect 479062 228218 479146 228454
rect 479382 228218 514826 228454
rect 515062 228218 515146 228454
rect 515382 228218 550826 228454
rect 551062 228218 551146 228454
rect 551382 228218 587262 228454
rect 587498 228218 587582 228454
rect 587818 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -3894 228134
rect -3658 227898 -3574 228134
rect -3338 227898 10826 228134
rect 11062 227898 11146 228134
rect 11382 227898 46826 228134
rect 47062 227898 47146 228134
rect 47382 227898 82826 228134
rect 83062 227898 83146 228134
rect 83382 227898 118826 228134
rect 119062 227898 119146 228134
rect 119382 227898 154826 228134
rect 155062 227898 155146 228134
rect 155382 227898 190826 228134
rect 191062 227898 191146 228134
rect 191382 227898 226826 228134
rect 227062 227898 227146 228134
rect 227382 227898 262826 228134
rect 263062 227898 263146 228134
rect 263382 227898 298826 228134
rect 299062 227898 299146 228134
rect 299382 227898 334826 228134
rect 335062 227898 335146 228134
rect 335382 227898 370826 228134
rect 371062 227898 371146 228134
rect 371382 227898 406826 228134
rect 407062 227898 407146 228134
rect 407382 227898 442826 228134
rect 443062 227898 443146 228134
rect 443382 227898 478826 228134
rect 479062 227898 479146 228134
rect 479382 227898 514826 228134
rect 515062 227898 515146 228134
rect 515382 227898 550826 228134
rect 551062 227898 551146 228134
rect 551382 227898 587262 228134
rect 587498 227898 587582 228134
rect 587818 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 223954 592650 223986
rect -8726 223718 -2934 223954
rect -2698 223718 -2614 223954
rect -2378 223718 6326 223954
rect 6562 223718 6646 223954
rect 6882 223718 42326 223954
rect 42562 223718 42646 223954
rect 42882 223718 78326 223954
rect 78562 223718 78646 223954
rect 78882 223718 114326 223954
rect 114562 223718 114646 223954
rect 114882 223718 150326 223954
rect 150562 223718 150646 223954
rect 150882 223718 186326 223954
rect 186562 223718 186646 223954
rect 186882 223718 222326 223954
rect 222562 223718 222646 223954
rect 222882 223718 258326 223954
rect 258562 223718 258646 223954
rect 258882 223718 294326 223954
rect 294562 223718 294646 223954
rect 294882 223718 330326 223954
rect 330562 223718 330646 223954
rect 330882 223718 366326 223954
rect 366562 223718 366646 223954
rect 366882 223718 402326 223954
rect 402562 223718 402646 223954
rect 402882 223718 438326 223954
rect 438562 223718 438646 223954
rect 438882 223718 474326 223954
rect 474562 223718 474646 223954
rect 474882 223718 510326 223954
rect 510562 223718 510646 223954
rect 510882 223718 546326 223954
rect 546562 223718 546646 223954
rect 546882 223718 582326 223954
rect 582562 223718 582646 223954
rect 582882 223718 586302 223954
rect 586538 223718 586622 223954
rect 586858 223718 592650 223954
rect -8726 223634 592650 223718
rect -8726 223398 -2934 223634
rect -2698 223398 -2614 223634
rect -2378 223398 6326 223634
rect 6562 223398 6646 223634
rect 6882 223398 42326 223634
rect 42562 223398 42646 223634
rect 42882 223398 78326 223634
rect 78562 223398 78646 223634
rect 78882 223398 114326 223634
rect 114562 223398 114646 223634
rect 114882 223398 150326 223634
rect 150562 223398 150646 223634
rect 150882 223398 186326 223634
rect 186562 223398 186646 223634
rect 186882 223398 222326 223634
rect 222562 223398 222646 223634
rect 222882 223398 258326 223634
rect 258562 223398 258646 223634
rect 258882 223398 294326 223634
rect 294562 223398 294646 223634
rect 294882 223398 330326 223634
rect 330562 223398 330646 223634
rect 330882 223398 366326 223634
rect 366562 223398 366646 223634
rect 366882 223398 402326 223634
rect 402562 223398 402646 223634
rect 402882 223398 438326 223634
rect 438562 223398 438646 223634
rect 438882 223398 474326 223634
rect 474562 223398 474646 223634
rect 474882 223398 510326 223634
rect 510562 223398 510646 223634
rect 510882 223398 546326 223634
rect 546562 223398 546646 223634
rect 546882 223398 582326 223634
rect 582562 223398 582646 223634
rect 582882 223398 586302 223634
rect 586538 223398 586622 223634
rect 586858 223398 592650 223634
rect -8726 223366 592650 223398
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 214954 592650 214986
rect -8726 214718 -8694 214954
rect -8458 214718 -8374 214954
rect -8138 214718 33326 214954
rect 33562 214718 33646 214954
rect 33882 214718 249326 214954
rect 249562 214718 249646 214954
rect 249882 214718 285326 214954
rect 285562 214718 285646 214954
rect 285882 214718 357326 214954
rect 357562 214718 357646 214954
rect 357882 214718 393326 214954
rect 393562 214718 393646 214954
rect 393882 214718 429326 214954
rect 429562 214718 429646 214954
rect 429882 214718 465326 214954
rect 465562 214718 465646 214954
rect 465882 214718 501326 214954
rect 501562 214718 501646 214954
rect 501882 214718 537326 214954
rect 537562 214718 537646 214954
rect 537882 214718 573326 214954
rect 573562 214718 573646 214954
rect 573882 214718 592062 214954
rect 592298 214718 592382 214954
rect 592618 214718 592650 214954
rect -8726 214634 592650 214718
rect -8726 214398 -8694 214634
rect -8458 214398 -8374 214634
rect -8138 214398 33326 214634
rect 33562 214398 33646 214634
rect 33882 214398 249326 214634
rect 249562 214398 249646 214634
rect 249882 214398 285326 214634
rect 285562 214398 285646 214634
rect 285882 214398 357326 214634
rect 357562 214398 357646 214634
rect 357882 214398 393326 214634
rect 393562 214398 393646 214634
rect 393882 214398 429326 214634
rect 429562 214398 429646 214634
rect 429882 214398 465326 214634
rect 465562 214398 465646 214634
rect 465882 214398 501326 214634
rect 501562 214398 501646 214634
rect 501882 214398 537326 214634
rect 537562 214398 537646 214634
rect 537882 214398 573326 214634
rect 573562 214398 573646 214634
rect 573882 214398 592062 214634
rect 592298 214398 592382 214634
rect 592618 214398 592650 214634
rect -8726 214366 592650 214398
rect -8726 210454 592650 210486
rect -8726 210218 -7734 210454
rect -7498 210218 -7414 210454
rect -7178 210218 28826 210454
rect 29062 210218 29146 210454
rect 29382 210218 244826 210454
rect 245062 210218 245146 210454
rect 245382 210218 280826 210454
rect 281062 210218 281146 210454
rect 281382 210218 352826 210454
rect 353062 210218 353146 210454
rect 353382 210218 388826 210454
rect 389062 210218 389146 210454
rect 389382 210218 424826 210454
rect 425062 210218 425146 210454
rect 425382 210218 460826 210454
rect 461062 210218 461146 210454
rect 461382 210218 496826 210454
rect 497062 210218 497146 210454
rect 497382 210218 532826 210454
rect 533062 210218 533146 210454
rect 533382 210218 568826 210454
rect 569062 210218 569146 210454
rect 569382 210218 591102 210454
rect 591338 210218 591422 210454
rect 591658 210218 592650 210454
rect -8726 210134 592650 210218
rect -8726 209898 -7734 210134
rect -7498 209898 -7414 210134
rect -7178 209898 28826 210134
rect 29062 209898 29146 210134
rect 29382 209898 244826 210134
rect 245062 209898 245146 210134
rect 245382 209898 280826 210134
rect 281062 209898 281146 210134
rect 281382 209898 352826 210134
rect 353062 209898 353146 210134
rect 353382 209898 388826 210134
rect 389062 209898 389146 210134
rect 389382 209898 424826 210134
rect 425062 209898 425146 210134
rect 425382 209898 460826 210134
rect 461062 209898 461146 210134
rect 461382 209898 496826 210134
rect 497062 209898 497146 210134
rect 497382 209898 532826 210134
rect 533062 209898 533146 210134
rect 533382 209898 568826 210134
rect 569062 209898 569146 210134
rect 569382 209898 591102 210134
rect 591338 209898 591422 210134
rect 591658 209898 592650 210134
rect -8726 209866 592650 209898
rect -8726 205954 592650 205986
rect -8726 205718 -6774 205954
rect -6538 205718 -6454 205954
rect -6218 205718 24326 205954
rect 24562 205718 24646 205954
rect 24882 205718 240326 205954
rect 240562 205718 240646 205954
rect 240882 205718 276326 205954
rect 276562 205718 276646 205954
rect 276882 205718 348326 205954
rect 348562 205718 348646 205954
rect 348882 205718 384326 205954
rect 384562 205718 384646 205954
rect 384882 205718 420326 205954
rect 420562 205718 420646 205954
rect 420882 205718 456326 205954
rect 456562 205718 456646 205954
rect 456882 205718 492326 205954
rect 492562 205718 492646 205954
rect 492882 205718 528326 205954
rect 528562 205718 528646 205954
rect 528882 205718 564326 205954
rect 564562 205718 564646 205954
rect 564882 205718 590142 205954
rect 590378 205718 590462 205954
rect 590698 205718 592650 205954
rect -8726 205634 592650 205718
rect -8726 205398 -6774 205634
rect -6538 205398 -6454 205634
rect -6218 205398 24326 205634
rect 24562 205398 24646 205634
rect 24882 205398 240326 205634
rect 240562 205398 240646 205634
rect 240882 205398 276326 205634
rect 276562 205398 276646 205634
rect 276882 205398 348326 205634
rect 348562 205398 348646 205634
rect 348882 205398 384326 205634
rect 384562 205398 384646 205634
rect 384882 205398 420326 205634
rect 420562 205398 420646 205634
rect 420882 205398 456326 205634
rect 456562 205398 456646 205634
rect 456882 205398 492326 205634
rect 492562 205398 492646 205634
rect 492882 205398 528326 205634
rect 528562 205398 528646 205634
rect 528882 205398 564326 205634
rect 564562 205398 564646 205634
rect 564882 205398 590142 205634
rect 590378 205398 590462 205634
rect 590698 205398 592650 205634
rect -8726 205366 592650 205398
rect -8726 201454 592650 201486
rect -8726 201218 -5814 201454
rect -5578 201218 -5494 201454
rect -5258 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 589182 201454
rect 589418 201218 589502 201454
rect 589738 201218 592650 201454
rect -8726 201134 592650 201218
rect -8726 200898 -5814 201134
rect -5578 200898 -5494 201134
rect -5258 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 589182 201134
rect 589418 200898 589502 201134
rect 589738 200898 592650 201134
rect -8726 200866 592650 200898
rect -8726 196954 592650 196986
rect -8726 196718 -4854 196954
rect -4618 196718 -4534 196954
rect -4298 196718 15326 196954
rect 15562 196718 15646 196954
rect 15882 196718 51326 196954
rect 51562 196718 51646 196954
rect 51882 196718 231326 196954
rect 231562 196718 231646 196954
rect 231882 196718 267326 196954
rect 267562 196718 267646 196954
rect 267882 196718 375326 196954
rect 375562 196718 375646 196954
rect 375882 196718 411326 196954
rect 411562 196718 411646 196954
rect 411882 196718 447326 196954
rect 447562 196718 447646 196954
rect 447882 196718 483326 196954
rect 483562 196718 483646 196954
rect 483882 196718 519326 196954
rect 519562 196718 519646 196954
rect 519882 196718 555326 196954
rect 555562 196718 555646 196954
rect 555882 196718 588222 196954
rect 588458 196718 588542 196954
rect 588778 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -4854 196634
rect -4618 196398 -4534 196634
rect -4298 196398 15326 196634
rect 15562 196398 15646 196634
rect 15882 196398 51326 196634
rect 51562 196398 51646 196634
rect 51882 196398 231326 196634
rect 231562 196398 231646 196634
rect 231882 196398 267326 196634
rect 267562 196398 267646 196634
rect 267882 196398 375326 196634
rect 375562 196398 375646 196634
rect 375882 196398 411326 196634
rect 411562 196398 411646 196634
rect 411882 196398 447326 196634
rect 447562 196398 447646 196634
rect 447882 196398 483326 196634
rect 483562 196398 483646 196634
rect 483882 196398 519326 196634
rect 519562 196398 519646 196634
rect 519882 196398 555326 196634
rect 555562 196398 555646 196634
rect 555882 196398 588222 196634
rect 588458 196398 588542 196634
rect 588778 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -3894 192454
rect -3658 192218 -3574 192454
rect -3338 192218 10826 192454
rect 11062 192218 11146 192454
rect 11382 192218 46826 192454
rect 47062 192218 47146 192454
rect 47382 192218 226826 192454
rect 227062 192218 227146 192454
rect 227382 192218 262826 192454
rect 263062 192218 263146 192454
rect 263382 192218 370826 192454
rect 371062 192218 371146 192454
rect 371382 192218 406826 192454
rect 407062 192218 407146 192454
rect 407382 192218 442826 192454
rect 443062 192218 443146 192454
rect 443382 192218 478826 192454
rect 479062 192218 479146 192454
rect 479382 192218 514826 192454
rect 515062 192218 515146 192454
rect 515382 192218 550826 192454
rect 551062 192218 551146 192454
rect 551382 192218 587262 192454
rect 587498 192218 587582 192454
rect 587818 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -3894 192134
rect -3658 191898 -3574 192134
rect -3338 191898 10826 192134
rect 11062 191898 11146 192134
rect 11382 191898 46826 192134
rect 47062 191898 47146 192134
rect 47382 191898 226826 192134
rect 227062 191898 227146 192134
rect 227382 191898 262826 192134
rect 263062 191898 263146 192134
rect 263382 191898 370826 192134
rect 371062 191898 371146 192134
rect 371382 191898 406826 192134
rect 407062 191898 407146 192134
rect 407382 191898 442826 192134
rect 443062 191898 443146 192134
rect 443382 191898 478826 192134
rect 479062 191898 479146 192134
rect 479382 191898 514826 192134
rect 515062 191898 515146 192134
rect 515382 191898 550826 192134
rect 551062 191898 551146 192134
rect 551382 191898 587262 192134
rect 587498 191898 587582 192134
rect 587818 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 187954 592650 187986
rect -8726 187718 -2934 187954
rect -2698 187718 -2614 187954
rect -2378 187718 6326 187954
rect 6562 187718 6646 187954
rect 6882 187718 42326 187954
rect 42562 187718 42646 187954
rect 42882 187718 79610 187954
rect 79846 187718 110330 187954
rect 110566 187718 141050 187954
rect 141286 187718 171770 187954
rect 172006 187718 202490 187954
rect 202726 187718 258326 187954
rect 258562 187718 258646 187954
rect 258882 187718 294326 187954
rect 294562 187718 294646 187954
rect 294882 187718 319610 187954
rect 319846 187718 366326 187954
rect 366562 187718 366646 187954
rect 366882 187718 402326 187954
rect 402562 187718 402646 187954
rect 402882 187718 438326 187954
rect 438562 187718 438646 187954
rect 438882 187718 474326 187954
rect 474562 187718 474646 187954
rect 474882 187718 510326 187954
rect 510562 187718 510646 187954
rect 510882 187718 546326 187954
rect 546562 187718 546646 187954
rect 546882 187718 582326 187954
rect 582562 187718 582646 187954
rect 582882 187718 586302 187954
rect 586538 187718 586622 187954
rect 586858 187718 592650 187954
rect -8726 187634 592650 187718
rect -8726 187398 -2934 187634
rect -2698 187398 -2614 187634
rect -2378 187398 6326 187634
rect 6562 187398 6646 187634
rect 6882 187398 42326 187634
rect 42562 187398 42646 187634
rect 42882 187398 79610 187634
rect 79846 187398 110330 187634
rect 110566 187398 141050 187634
rect 141286 187398 171770 187634
rect 172006 187398 202490 187634
rect 202726 187398 258326 187634
rect 258562 187398 258646 187634
rect 258882 187398 294326 187634
rect 294562 187398 294646 187634
rect 294882 187398 319610 187634
rect 319846 187398 366326 187634
rect 366562 187398 366646 187634
rect 366882 187398 402326 187634
rect 402562 187398 402646 187634
rect 402882 187398 438326 187634
rect 438562 187398 438646 187634
rect 438882 187398 474326 187634
rect 474562 187398 474646 187634
rect 474882 187398 510326 187634
rect 510562 187398 510646 187634
rect 510882 187398 546326 187634
rect 546562 187398 546646 187634
rect 546882 187398 582326 187634
rect 582562 187398 582646 187634
rect 582882 187398 586302 187634
rect 586538 187398 586622 187634
rect 586858 187398 592650 187634
rect -8726 187366 592650 187398
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 64250 183454
rect 64486 183218 94970 183454
rect 95206 183218 125690 183454
rect 125926 183218 156410 183454
rect 156646 183218 187130 183454
rect 187366 183218 217850 183454
rect 218086 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 304250 183454
rect 304486 183218 334970 183454
rect 335206 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 64250 183134
rect 64486 182898 94970 183134
rect 95206 182898 125690 183134
rect 125926 182898 156410 183134
rect 156646 182898 187130 183134
rect 187366 182898 217850 183134
rect 218086 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 304250 183134
rect 304486 182898 334970 183134
rect 335206 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 178954 592650 178986
rect -8726 178718 -8694 178954
rect -8458 178718 -8374 178954
rect -8138 178718 33326 178954
rect 33562 178718 33646 178954
rect 33882 178718 249326 178954
rect 249562 178718 249646 178954
rect 249882 178718 285326 178954
rect 285562 178718 285646 178954
rect 285882 178718 357326 178954
rect 357562 178718 357646 178954
rect 357882 178718 393326 178954
rect 393562 178718 393646 178954
rect 393882 178718 429326 178954
rect 429562 178718 429646 178954
rect 429882 178718 465326 178954
rect 465562 178718 465646 178954
rect 465882 178718 501326 178954
rect 501562 178718 501646 178954
rect 501882 178718 537326 178954
rect 537562 178718 537646 178954
rect 537882 178718 573326 178954
rect 573562 178718 573646 178954
rect 573882 178718 592062 178954
rect 592298 178718 592382 178954
rect 592618 178718 592650 178954
rect -8726 178634 592650 178718
rect -8726 178398 -8694 178634
rect -8458 178398 -8374 178634
rect -8138 178398 33326 178634
rect 33562 178398 33646 178634
rect 33882 178398 249326 178634
rect 249562 178398 249646 178634
rect 249882 178398 285326 178634
rect 285562 178398 285646 178634
rect 285882 178398 357326 178634
rect 357562 178398 357646 178634
rect 357882 178398 393326 178634
rect 393562 178398 393646 178634
rect 393882 178398 429326 178634
rect 429562 178398 429646 178634
rect 429882 178398 465326 178634
rect 465562 178398 465646 178634
rect 465882 178398 501326 178634
rect 501562 178398 501646 178634
rect 501882 178398 537326 178634
rect 537562 178398 537646 178634
rect 537882 178398 573326 178634
rect 573562 178398 573646 178634
rect 573882 178398 592062 178634
rect 592298 178398 592382 178634
rect 592618 178398 592650 178634
rect -8726 178366 592650 178398
rect -8726 174454 592650 174486
rect -8726 174218 -7734 174454
rect -7498 174218 -7414 174454
rect -7178 174218 28826 174454
rect 29062 174218 29146 174454
rect 29382 174218 244826 174454
rect 245062 174218 245146 174454
rect 245382 174218 280826 174454
rect 281062 174218 281146 174454
rect 281382 174218 352826 174454
rect 353062 174218 353146 174454
rect 353382 174218 388826 174454
rect 389062 174218 389146 174454
rect 389382 174218 424826 174454
rect 425062 174218 425146 174454
rect 425382 174218 460826 174454
rect 461062 174218 461146 174454
rect 461382 174218 496826 174454
rect 497062 174218 497146 174454
rect 497382 174218 532826 174454
rect 533062 174218 533146 174454
rect 533382 174218 568826 174454
rect 569062 174218 569146 174454
rect 569382 174218 591102 174454
rect 591338 174218 591422 174454
rect 591658 174218 592650 174454
rect -8726 174134 592650 174218
rect -8726 173898 -7734 174134
rect -7498 173898 -7414 174134
rect -7178 173898 28826 174134
rect 29062 173898 29146 174134
rect 29382 173898 244826 174134
rect 245062 173898 245146 174134
rect 245382 173898 280826 174134
rect 281062 173898 281146 174134
rect 281382 173898 352826 174134
rect 353062 173898 353146 174134
rect 353382 173898 388826 174134
rect 389062 173898 389146 174134
rect 389382 173898 424826 174134
rect 425062 173898 425146 174134
rect 425382 173898 460826 174134
rect 461062 173898 461146 174134
rect 461382 173898 496826 174134
rect 497062 173898 497146 174134
rect 497382 173898 532826 174134
rect 533062 173898 533146 174134
rect 533382 173898 568826 174134
rect 569062 173898 569146 174134
rect 569382 173898 591102 174134
rect 591338 173898 591422 174134
rect 591658 173898 592650 174134
rect -8726 173866 592650 173898
rect -8726 169954 592650 169986
rect -8726 169718 -6774 169954
rect -6538 169718 -6454 169954
rect -6218 169718 24326 169954
rect 24562 169718 24646 169954
rect 24882 169718 240326 169954
rect 240562 169718 240646 169954
rect 240882 169718 276326 169954
rect 276562 169718 276646 169954
rect 276882 169718 348326 169954
rect 348562 169718 348646 169954
rect 348882 169718 384326 169954
rect 384562 169718 384646 169954
rect 384882 169718 420326 169954
rect 420562 169718 420646 169954
rect 420882 169718 456326 169954
rect 456562 169718 456646 169954
rect 456882 169718 492326 169954
rect 492562 169718 492646 169954
rect 492882 169718 528326 169954
rect 528562 169718 528646 169954
rect 528882 169718 564326 169954
rect 564562 169718 564646 169954
rect 564882 169718 590142 169954
rect 590378 169718 590462 169954
rect 590698 169718 592650 169954
rect -8726 169634 592650 169718
rect -8726 169398 -6774 169634
rect -6538 169398 -6454 169634
rect -6218 169398 24326 169634
rect 24562 169398 24646 169634
rect 24882 169398 240326 169634
rect 240562 169398 240646 169634
rect 240882 169398 276326 169634
rect 276562 169398 276646 169634
rect 276882 169398 348326 169634
rect 348562 169398 348646 169634
rect 348882 169398 384326 169634
rect 384562 169398 384646 169634
rect 384882 169398 420326 169634
rect 420562 169398 420646 169634
rect 420882 169398 456326 169634
rect 456562 169398 456646 169634
rect 456882 169398 492326 169634
rect 492562 169398 492646 169634
rect 492882 169398 528326 169634
rect 528562 169398 528646 169634
rect 528882 169398 564326 169634
rect 564562 169398 564646 169634
rect 564882 169398 590142 169634
rect 590378 169398 590462 169634
rect 590698 169398 592650 169634
rect -8726 169366 592650 169398
rect -8726 165454 592650 165486
rect -8726 165218 -5814 165454
rect -5578 165218 -5494 165454
rect -5258 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 589182 165454
rect 589418 165218 589502 165454
rect 589738 165218 592650 165454
rect -8726 165134 592650 165218
rect -8726 164898 -5814 165134
rect -5578 164898 -5494 165134
rect -5258 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 589182 165134
rect 589418 164898 589502 165134
rect 589738 164898 592650 165134
rect -8726 164866 592650 164898
rect -8726 160954 592650 160986
rect -8726 160718 -4854 160954
rect -4618 160718 -4534 160954
rect -4298 160718 15326 160954
rect 15562 160718 15646 160954
rect 15882 160718 51326 160954
rect 51562 160718 51646 160954
rect 51882 160718 231326 160954
rect 231562 160718 231646 160954
rect 231882 160718 267326 160954
rect 267562 160718 267646 160954
rect 267882 160718 375326 160954
rect 375562 160718 375646 160954
rect 375882 160718 411326 160954
rect 411562 160718 411646 160954
rect 411882 160718 447326 160954
rect 447562 160718 447646 160954
rect 447882 160718 483326 160954
rect 483562 160718 483646 160954
rect 483882 160718 519326 160954
rect 519562 160718 519646 160954
rect 519882 160718 555326 160954
rect 555562 160718 555646 160954
rect 555882 160718 588222 160954
rect 588458 160718 588542 160954
rect 588778 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -4854 160634
rect -4618 160398 -4534 160634
rect -4298 160398 15326 160634
rect 15562 160398 15646 160634
rect 15882 160398 51326 160634
rect 51562 160398 51646 160634
rect 51882 160398 231326 160634
rect 231562 160398 231646 160634
rect 231882 160398 267326 160634
rect 267562 160398 267646 160634
rect 267882 160398 375326 160634
rect 375562 160398 375646 160634
rect 375882 160398 411326 160634
rect 411562 160398 411646 160634
rect 411882 160398 447326 160634
rect 447562 160398 447646 160634
rect 447882 160398 483326 160634
rect 483562 160398 483646 160634
rect 483882 160398 519326 160634
rect 519562 160398 519646 160634
rect 519882 160398 555326 160634
rect 555562 160398 555646 160634
rect 555882 160398 588222 160634
rect 588458 160398 588542 160634
rect 588778 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -3894 156454
rect -3658 156218 -3574 156454
rect -3338 156218 10826 156454
rect 11062 156218 11146 156454
rect 11382 156218 46826 156454
rect 47062 156218 47146 156454
rect 47382 156218 226826 156454
rect 227062 156218 227146 156454
rect 227382 156218 262826 156454
rect 263062 156218 263146 156454
rect 263382 156218 370826 156454
rect 371062 156218 371146 156454
rect 371382 156218 406826 156454
rect 407062 156218 407146 156454
rect 407382 156218 442826 156454
rect 443062 156218 443146 156454
rect 443382 156218 478826 156454
rect 479062 156218 479146 156454
rect 479382 156218 514826 156454
rect 515062 156218 515146 156454
rect 515382 156218 550826 156454
rect 551062 156218 551146 156454
rect 551382 156218 587262 156454
rect 587498 156218 587582 156454
rect 587818 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -3894 156134
rect -3658 155898 -3574 156134
rect -3338 155898 10826 156134
rect 11062 155898 11146 156134
rect 11382 155898 46826 156134
rect 47062 155898 47146 156134
rect 47382 155898 226826 156134
rect 227062 155898 227146 156134
rect 227382 155898 262826 156134
rect 263062 155898 263146 156134
rect 263382 155898 370826 156134
rect 371062 155898 371146 156134
rect 371382 155898 406826 156134
rect 407062 155898 407146 156134
rect 407382 155898 442826 156134
rect 443062 155898 443146 156134
rect 443382 155898 478826 156134
rect 479062 155898 479146 156134
rect 479382 155898 514826 156134
rect 515062 155898 515146 156134
rect 515382 155898 550826 156134
rect 551062 155898 551146 156134
rect 551382 155898 587262 156134
rect 587498 155898 587582 156134
rect 587818 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 151954 592650 151986
rect -8726 151718 -2934 151954
rect -2698 151718 -2614 151954
rect -2378 151718 6326 151954
rect 6562 151718 6646 151954
rect 6882 151718 42326 151954
rect 42562 151718 42646 151954
rect 42882 151718 79610 151954
rect 79846 151718 110330 151954
rect 110566 151718 141050 151954
rect 141286 151718 171770 151954
rect 172006 151718 202490 151954
rect 202726 151718 258326 151954
rect 258562 151718 258646 151954
rect 258882 151718 294326 151954
rect 294562 151718 294646 151954
rect 294882 151718 319610 151954
rect 319846 151718 366326 151954
rect 366562 151718 366646 151954
rect 366882 151718 402326 151954
rect 402562 151718 402646 151954
rect 402882 151718 438326 151954
rect 438562 151718 438646 151954
rect 438882 151718 474326 151954
rect 474562 151718 474646 151954
rect 474882 151718 510326 151954
rect 510562 151718 510646 151954
rect 510882 151718 546326 151954
rect 546562 151718 546646 151954
rect 546882 151718 582326 151954
rect 582562 151718 582646 151954
rect 582882 151718 586302 151954
rect 586538 151718 586622 151954
rect 586858 151718 592650 151954
rect -8726 151634 592650 151718
rect -8726 151398 -2934 151634
rect -2698 151398 -2614 151634
rect -2378 151398 6326 151634
rect 6562 151398 6646 151634
rect 6882 151398 42326 151634
rect 42562 151398 42646 151634
rect 42882 151398 79610 151634
rect 79846 151398 110330 151634
rect 110566 151398 141050 151634
rect 141286 151398 171770 151634
rect 172006 151398 202490 151634
rect 202726 151398 258326 151634
rect 258562 151398 258646 151634
rect 258882 151398 294326 151634
rect 294562 151398 294646 151634
rect 294882 151398 319610 151634
rect 319846 151398 366326 151634
rect 366562 151398 366646 151634
rect 366882 151398 402326 151634
rect 402562 151398 402646 151634
rect 402882 151398 438326 151634
rect 438562 151398 438646 151634
rect 438882 151398 474326 151634
rect 474562 151398 474646 151634
rect 474882 151398 510326 151634
rect 510562 151398 510646 151634
rect 510882 151398 546326 151634
rect 546562 151398 546646 151634
rect 546882 151398 582326 151634
rect 582562 151398 582646 151634
rect 582882 151398 586302 151634
rect 586538 151398 586622 151634
rect 586858 151398 592650 151634
rect -8726 151366 592650 151398
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 304250 147454
rect 304486 147218 334970 147454
rect 335206 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 304250 147134
rect 304486 146898 334970 147134
rect 335206 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 142954 592650 142986
rect -8726 142718 -8694 142954
rect -8458 142718 -8374 142954
rect -8138 142718 33326 142954
rect 33562 142718 33646 142954
rect 33882 142718 249326 142954
rect 249562 142718 249646 142954
rect 249882 142718 285326 142954
rect 285562 142718 285646 142954
rect 285882 142718 357326 142954
rect 357562 142718 357646 142954
rect 357882 142718 393326 142954
rect 393562 142718 393646 142954
rect 393882 142718 429326 142954
rect 429562 142718 429646 142954
rect 429882 142718 465326 142954
rect 465562 142718 465646 142954
rect 465882 142718 501326 142954
rect 501562 142718 501646 142954
rect 501882 142718 537326 142954
rect 537562 142718 537646 142954
rect 537882 142718 573326 142954
rect 573562 142718 573646 142954
rect 573882 142718 592062 142954
rect 592298 142718 592382 142954
rect 592618 142718 592650 142954
rect -8726 142634 592650 142718
rect -8726 142398 -8694 142634
rect -8458 142398 -8374 142634
rect -8138 142398 33326 142634
rect 33562 142398 33646 142634
rect 33882 142398 249326 142634
rect 249562 142398 249646 142634
rect 249882 142398 285326 142634
rect 285562 142398 285646 142634
rect 285882 142398 357326 142634
rect 357562 142398 357646 142634
rect 357882 142398 393326 142634
rect 393562 142398 393646 142634
rect 393882 142398 429326 142634
rect 429562 142398 429646 142634
rect 429882 142398 465326 142634
rect 465562 142398 465646 142634
rect 465882 142398 501326 142634
rect 501562 142398 501646 142634
rect 501882 142398 537326 142634
rect 537562 142398 537646 142634
rect 537882 142398 573326 142634
rect 573562 142398 573646 142634
rect 573882 142398 592062 142634
rect 592298 142398 592382 142634
rect 592618 142398 592650 142634
rect -8726 142366 592650 142398
rect -8726 138454 592650 138486
rect -8726 138218 -7734 138454
rect -7498 138218 -7414 138454
rect -7178 138218 28826 138454
rect 29062 138218 29146 138454
rect 29382 138218 244826 138454
rect 245062 138218 245146 138454
rect 245382 138218 280826 138454
rect 281062 138218 281146 138454
rect 281382 138218 352826 138454
rect 353062 138218 353146 138454
rect 353382 138218 388826 138454
rect 389062 138218 389146 138454
rect 389382 138218 424826 138454
rect 425062 138218 425146 138454
rect 425382 138218 460826 138454
rect 461062 138218 461146 138454
rect 461382 138218 496826 138454
rect 497062 138218 497146 138454
rect 497382 138218 532826 138454
rect 533062 138218 533146 138454
rect 533382 138218 568826 138454
rect 569062 138218 569146 138454
rect 569382 138218 591102 138454
rect 591338 138218 591422 138454
rect 591658 138218 592650 138454
rect -8726 138134 592650 138218
rect -8726 137898 -7734 138134
rect -7498 137898 -7414 138134
rect -7178 137898 28826 138134
rect 29062 137898 29146 138134
rect 29382 137898 244826 138134
rect 245062 137898 245146 138134
rect 245382 137898 280826 138134
rect 281062 137898 281146 138134
rect 281382 137898 352826 138134
rect 353062 137898 353146 138134
rect 353382 137898 388826 138134
rect 389062 137898 389146 138134
rect 389382 137898 424826 138134
rect 425062 137898 425146 138134
rect 425382 137898 460826 138134
rect 461062 137898 461146 138134
rect 461382 137898 496826 138134
rect 497062 137898 497146 138134
rect 497382 137898 532826 138134
rect 533062 137898 533146 138134
rect 533382 137898 568826 138134
rect 569062 137898 569146 138134
rect 569382 137898 591102 138134
rect 591338 137898 591422 138134
rect 591658 137898 592650 138134
rect -8726 137866 592650 137898
rect -8726 133954 592650 133986
rect -8726 133718 -6774 133954
rect -6538 133718 -6454 133954
rect -6218 133718 24326 133954
rect 24562 133718 24646 133954
rect 24882 133718 240326 133954
rect 240562 133718 240646 133954
rect 240882 133718 276326 133954
rect 276562 133718 276646 133954
rect 276882 133718 348326 133954
rect 348562 133718 348646 133954
rect 348882 133718 384326 133954
rect 384562 133718 384646 133954
rect 384882 133718 420326 133954
rect 420562 133718 420646 133954
rect 420882 133718 456326 133954
rect 456562 133718 456646 133954
rect 456882 133718 492326 133954
rect 492562 133718 492646 133954
rect 492882 133718 528326 133954
rect 528562 133718 528646 133954
rect 528882 133718 564326 133954
rect 564562 133718 564646 133954
rect 564882 133718 590142 133954
rect 590378 133718 590462 133954
rect 590698 133718 592650 133954
rect -8726 133634 592650 133718
rect -8726 133398 -6774 133634
rect -6538 133398 -6454 133634
rect -6218 133398 24326 133634
rect 24562 133398 24646 133634
rect 24882 133398 240326 133634
rect 240562 133398 240646 133634
rect 240882 133398 276326 133634
rect 276562 133398 276646 133634
rect 276882 133398 348326 133634
rect 348562 133398 348646 133634
rect 348882 133398 384326 133634
rect 384562 133398 384646 133634
rect 384882 133398 420326 133634
rect 420562 133398 420646 133634
rect 420882 133398 456326 133634
rect 456562 133398 456646 133634
rect 456882 133398 492326 133634
rect 492562 133398 492646 133634
rect 492882 133398 528326 133634
rect 528562 133398 528646 133634
rect 528882 133398 564326 133634
rect 564562 133398 564646 133634
rect 564882 133398 590142 133634
rect 590378 133398 590462 133634
rect 590698 133398 592650 133634
rect -8726 133366 592650 133398
rect -8726 129454 592650 129486
rect -8726 129218 -5814 129454
rect -5578 129218 -5494 129454
rect -5258 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 589182 129454
rect 589418 129218 589502 129454
rect 589738 129218 592650 129454
rect -8726 129134 592650 129218
rect -8726 128898 -5814 129134
rect -5578 128898 -5494 129134
rect -5258 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 589182 129134
rect 589418 128898 589502 129134
rect 589738 128898 592650 129134
rect -8726 128866 592650 128898
rect -8726 124954 592650 124986
rect -8726 124718 -4854 124954
rect -4618 124718 -4534 124954
rect -4298 124718 15326 124954
rect 15562 124718 15646 124954
rect 15882 124718 51326 124954
rect 51562 124718 51646 124954
rect 51882 124718 231326 124954
rect 231562 124718 231646 124954
rect 231882 124718 267326 124954
rect 267562 124718 267646 124954
rect 267882 124718 375326 124954
rect 375562 124718 375646 124954
rect 375882 124718 411326 124954
rect 411562 124718 411646 124954
rect 411882 124718 447326 124954
rect 447562 124718 447646 124954
rect 447882 124718 483326 124954
rect 483562 124718 483646 124954
rect 483882 124718 519326 124954
rect 519562 124718 519646 124954
rect 519882 124718 555326 124954
rect 555562 124718 555646 124954
rect 555882 124718 588222 124954
rect 588458 124718 588542 124954
rect 588778 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -4854 124634
rect -4618 124398 -4534 124634
rect -4298 124398 15326 124634
rect 15562 124398 15646 124634
rect 15882 124398 51326 124634
rect 51562 124398 51646 124634
rect 51882 124398 231326 124634
rect 231562 124398 231646 124634
rect 231882 124398 267326 124634
rect 267562 124398 267646 124634
rect 267882 124398 375326 124634
rect 375562 124398 375646 124634
rect 375882 124398 411326 124634
rect 411562 124398 411646 124634
rect 411882 124398 447326 124634
rect 447562 124398 447646 124634
rect 447882 124398 483326 124634
rect 483562 124398 483646 124634
rect 483882 124398 519326 124634
rect 519562 124398 519646 124634
rect 519882 124398 555326 124634
rect 555562 124398 555646 124634
rect 555882 124398 588222 124634
rect 588458 124398 588542 124634
rect 588778 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -3894 120454
rect -3658 120218 -3574 120454
rect -3338 120218 10826 120454
rect 11062 120218 11146 120454
rect 11382 120218 46826 120454
rect 47062 120218 47146 120454
rect 47382 120218 226826 120454
rect 227062 120218 227146 120454
rect 227382 120218 262826 120454
rect 263062 120218 263146 120454
rect 263382 120218 370826 120454
rect 371062 120218 371146 120454
rect 371382 120218 406826 120454
rect 407062 120218 407146 120454
rect 407382 120218 442826 120454
rect 443062 120218 443146 120454
rect 443382 120218 478826 120454
rect 479062 120218 479146 120454
rect 479382 120218 514826 120454
rect 515062 120218 515146 120454
rect 515382 120218 550826 120454
rect 551062 120218 551146 120454
rect 551382 120218 587262 120454
rect 587498 120218 587582 120454
rect 587818 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -3894 120134
rect -3658 119898 -3574 120134
rect -3338 119898 10826 120134
rect 11062 119898 11146 120134
rect 11382 119898 46826 120134
rect 47062 119898 47146 120134
rect 47382 119898 226826 120134
rect 227062 119898 227146 120134
rect 227382 119898 262826 120134
rect 263062 119898 263146 120134
rect 263382 119898 370826 120134
rect 371062 119898 371146 120134
rect 371382 119898 406826 120134
rect 407062 119898 407146 120134
rect 407382 119898 442826 120134
rect 443062 119898 443146 120134
rect 443382 119898 478826 120134
rect 479062 119898 479146 120134
rect 479382 119898 514826 120134
rect 515062 119898 515146 120134
rect 515382 119898 550826 120134
rect 551062 119898 551146 120134
rect 551382 119898 587262 120134
rect 587498 119898 587582 120134
rect 587818 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 115954 592650 115986
rect -8726 115718 -2934 115954
rect -2698 115718 -2614 115954
rect -2378 115718 6326 115954
rect 6562 115718 6646 115954
rect 6882 115718 42326 115954
rect 42562 115718 42646 115954
rect 42882 115718 79610 115954
rect 79846 115718 110330 115954
rect 110566 115718 141050 115954
rect 141286 115718 171770 115954
rect 172006 115718 202490 115954
rect 202726 115718 258326 115954
rect 258562 115718 258646 115954
rect 258882 115718 294326 115954
rect 294562 115718 294646 115954
rect 294882 115718 319610 115954
rect 319846 115718 366326 115954
rect 366562 115718 366646 115954
rect 366882 115718 402326 115954
rect 402562 115718 402646 115954
rect 402882 115718 438326 115954
rect 438562 115718 438646 115954
rect 438882 115718 474326 115954
rect 474562 115718 474646 115954
rect 474882 115718 510326 115954
rect 510562 115718 510646 115954
rect 510882 115718 546326 115954
rect 546562 115718 546646 115954
rect 546882 115718 582326 115954
rect 582562 115718 582646 115954
rect 582882 115718 586302 115954
rect 586538 115718 586622 115954
rect 586858 115718 592650 115954
rect -8726 115634 592650 115718
rect -8726 115398 -2934 115634
rect -2698 115398 -2614 115634
rect -2378 115398 6326 115634
rect 6562 115398 6646 115634
rect 6882 115398 42326 115634
rect 42562 115398 42646 115634
rect 42882 115398 79610 115634
rect 79846 115398 110330 115634
rect 110566 115398 141050 115634
rect 141286 115398 171770 115634
rect 172006 115398 202490 115634
rect 202726 115398 258326 115634
rect 258562 115398 258646 115634
rect 258882 115398 294326 115634
rect 294562 115398 294646 115634
rect 294882 115398 319610 115634
rect 319846 115398 366326 115634
rect 366562 115398 366646 115634
rect 366882 115398 402326 115634
rect 402562 115398 402646 115634
rect 402882 115398 438326 115634
rect 438562 115398 438646 115634
rect 438882 115398 474326 115634
rect 474562 115398 474646 115634
rect 474882 115398 510326 115634
rect 510562 115398 510646 115634
rect 510882 115398 546326 115634
rect 546562 115398 546646 115634
rect 546882 115398 582326 115634
rect 582562 115398 582646 115634
rect 582882 115398 586302 115634
rect 586538 115398 586622 115634
rect 586858 115398 592650 115634
rect -8726 115366 592650 115398
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 304250 111454
rect 304486 111218 334970 111454
rect 335206 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 304250 111134
rect 304486 110898 334970 111134
rect 335206 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 106954 592650 106986
rect -8726 106718 -8694 106954
rect -8458 106718 -8374 106954
rect -8138 106718 33326 106954
rect 33562 106718 33646 106954
rect 33882 106718 249326 106954
rect 249562 106718 249646 106954
rect 249882 106718 285326 106954
rect 285562 106718 285646 106954
rect 285882 106718 357326 106954
rect 357562 106718 357646 106954
rect 357882 106718 393326 106954
rect 393562 106718 393646 106954
rect 393882 106718 429326 106954
rect 429562 106718 429646 106954
rect 429882 106718 465326 106954
rect 465562 106718 465646 106954
rect 465882 106718 501326 106954
rect 501562 106718 501646 106954
rect 501882 106718 537326 106954
rect 537562 106718 537646 106954
rect 537882 106718 573326 106954
rect 573562 106718 573646 106954
rect 573882 106718 592062 106954
rect 592298 106718 592382 106954
rect 592618 106718 592650 106954
rect -8726 106634 592650 106718
rect -8726 106398 -8694 106634
rect -8458 106398 -8374 106634
rect -8138 106398 33326 106634
rect 33562 106398 33646 106634
rect 33882 106398 249326 106634
rect 249562 106398 249646 106634
rect 249882 106398 285326 106634
rect 285562 106398 285646 106634
rect 285882 106398 357326 106634
rect 357562 106398 357646 106634
rect 357882 106398 393326 106634
rect 393562 106398 393646 106634
rect 393882 106398 429326 106634
rect 429562 106398 429646 106634
rect 429882 106398 465326 106634
rect 465562 106398 465646 106634
rect 465882 106398 501326 106634
rect 501562 106398 501646 106634
rect 501882 106398 537326 106634
rect 537562 106398 537646 106634
rect 537882 106398 573326 106634
rect 573562 106398 573646 106634
rect 573882 106398 592062 106634
rect 592298 106398 592382 106634
rect 592618 106398 592650 106634
rect -8726 106366 592650 106398
rect -8726 102454 592650 102486
rect -8726 102218 -7734 102454
rect -7498 102218 -7414 102454
rect -7178 102218 28826 102454
rect 29062 102218 29146 102454
rect 29382 102218 244826 102454
rect 245062 102218 245146 102454
rect 245382 102218 280826 102454
rect 281062 102218 281146 102454
rect 281382 102218 352826 102454
rect 353062 102218 353146 102454
rect 353382 102218 388826 102454
rect 389062 102218 389146 102454
rect 389382 102218 424826 102454
rect 425062 102218 425146 102454
rect 425382 102218 460826 102454
rect 461062 102218 461146 102454
rect 461382 102218 496826 102454
rect 497062 102218 497146 102454
rect 497382 102218 532826 102454
rect 533062 102218 533146 102454
rect 533382 102218 568826 102454
rect 569062 102218 569146 102454
rect 569382 102218 591102 102454
rect 591338 102218 591422 102454
rect 591658 102218 592650 102454
rect -8726 102134 592650 102218
rect -8726 101898 -7734 102134
rect -7498 101898 -7414 102134
rect -7178 101898 28826 102134
rect 29062 101898 29146 102134
rect 29382 101898 244826 102134
rect 245062 101898 245146 102134
rect 245382 101898 280826 102134
rect 281062 101898 281146 102134
rect 281382 101898 352826 102134
rect 353062 101898 353146 102134
rect 353382 101898 388826 102134
rect 389062 101898 389146 102134
rect 389382 101898 424826 102134
rect 425062 101898 425146 102134
rect 425382 101898 460826 102134
rect 461062 101898 461146 102134
rect 461382 101898 496826 102134
rect 497062 101898 497146 102134
rect 497382 101898 532826 102134
rect 533062 101898 533146 102134
rect 533382 101898 568826 102134
rect 569062 101898 569146 102134
rect 569382 101898 591102 102134
rect 591338 101898 591422 102134
rect 591658 101898 592650 102134
rect -8726 101866 592650 101898
rect -8726 97954 592650 97986
rect -8726 97718 -6774 97954
rect -6538 97718 -6454 97954
rect -6218 97718 24326 97954
rect 24562 97718 24646 97954
rect 24882 97718 240326 97954
rect 240562 97718 240646 97954
rect 240882 97718 276326 97954
rect 276562 97718 276646 97954
rect 276882 97718 348326 97954
rect 348562 97718 348646 97954
rect 348882 97718 384326 97954
rect 384562 97718 384646 97954
rect 384882 97718 420326 97954
rect 420562 97718 420646 97954
rect 420882 97718 456326 97954
rect 456562 97718 456646 97954
rect 456882 97718 492326 97954
rect 492562 97718 492646 97954
rect 492882 97718 528326 97954
rect 528562 97718 528646 97954
rect 528882 97718 564326 97954
rect 564562 97718 564646 97954
rect 564882 97718 590142 97954
rect 590378 97718 590462 97954
rect 590698 97718 592650 97954
rect -8726 97634 592650 97718
rect -8726 97398 -6774 97634
rect -6538 97398 -6454 97634
rect -6218 97398 24326 97634
rect 24562 97398 24646 97634
rect 24882 97398 240326 97634
rect 240562 97398 240646 97634
rect 240882 97398 276326 97634
rect 276562 97398 276646 97634
rect 276882 97398 348326 97634
rect 348562 97398 348646 97634
rect 348882 97398 384326 97634
rect 384562 97398 384646 97634
rect 384882 97398 420326 97634
rect 420562 97398 420646 97634
rect 420882 97398 456326 97634
rect 456562 97398 456646 97634
rect 456882 97398 492326 97634
rect 492562 97398 492646 97634
rect 492882 97398 528326 97634
rect 528562 97398 528646 97634
rect 528882 97398 564326 97634
rect 564562 97398 564646 97634
rect 564882 97398 590142 97634
rect 590378 97398 590462 97634
rect 590698 97398 592650 97634
rect -8726 97366 592650 97398
rect -8726 93454 592650 93486
rect -8726 93218 -5814 93454
rect -5578 93218 -5494 93454
rect -5258 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 589182 93454
rect 589418 93218 589502 93454
rect 589738 93218 592650 93454
rect -8726 93134 592650 93218
rect -8726 92898 -5814 93134
rect -5578 92898 -5494 93134
rect -5258 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 589182 93134
rect 589418 92898 589502 93134
rect 589738 92898 592650 93134
rect -8726 92866 592650 92898
rect -8726 88954 592650 88986
rect -8726 88718 -4854 88954
rect -4618 88718 -4534 88954
rect -4298 88718 15326 88954
rect 15562 88718 15646 88954
rect 15882 88718 51326 88954
rect 51562 88718 51646 88954
rect 51882 88718 231326 88954
rect 231562 88718 231646 88954
rect 231882 88718 267326 88954
rect 267562 88718 267646 88954
rect 267882 88718 375326 88954
rect 375562 88718 375646 88954
rect 375882 88718 411326 88954
rect 411562 88718 411646 88954
rect 411882 88718 447326 88954
rect 447562 88718 447646 88954
rect 447882 88718 483326 88954
rect 483562 88718 483646 88954
rect 483882 88718 519326 88954
rect 519562 88718 519646 88954
rect 519882 88718 555326 88954
rect 555562 88718 555646 88954
rect 555882 88718 588222 88954
rect 588458 88718 588542 88954
rect 588778 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -4854 88634
rect -4618 88398 -4534 88634
rect -4298 88398 15326 88634
rect 15562 88398 15646 88634
rect 15882 88398 51326 88634
rect 51562 88398 51646 88634
rect 51882 88398 231326 88634
rect 231562 88398 231646 88634
rect 231882 88398 267326 88634
rect 267562 88398 267646 88634
rect 267882 88398 375326 88634
rect 375562 88398 375646 88634
rect 375882 88398 411326 88634
rect 411562 88398 411646 88634
rect 411882 88398 447326 88634
rect 447562 88398 447646 88634
rect 447882 88398 483326 88634
rect 483562 88398 483646 88634
rect 483882 88398 519326 88634
rect 519562 88398 519646 88634
rect 519882 88398 555326 88634
rect 555562 88398 555646 88634
rect 555882 88398 588222 88634
rect 588458 88398 588542 88634
rect 588778 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -3894 84454
rect -3658 84218 -3574 84454
rect -3338 84218 10826 84454
rect 11062 84218 11146 84454
rect 11382 84218 46826 84454
rect 47062 84218 47146 84454
rect 47382 84218 226826 84454
rect 227062 84218 227146 84454
rect 227382 84218 262826 84454
rect 263062 84218 263146 84454
rect 263382 84218 370826 84454
rect 371062 84218 371146 84454
rect 371382 84218 406826 84454
rect 407062 84218 407146 84454
rect 407382 84218 442826 84454
rect 443062 84218 443146 84454
rect 443382 84218 478826 84454
rect 479062 84218 479146 84454
rect 479382 84218 514826 84454
rect 515062 84218 515146 84454
rect 515382 84218 550826 84454
rect 551062 84218 551146 84454
rect 551382 84218 587262 84454
rect 587498 84218 587582 84454
rect 587818 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -3894 84134
rect -3658 83898 -3574 84134
rect -3338 83898 10826 84134
rect 11062 83898 11146 84134
rect 11382 83898 46826 84134
rect 47062 83898 47146 84134
rect 47382 83898 226826 84134
rect 227062 83898 227146 84134
rect 227382 83898 262826 84134
rect 263062 83898 263146 84134
rect 263382 83898 370826 84134
rect 371062 83898 371146 84134
rect 371382 83898 406826 84134
rect 407062 83898 407146 84134
rect 407382 83898 442826 84134
rect 443062 83898 443146 84134
rect 443382 83898 478826 84134
rect 479062 83898 479146 84134
rect 479382 83898 514826 84134
rect 515062 83898 515146 84134
rect 515382 83898 550826 84134
rect 551062 83898 551146 84134
rect 551382 83898 587262 84134
rect 587498 83898 587582 84134
rect 587818 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 79954 592650 79986
rect -8726 79718 -2934 79954
rect -2698 79718 -2614 79954
rect -2378 79718 6326 79954
rect 6562 79718 6646 79954
rect 6882 79718 42326 79954
rect 42562 79718 42646 79954
rect 42882 79718 79610 79954
rect 79846 79718 110330 79954
rect 110566 79718 141050 79954
rect 141286 79718 171770 79954
rect 172006 79718 202490 79954
rect 202726 79718 258326 79954
rect 258562 79718 258646 79954
rect 258882 79718 294326 79954
rect 294562 79718 294646 79954
rect 294882 79718 319610 79954
rect 319846 79718 366326 79954
rect 366562 79718 366646 79954
rect 366882 79718 402326 79954
rect 402562 79718 402646 79954
rect 402882 79718 438326 79954
rect 438562 79718 438646 79954
rect 438882 79718 474326 79954
rect 474562 79718 474646 79954
rect 474882 79718 510326 79954
rect 510562 79718 510646 79954
rect 510882 79718 546326 79954
rect 546562 79718 546646 79954
rect 546882 79718 582326 79954
rect 582562 79718 582646 79954
rect 582882 79718 586302 79954
rect 586538 79718 586622 79954
rect 586858 79718 592650 79954
rect -8726 79634 592650 79718
rect -8726 79398 -2934 79634
rect -2698 79398 -2614 79634
rect -2378 79398 6326 79634
rect 6562 79398 6646 79634
rect 6882 79398 42326 79634
rect 42562 79398 42646 79634
rect 42882 79398 79610 79634
rect 79846 79398 110330 79634
rect 110566 79398 141050 79634
rect 141286 79398 171770 79634
rect 172006 79398 202490 79634
rect 202726 79398 258326 79634
rect 258562 79398 258646 79634
rect 258882 79398 294326 79634
rect 294562 79398 294646 79634
rect 294882 79398 319610 79634
rect 319846 79398 366326 79634
rect 366562 79398 366646 79634
rect 366882 79398 402326 79634
rect 402562 79398 402646 79634
rect 402882 79398 438326 79634
rect 438562 79398 438646 79634
rect 438882 79398 474326 79634
rect 474562 79398 474646 79634
rect 474882 79398 510326 79634
rect 510562 79398 510646 79634
rect 510882 79398 546326 79634
rect 546562 79398 546646 79634
rect 546882 79398 582326 79634
rect 582562 79398 582646 79634
rect 582882 79398 586302 79634
rect 586538 79398 586622 79634
rect 586858 79398 592650 79634
rect -8726 79366 592650 79398
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 304250 75454
rect 304486 75218 334970 75454
rect 335206 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 304250 75134
rect 304486 74898 334970 75134
rect 335206 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 70954 592650 70986
rect -8726 70718 -8694 70954
rect -8458 70718 -8374 70954
rect -8138 70718 33326 70954
rect 33562 70718 33646 70954
rect 33882 70718 249326 70954
rect 249562 70718 249646 70954
rect 249882 70718 285326 70954
rect 285562 70718 285646 70954
rect 285882 70718 357326 70954
rect 357562 70718 357646 70954
rect 357882 70718 393326 70954
rect 393562 70718 393646 70954
rect 393882 70718 429326 70954
rect 429562 70718 429646 70954
rect 429882 70718 465326 70954
rect 465562 70718 465646 70954
rect 465882 70718 501326 70954
rect 501562 70718 501646 70954
rect 501882 70718 537326 70954
rect 537562 70718 537646 70954
rect 537882 70718 573326 70954
rect 573562 70718 573646 70954
rect 573882 70718 592062 70954
rect 592298 70718 592382 70954
rect 592618 70718 592650 70954
rect -8726 70634 592650 70718
rect -8726 70398 -8694 70634
rect -8458 70398 -8374 70634
rect -8138 70398 33326 70634
rect 33562 70398 33646 70634
rect 33882 70398 249326 70634
rect 249562 70398 249646 70634
rect 249882 70398 285326 70634
rect 285562 70398 285646 70634
rect 285882 70398 357326 70634
rect 357562 70398 357646 70634
rect 357882 70398 393326 70634
rect 393562 70398 393646 70634
rect 393882 70398 429326 70634
rect 429562 70398 429646 70634
rect 429882 70398 465326 70634
rect 465562 70398 465646 70634
rect 465882 70398 501326 70634
rect 501562 70398 501646 70634
rect 501882 70398 537326 70634
rect 537562 70398 537646 70634
rect 537882 70398 573326 70634
rect 573562 70398 573646 70634
rect 573882 70398 592062 70634
rect 592298 70398 592382 70634
rect 592618 70398 592650 70634
rect -8726 70366 592650 70398
rect -8726 66454 592650 66486
rect -8726 66218 -7734 66454
rect -7498 66218 -7414 66454
rect -7178 66218 28826 66454
rect 29062 66218 29146 66454
rect 29382 66218 244826 66454
rect 245062 66218 245146 66454
rect 245382 66218 280826 66454
rect 281062 66218 281146 66454
rect 281382 66218 352826 66454
rect 353062 66218 353146 66454
rect 353382 66218 388826 66454
rect 389062 66218 389146 66454
rect 389382 66218 424826 66454
rect 425062 66218 425146 66454
rect 425382 66218 460826 66454
rect 461062 66218 461146 66454
rect 461382 66218 496826 66454
rect 497062 66218 497146 66454
rect 497382 66218 532826 66454
rect 533062 66218 533146 66454
rect 533382 66218 568826 66454
rect 569062 66218 569146 66454
rect 569382 66218 591102 66454
rect 591338 66218 591422 66454
rect 591658 66218 592650 66454
rect -8726 66134 592650 66218
rect -8726 65898 -7734 66134
rect -7498 65898 -7414 66134
rect -7178 65898 28826 66134
rect 29062 65898 29146 66134
rect 29382 65898 244826 66134
rect 245062 65898 245146 66134
rect 245382 65898 280826 66134
rect 281062 65898 281146 66134
rect 281382 65898 352826 66134
rect 353062 65898 353146 66134
rect 353382 65898 388826 66134
rect 389062 65898 389146 66134
rect 389382 65898 424826 66134
rect 425062 65898 425146 66134
rect 425382 65898 460826 66134
rect 461062 65898 461146 66134
rect 461382 65898 496826 66134
rect 497062 65898 497146 66134
rect 497382 65898 532826 66134
rect 533062 65898 533146 66134
rect 533382 65898 568826 66134
rect 569062 65898 569146 66134
rect 569382 65898 591102 66134
rect 591338 65898 591422 66134
rect 591658 65898 592650 66134
rect -8726 65866 592650 65898
rect -8726 61954 592650 61986
rect -8726 61718 -6774 61954
rect -6538 61718 -6454 61954
rect -6218 61718 24326 61954
rect 24562 61718 24646 61954
rect 24882 61718 240326 61954
rect 240562 61718 240646 61954
rect 240882 61718 276326 61954
rect 276562 61718 276646 61954
rect 276882 61718 348326 61954
rect 348562 61718 348646 61954
rect 348882 61718 384326 61954
rect 384562 61718 384646 61954
rect 384882 61718 420326 61954
rect 420562 61718 420646 61954
rect 420882 61718 456326 61954
rect 456562 61718 456646 61954
rect 456882 61718 492326 61954
rect 492562 61718 492646 61954
rect 492882 61718 528326 61954
rect 528562 61718 528646 61954
rect 528882 61718 564326 61954
rect 564562 61718 564646 61954
rect 564882 61718 590142 61954
rect 590378 61718 590462 61954
rect 590698 61718 592650 61954
rect -8726 61634 592650 61718
rect -8726 61398 -6774 61634
rect -6538 61398 -6454 61634
rect -6218 61398 24326 61634
rect 24562 61398 24646 61634
rect 24882 61398 240326 61634
rect 240562 61398 240646 61634
rect 240882 61398 276326 61634
rect 276562 61398 276646 61634
rect 276882 61398 348326 61634
rect 348562 61398 348646 61634
rect 348882 61398 384326 61634
rect 384562 61398 384646 61634
rect 384882 61398 420326 61634
rect 420562 61398 420646 61634
rect 420882 61398 456326 61634
rect 456562 61398 456646 61634
rect 456882 61398 492326 61634
rect 492562 61398 492646 61634
rect 492882 61398 528326 61634
rect 528562 61398 528646 61634
rect 528882 61398 564326 61634
rect 564562 61398 564646 61634
rect 564882 61398 590142 61634
rect 590378 61398 590462 61634
rect 590698 61398 592650 61634
rect -8726 61366 592650 61398
rect -8726 57454 592650 57486
rect -8726 57218 -5814 57454
rect -5578 57218 -5494 57454
rect -5258 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 589182 57454
rect 589418 57218 589502 57454
rect 589738 57218 592650 57454
rect -8726 57134 592650 57218
rect -8726 56898 -5814 57134
rect -5578 56898 -5494 57134
rect -5258 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 589182 57134
rect 589418 56898 589502 57134
rect 589738 56898 592650 57134
rect -8726 56866 592650 56898
rect -8726 52954 592650 52986
rect -8726 52718 -4854 52954
rect -4618 52718 -4534 52954
rect -4298 52718 15326 52954
rect 15562 52718 15646 52954
rect 15882 52718 51326 52954
rect 51562 52718 51646 52954
rect 51882 52718 87326 52954
rect 87562 52718 87646 52954
rect 87882 52718 123326 52954
rect 123562 52718 123646 52954
rect 123882 52718 159326 52954
rect 159562 52718 159646 52954
rect 159882 52718 195326 52954
rect 195562 52718 195646 52954
rect 195882 52718 231326 52954
rect 231562 52718 231646 52954
rect 231882 52718 267326 52954
rect 267562 52718 267646 52954
rect 267882 52718 303326 52954
rect 303562 52718 303646 52954
rect 303882 52718 339326 52954
rect 339562 52718 339646 52954
rect 339882 52718 375326 52954
rect 375562 52718 375646 52954
rect 375882 52718 411326 52954
rect 411562 52718 411646 52954
rect 411882 52718 447326 52954
rect 447562 52718 447646 52954
rect 447882 52718 483326 52954
rect 483562 52718 483646 52954
rect 483882 52718 519326 52954
rect 519562 52718 519646 52954
rect 519882 52718 555326 52954
rect 555562 52718 555646 52954
rect 555882 52718 588222 52954
rect 588458 52718 588542 52954
rect 588778 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -4854 52634
rect -4618 52398 -4534 52634
rect -4298 52398 15326 52634
rect 15562 52398 15646 52634
rect 15882 52398 51326 52634
rect 51562 52398 51646 52634
rect 51882 52398 87326 52634
rect 87562 52398 87646 52634
rect 87882 52398 123326 52634
rect 123562 52398 123646 52634
rect 123882 52398 159326 52634
rect 159562 52398 159646 52634
rect 159882 52398 195326 52634
rect 195562 52398 195646 52634
rect 195882 52398 231326 52634
rect 231562 52398 231646 52634
rect 231882 52398 267326 52634
rect 267562 52398 267646 52634
rect 267882 52398 303326 52634
rect 303562 52398 303646 52634
rect 303882 52398 339326 52634
rect 339562 52398 339646 52634
rect 339882 52398 375326 52634
rect 375562 52398 375646 52634
rect 375882 52398 411326 52634
rect 411562 52398 411646 52634
rect 411882 52398 447326 52634
rect 447562 52398 447646 52634
rect 447882 52398 483326 52634
rect 483562 52398 483646 52634
rect 483882 52398 519326 52634
rect 519562 52398 519646 52634
rect 519882 52398 555326 52634
rect 555562 52398 555646 52634
rect 555882 52398 588222 52634
rect 588458 52398 588542 52634
rect 588778 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -3894 48454
rect -3658 48218 -3574 48454
rect -3338 48218 10826 48454
rect 11062 48218 11146 48454
rect 11382 48218 46826 48454
rect 47062 48218 47146 48454
rect 47382 48218 82826 48454
rect 83062 48218 83146 48454
rect 83382 48218 118826 48454
rect 119062 48218 119146 48454
rect 119382 48218 154826 48454
rect 155062 48218 155146 48454
rect 155382 48218 190826 48454
rect 191062 48218 191146 48454
rect 191382 48218 226826 48454
rect 227062 48218 227146 48454
rect 227382 48218 262826 48454
rect 263062 48218 263146 48454
rect 263382 48218 298826 48454
rect 299062 48218 299146 48454
rect 299382 48218 334826 48454
rect 335062 48218 335146 48454
rect 335382 48218 370826 48454
rect 371062 48218 371146 48454
rect 371382 48218 406826 48454
rect 407062 48218 407146 48454
rect 407382 48218 442826 48454
rect 443062 48218 443146 48454
rect 443382 48218 478826 48454
rect 479062 48218 479146 48454
rect 479382 48218 514826 48454
rect 515062 48218 515146 48454
rect 515382 48218 550826 48454
rect 551062 48218 551146 48454
rect 551382 48218 587262 48454
rect 587498 48218 587582 48454
rect 587818 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -3894 48134
rect -3658 47898 -3574 48134
rect -3338 47898 10826 48134
rect 11062 47898 11146 48134
rect 11382 47898 46826 48134
rect 47062 47898 47146 48134
rect 47382 47898 82826 48134
rect 83062 47898 83146 48134
rect 83382 47898 118826 48134
rect 119062 47898 119146 48134
rect 119382 47898 154826 48134
rect 155062 47898 155146 48134
rect 155382 47898 190826 48134
rect 191062 47898 191146 48134
rect 191382 47898 226826 48134
rect 227062 47898 227146 48134
rect 227382 47898 262826 48134
rect 263062 47898 263146 48134
rect 263382 47898 298826 48134
rect 299062 47898 299146 48134
rect 299382 47898 334826 48134
rect 335062 47898 335146 48134
rect 335382 47898 370826 48134
rect 371062 47898 371146 48134
rect 371382 47898 406826 48134
rect 407062 47898 407146 48134
rect 407382 47898 442826 48134
rect 443062 47898 443146 48134
rect 443382 47898 478826 48134
rect 479062 47898 479146 48134
rect 479382 47898 514826 48134
rect 515062 47898 515146 48134
rect 515382 47898 550826 48134
rect 551062 47898 551146 48134
rect 551382 47898 587262 48134
rect 587498 47898 587582 48134
rect 587818 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 43954 592650 43986
rect -8726 43718 -2934 43954
rect -2698 43718 -2614 43954
rect -2378 43718 6326 43954
rect 6562 43718 6646 43954
rect 6882 43718 42326 43954
rect 42562 43718 42646 43954
rect 42882 43718 78326 43954
rect 78562 43718 78646 43954
rect 78882 43718 114326 43954
rect 114562 43718 114646 43954
rect 114882 43718 150326 43954
rect 150562 43718 150646 43954
rect 150882 43718 186326 43954
rect 186562 43718 186646 43954
rect 186882 43718 222326 43954
rect 222562 43718 222646 43954
rect 222882 43718 258326 43954
rect 258562 43718 258646 43954
rect 258882 43718 294326 43954
rect 294562 43718 294646 43954
rect 294882 43718 330326 43954
rect 330562 43718 330646 43954
rect 330882 43718 366326 43954
rect 366562 43718 366646 43954
rect 366882 43718 402326 43954
rect 402562 43718 402646 43954
rect 402882 43718 438326 43954
rect 438562 43718 438646 43954
rect 438882 43718 474326 43954
rect 474562 43718 474646 43954
rect 474882 43718 510326 43954
rect 510562 43718 510646 43954
rect 510882 43718 546326 43954
rect 546562 43718 546646 43954
rect 546882 43718 582326 43954
rect 582562 43718 582646 43954
rect 582882 43718 586302 43954
rect 586538 43718 586622 43954
rect 586858 43718 592650 43954
rect -8726 43634 592650 43718
rect -8726 43398 -2934 43634
rect -2698 43398 -2614 43634
rect -2378 43398 6326 43634
rect 6562 43398 6646 43634
rect 6882 43398 42326 43634
rect 42562 43398 42646 43634
rect 42882 43398 78326 43634
rect 78562 43398 78646 43634
rect 78882 43398 114326 43634
rect 114562 43398 114646 43634
rect 114882 43398 150326 43634
rect 150562 43398 150646 43634
rect 150882 43398 186326 43634
rect 186562 43398 186646 43634
rect 186882 43398 222326 43634
rect 222562 43398 222646 43634
rect 222882 43398 258326 43634
rect 258562 43398 258646 43634
rect 258882 43398 294326 43634
rect 294562 43398 294646 43634
rect 294882 43398 330326 43634
rect 330562 43398 330646 43634
rect 330882 43398 366326 43634
rect 366562 43398 366646 43634
rect 366882 43398 402326 43634
rect 402562 43398 402646 43634
rect 402882 43398 438326 43634
rect 438562 43398 438646 43634
rect 438882 43398 474326 43634
rect 474562 43398 474646 43634
rect 474882 43398 510326 43634
rect 510562 43398 510646 43634
rect 510882 43398 546326 43634
rect 546562 43398 546646 43634
rect 546882 43398 582326 43634
rect 582562 43398 582646 43634
rect 582882 43398 586302 43634
rect 586538 43398 586622 43634
rect 586858 43398 592650 43634
rect -8726 43366 592650 43398
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 34954 592650 34986
rect -8726 34718 -8694 34954
rect -8458 34718 -8374 34954
rect -8138 34718 33326 34954
rect 33562 34718 33646 34954
rect 33882 34718 69326 34954
rect 69562 34718 69646 34954
rect 69882 34718 105326 34954
rect 105562 34718 105646 34954
rect 105882 34718 141326 34954
rect 141562 34718 141646 34954
rect 141882 34718 177326 34954
rect 177562 34718 177646 34954
rect 177882 34718 213326 34954
rect 213562 34718 213646 34954
rect 213882 34718 249326 34954
rect 249562 34718 249646 34954
rect 249882 34718 285326 34954
rect 285562 34718 285646 34954
rect 285882 34718 321326 34954
rect 321562 34718 321646 34954
rect 321882 34718 357326 34954
rect 357562 34718 357646 34954
rect 357882 34718 393326 34954
rect 393562 34718 393646 34954
rect 393882 34718 429326 34954
rect 429562 34718 429646 34954
rect 429882 34718 465326 34954
rect 465562 34718 465646 34954
rect 465882 34718 501326 34954
rect 501562 34718 501646 34954
rect 501882 34718 537326 34954
rect 537562 34718 537646 34954
rect 537882 34718 573326 34954
rect 573562 34718 573646 34954
rect 573882 34718 592062 34954
rect 592298 34718 592382 34954
rect 592618 34718 592650 34954
rect -8726 34634 592650 34718
rect -8726 34398 -8694 34634
rect -8458 34398 -8374 34634
rect -8138 34398 33326 34634
rect 33562 34398 33646 34634
rect 33882 34398 69326 34634
rect 69562 34398 69646 34634
rect 69882 34398 105326 34634
rect 105562 34398 105646 34634
rect 105882 34398 141326 34634
rect 141562 34398 141646 34634
rect 141882 34398 177326 34634
rect 177562 34398 177646 34634
rect 177882 34398 213326 34634
rect 213562 34398 213646 34634
rect 213882 34398 249326 34634
rect 249562 34398 249646 34634
rect 249882 34398 285326 34634
rect 285562 34398 285646 34634
rect 285882 34398 321326 34634
rect 321562 34398 321646 34634
rect 321882 34398 357326 34634
rect 357562 34398 357646 34634
rect 357882 34398 393326 34634
rect 393562 34398 393646 34634
rect 393882 34398 429326 34634
rect 429562 34398 429646 34634
rect 429882 34398 465326 34634
rect 465562 34398 465646 34634
rect 465882 34398 501326 34634
rect 501562 34398 501646 34634
rect 501882 34398 537326 34634
rect 537562 34398 537646 34634
rect 537882 34398 573326 34634
rect 573562 34398 573646 34634
rect 573882 34398 592062 34634
rect 592298 34398 592382 34634
rect 592618 34398 592650 34634
rect -8726 34366 592650 34398
rect -8726 30454 592650 30486
rect -8726 30218 -7734 30454
rect -7498 30218 -7414 30454
rect -7178 30218 28826 30454
rect 29062 30218 29146 30454
rect 29382 30218 64826 30454
rect 65062 30218 65146 30454
rect 65382 30218 100826 30454
rect 101062 30218 101146 30454
rect 101382 30218 136826 30454
rect 137062 30218 137146 30454
rect 137382 30218 172826 30454
rect 173062 30218 173146 30454
rect 173382 30218 208826 30454
rect 209062 30218 209146 30454
rect 209382 30218 244826 30454
rect 245062 30218 245146 30454
rect 245382 30218 280826 30454
rect 281062 30218 281146 30454
rect 281382 30218 316826 30454
rect 317062 30218 317146 30454
rect 317382 30218 352826 30454
rect 353062 30218 353146 30454
rect 353382 30218 388826 30454
rect 389062 30218 389146 30454
rect 389382 30218 424826 30454
rect 425062 30218 425146 30454
rect 425382 30218 460826 30454
rect 461062 30218 461146 30454
rect 461382 30218 496826 30454
rect 497062 30218 497146 30454
rect 497382 30218 532826 30454
rect 533062 30218 533146 30454
rect 533382 30218 568826 30454
rect 569062 30218 569146 30454
rect 569382 30218 591102 30454
rect 591338 30218 591422 30454
rect 591658 30218 592650 30454
rect -8726 30134 592650 30218
rect -8726 29898 -7734 30134
rect -7498 29898 -7414 30134
rect -7178 29898 28826 30134
rect 29062 29898 29146 30134
rect 29382 29898 64826 30134
rect 65062 29898 65146 30134
rect 65382 29898 100826 30134
rect 101062 29898 101146 30134
rect 101382 29898 136826 30134
rect 137062 29898 137146 30134
rect 137382 29898 172826 30134
rect 173062 29898 173146 30134
rect 173382 29898 208826 30134
rect 209062 29898 209146 30134
rect 209382 29898 244826 30134
rect 245062 29898 245146 30134
rect 245382 29898 280826 30134
rect 281062 29898 281146 30134
rect 281382 29898 316826 30134
rect 317062 29898 317146 30134
rect 317382 29898 352826 30134
rect 353062 29898 353146 30134
rect 353382 29898 388826 30134
rect 389062 29898 389146 30134
rect 389382 29898 424826 30134
rect 425062 29898 425146 30134
rect 425382 29898 460826 30134
rect 461062 29898 461146 30134
rect 461382 29898 496826 30134
rect 497062 29898 497146 30134
rect 497382 29898 532826 30134
rect 533062 29898 533146 30134
rect 533382 29898 568826 30134
rect 569062 29898 569146 30134
rect 569382 29898 591102 30134
rect 591338 29898 591422 30134
rect 591658 29898 592650 30134
rect -8726 29866 592650 29898
rect -8726 25954 592650 25986
rect -8726 25718 -6774 25954
rect -6538 25718 -6454 25954
rect -6218 25718 24326 25954
rect 24562 25718 24646 25954
rect 24882 25718 60326 25954
rect 60562 25718 60646 25954
rect 60882 25718 96326 25954
rect 96562 25718 96646 25954
rect 96882 25718 132326 25954
rect 132562 25718 132646 25954
rect 132882 25718 168326 25954
rect 168562 25718 168646 25954
rect 168882 25718 204326 25954
rect 204562 25718 204646 25954
rect 204882 25718 240326 25954
rect 240562 25718 240646 25954
rect 240882 25718 276326 25954
rect 276562 25718 276646 25954
rect 276882 25718 312326 25954
rect 312562 25718 312646 25954
rect 312882 25718 348326 25954
rect 348562 25718 348646 25954
rect 348882 25718 384326 25954
rect 384562 25718 384646 25954
rect 384882 25718 420326 25954
rect 420562 25718 420646 25954
rect 420882 25718 456326 25954
rect 456562 25718 456646 25954
rect 456882 25718 492326 25954
rect 492562 25718 492646 25954
rect 492882 25718 528326 25954
rect 528562 25718 528646 25954
rect 528882 25718 564326 25954
rect 564562 25718 564646 25954
rect 564882 25718 590142 25954
rect 590378 25718 590462 25954
rect 590698 25718 592650 25954
rect -8726 25634 592650 25718
rect -8726 25398 -6774 25634
rect -6538 25398 -6454 25634
rect -6218 25398 24326 25634
rect 24562 25398 24646 25634
rect 24882 25398 60326 25634
rect 60562 25398 60646 25634
rect 60882 25398 96326 25634
rect 96562 25398 96646 25634
rect 96882 25398 132326 25634
rect 132562 25398 132646 25634
rect 132882 25398 168326 25634
rect 168562 25398 168646 25634
rect 168882 25398 204326 25634
rect 204562 25398 204646 25634
rect 204882 25398 240326 25634
rect 240562 25398 240646 25634
rect 240882 25398 276326 25634
rect 276562 25398 276646 25634
rect 276882 25398 312326 25634
rect 312562 25398 312646 25634
rect 312882 25398 348326 25634
rect 348562 25398 348646 25634
rect 348882 25398 384326 25634
rect 384562 25398 384646 25634
rect 384882 25398 420326 25634
rect 420562 25398 420646 25634
rect 420882 25398 456326 25634
rect 456562 25398 456646 25634
rect 456882 25398 492326 25634
rect 492562 25398 492646 25634
rect 492882 25398 528326 25634
rect 528562 25398 528646 25634
rect 528882 25398 564326 25634
rect 564562 25398 564646 25634
rect 564882 25398 590142 25634
rect 590378 25398 590462 25634
rect 590698 25398 592650 25634
rect -8726 25366 592650 25398
rect -8726 21454 592650 21486
rect -8726 21218 -5814 21454
rect -5578 21218 -5494 21454
rect -5258 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 589182 21454
rect 589418 21218 589502 21454
rect 589738 21218 592650 21454
rect -8726 21134 592650 21218
rect -8726 20898 -5814 21134
rect -5578 20898 -5494 21134
rect -5258 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 589182 21134
rect 589418 20898 589502 21134
rect 589738 20898 592650 21134
rect -8726 20866 592650 20898
rect -8726 16954 592650 16986
rect -8726 16718 -4854 16954
rect -4618 16718 -4534 16954
rect -4298 16718 15326 16954
rect 15562 16718 15646 16954
rect 15882 16718 51326 16954
rect 51562 16718 51646 16954
rect 51882 16718 87326 16954
rect 87562 16718 87646 16954
rect 87882 16718 123326 16954
rect 123562 16718 123646 16954
rect 123882 16718 159326 16954
rect 159562 16718 159646 16954
rect 159882 16718 195326 16954
rect 195562 16718 195646 16954
rect 195882 16718 231326 16954
rect 231562 16718 231646 16954
rect 231882 16718 267326 16954
rect 267562 16718 267646 16954
rect 267882 16718 303326 16954
rect 303562 16718 303646 16954
rect 303882 16718 339326 16954
rect 339562 16718 339646 16954
rect 339882 16718 375326 16954
rect 375562 16718 375646 16954
rect 375882 16718 411326 16954
rect 411562 16718 411646 16954
rect 411882 16718 447326 16954
rect 447562 16718 447646 16954
rect 447882 16718 483326 16954
rect 483562 16718 483646 16954
rect 483882 16718 519326 16954
rect 519562 16718 519646 16954
rect 519882 16718 555326 16954
rect 555562 16718 555646 16954
rect 555882 16718 588222 16954
rect 588458 16718 588542 16954
rect 588778 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -4854 16634
rect -4618 16398 -4534 16634
rect -4298 16398 15326 16634
rect 15562 16398 15646 16634
rect 15882 16398 51326 16634
rect 51562 16398 51646 16634
rect 51882 16398 87326 16634
rect 87562 16398 87646 16634
rect 87882 16398 123326 16634
rect 123562 16398 123646 16634
rect 123882 16398 159326 16634
rect 159562 16398 159646 16634
rect 159882 16398 195326 16634
rect 195562 16398 195646 16634
rect 195882 16398 231326 16634
rect 231562 16398 231646 16634
rect 231882 16398 267326 16634
rect 267562 16398 267646 16634
rect 267882 16398 303326 16634
rect 303562 16398 303646 16634
rect 303882 16398 339326 16634
rect 339562 16398 339646 16634
rect 339882 16398 375326 16634
rect 375562 16398 375646 16634
rect 375882 16398 411326 16634
rect 411562 16398 411646 16634
rect 411882 16398 447326 16634
rect 447562 16398 447646 16634
rect 447882 16398 483326 16634
rect 483562 16398 483646 16634
rect 483882 16398 519326 16634
rect 519562 16398 519646 16634
rect 519882 16398 555326 16634
rect 555562 16398 555646 16634
rect 555882 16398 588222 16634
rect 588458 16398 588542 16634
rect 588778 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -3894 12454
rect -3658 12218 -3574 12454
rect -3338 12218 10826 12454
rect 11062 12218 11146 12454
rect 11382 12218 46826 12454
rect 47062 12218 47146 12454
rect 47382 12218 82826 12454
rect 83062 12218 83146 12454
rect 83382 12218 118826 12454
rect 119062 12218 119146 12454
rect 119382 12218 154826 12454
rect 155062 12218 155146 12454
rect 155382 12218 190826 12454
rect 191062 12218 191146 12454
rect 191382 12218 226826 12454
rect 227062 12218 227146 12454
rect 227382 12218 262826 12454
rect 263062 12218 263146 12454
rect 263382 12218 298826 12454
rect 299062 12218 299146 12454
rect 299382 12218 334826 12454
rect 335062 12218 335146 12454
rect 335382 12218 370826 12454
rect 371062 12218 371146 12454
rect 371382 12218 406826 12454
rect 407062 12218 407146 12454
rect 407382 12218 442826 12454
rect 443062 12218 443146 12454
rect 443382 12218 478826 12454
rect 479062 12218 479146 12454
rect 479382 12218 514826 12454
rect 515062 12218 515146 12454
rect 515382 12218 550826 12454
rect 551062 12218 551146 12454
rect 551382 12218 587262 12454
rect 587498 12218 587582 12454
rect 587818 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -3894 12134
rect -3658 11898 -3574 12134
rect -3338 11898 10826 12134
rect 11062 11898 11146 12134
rect 11382 11898 46826 12134
rect 47062 11898 47146 12134
rect 47382 11898 82826 12134
rect 83062 11898 83146 12134
rect 83382 11898 118826 12134
rect 119062 11898 119146 12134
rect 119382 11898 154826 12134
rect 155062 11898 155146 12134
rect 155382 11898 190826 12134
rect 191062 11898 191146 12134
rect 191382 11898 226826 12134
rect 227062 11898 227146 12134
rect 227382 11898 262826 12134
rect 263062 11898 263146 12134
rect 263382 11898 298826 12134
rect 299062 11898 299146 12134
rect 299382 11898 334826 12134
rect 335062 11898 335146 12134
rect 335382 11898 370826 12134
rect 371062 11898 371146 12134
rect 371382 11898 406826 12134
rect 407062 11898 407146 12134
rect 407382 11898 442826 12134
rect 443062 11898 443146 12134
rect 443382 11898 478826 12134
rect 479062 11898 479146 12134
rect 479382 11898 514826 12134
rect 515062 11898 515146 12134
rect 515382 11898 550826 12134
rect 551062 11898 551146 12134
rect 551382 11898 587262 12134
rect 587498 11898 587582 12134
rect 587818 11898 592650 12134
rect -8726 11866 592650 11898
rect -8726 7954 592650 7986
rect -8726 7718 -2934 7954
rect -2698 7718 -2614 7954
rect -2378 7718 6326 7954
rect 6562 7718 6646 7954
rect 6882 7718 42326 7954
rect 42562 7718 42646 7954
rect 42882 7718 78326 7954
rect 78562 7718 78646 7954
rect 78882 7718 114326 7954
rect 114562 7718 114646 7954
rect 114882 7718 150326 7954
rect 150562 7718 150646 7954
rect 150882 7718 186326 7954
rect 186562 7718 186646 7954
rect 186882 7718 222326 7954
rect 222562 7718 222646 7954
rect 222882 7718 258326 7954
rect 258562 7718 258646 7954
rect 258882 7718 294326 7954
rect 294562 7718 294646 7954
rect 294882 7718 330326 7954
rect 330562 7718 330646 7954
rect 330882 7718 366326 7954
rect 366562 7718 366646 7954
rect 366882 7718 402326 7954
rect 402562 7718 402646 7954
rect 402882 7718 438326 7954
rect 438562 7718 438646 7954
rect 438882 7718 474326 7954
rect 474562 7718 474646 7954
rect 474882 7718 510326 7954
rect 510562 7718 510646 7954
rect 510882 7718 546326 7954
rect 546562 7718 546646 7954
rect 546882 7718 582326 7954
rect 582562 7718 582646 7954
rect 582882 7718 586302 7954
rect 586538 7718 586622 7954
rect 586858 7718 592650 7954
rect -8726 7634 592650 7718
rect -8726 7398 -2934 7634
rect -2698 7398 -2614 7634
rect -2378 7398 6326 7634
rect 6562 7398 6646 7634
rect 6882 7398 42326 7634
rect 42562 7398 42646 7634
rect 42882 7398 78326 7634
rect 78562 7398 78646 7634
rect 78882 7398 114326 7634
rect 114562 7398 114646 7634
rect 114882 7398 150326 7634
rect 150562 7398 150646 7634
rect 150882 7398 186326 7634
rect 186562 7398 186646 7634
rect 186882 7398 222326 7634
rect 222562 7398 222646 7634
rect 222882 7398 258326 7634
rect 258562 7398 258646 7634
rect 258882 7398 294326 7634
rect 294562 7398 294646 7634
rect 294882 7398 330326 7634
rect 330562 7398 330646 7634
rect 330882 7398 366326 7634
rect 366562 7398 366646 7634
rect 366882 7398 402326 7634
rect 402562 7398 402646 7634
rect 402882 7398 438326 7634
rect 438562 7398 438646 7634
rect 438882 7398 474326 7634
rect 474562 7398 474646 7634
rect 474882 7398 510326 7634
rect 510562 7398 510646 7634
rect 510882 7398 546326 7634
rect 546562 7398 546646 7634
rect 546882 7398 582326 7634
rect 582562 7398 582646 7634
rect 582882 7398 586302 7634
rect 586538 7398 586622 7634
rect 586858 7398 592650 7634
rect -8726 7366 592650 7398
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 6326 -1306
rect 6562 -1542 6646 -1306
rect 6882 -1542 42326 -1306
rect 42562 -1542 42646 -1306
rect 42882 -1542 78326 -1306
rect 78562 -1542 78646 -1306
rect 78882 -1542 114326 -1306
rect 114562 -1542 114646 -1306
rect 114882 -1542 150326 -1306
rect 150562 -1542 150646 -1306
rect 150882 -1542 186326 -1306
rect 186562 -1542 186646 -1306
rect 186882 -1542 222326 -1306
rect 222562 -1542 222646 -1306
rect 222882 -1542 258326 -1306
rect 258562 -1542 258646 -1306
rect 258882 -1542 294326 -1306
rect 294562 -1542 294646 -1306
rect 294882 -1542 330326 -1306
rect 330562 -1542 330646 -1306
rect 330882 -1542 366326 -1306
rect 366562 -1542 366646 -1306
rect 366882 -1542 402326 -1306
rect 402562 -1542 402646 -1306
rect 402882 -1542 438326 -1306
rect 438562 -1542 438646 -1306
rect 438882 -1542 474326 -1306
rect 474562 -1542 474646 -1306
rect 474882 -1542 510326 -1306
rect 510562 -1542 510646 -1306
rect 510882 -1542 546326 -1306
rect 546562 -1542 546646 -1306
rect 546882 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 6326 -1626
rect 6562 -1862 6646 -1626
rect 6882 -1862 42326 -1626
rect 42562 -1862 42646 -1626
rect 42882 -1862 78326 -1626
rect 78562 -1862 78646 -1626
rect 78882 -1862 114326 -1626
rect 114562 -1862 114646 -1626
rect 114882 -1862 150326 -1626
rect 150562 -1862 150646 -1626
rect 150882 -1862 186326 -1626
rect 186562 -1862 186646 -1626
rect 186882 -1862 222326 -1626
rect 222562 -1862 222646 -1626
rect 222882 -1862 258326 -1626
rect 258562 -1862 258646 -1626
rect 258882 -1862 294326 -1626
rect 294562 -1862 294646 -1626
rect 294882 -1862 330326 -1626
rect 330562 -1862 330646 -1626
rect 330882 -1862 366326 -1626
rect 366562 -1862 366646 -1626
rect 366882 -1862 402326 -1626
rect 402562 -1862 402646 -1626
rect 402882 -1862 438326 -1626
rect 438562 -1862 438646 -1626
rect 438882 -1862 474326 -1626
rect 474562 -1862 474646 -1626
rect 474882 -1862 510326 -1626
rect 510562 -1862 510646 -1626
rect 510882 -1862 546326 -1626
rect 546562 -1862 546646 -1626
rect 546882 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 10826 -2266
rect 11062 -2502 11146 -2266
rect 11382 -2502 46826 -2266
rect 47062 -2502 47146 -2266
rect 47382 -2502 82826 -2266
rect 83062 -2502 83146 -2266
rect 83382 -2502 118826 -2266
rect 119062 -2502 119146 -2266
rect 119382 -2502 154826 -2266
rect 155062 -2502 155146 -2266
rect 155382 -2502 190826 -2266
rect 191062 -2502 191146 -2266
rect 191382 -2502 226826 -2266
rect 227062 -2502 227146 -2266
rect 227382 -2502 262826 -2266
rect 263062 -2502 263146 -2266
rect 263382 -2502 298826 -2266
rect 299062 -2502 299146 -2266
rect 299382 -2502 334826 -2266
rect 335062 -2502 335146 -2266
rect 335382 -2502 370826 -2266
rect 371062 -2502 371146 -2266
rect 371382 -2502 406826 -2266
rect 407062 -2502 407146 -2266
rect 407382 -2502 442826 -2266
rect 443062 -2502 443146 -2266
rect 443382 -2502 478826 -2266
rect 479062 -2502 479146 -2266
rect 479382 -2502 514826 -2266
rect 515062 -2502 515146 -2266
rect 515382 -2502 550826 -2266
rect 551062 -2502 551146 -2266
rect 551382 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 10826 -2586
rect 11062 -2822 11146 -2586
rect 11382 -2822 46826 -2586
rect 47062 -2822 47146 -2586
rect 47382 -2822 82826 -2586
rect 83062 -2822 83146 -2586
rect 83382 -2822 118826 -2586
rect 119062 -2822 119146 -2586
rect 119382 -2822 154826 -2586
rect 155062 -2822 155146 -2586
rect 155382 -2822 190826 -2586
rect 191062 -2822 191146 -2586
rect 191382 -2822 226826 -2586
rect 227062 -2822 227146 -2586
rect 227382 -2822 262826 -2586
rect 263062 -2822 263146 -2586
rect 263382 -2822 298826 -2586
rect 299062 -2822 299146 -2586
rect 299382 -2822 334826 -2586
rect 335062 -2822 335146 -2586
rect 335382 -2822 370826 -2586
rect 371062 -2822 371146 -2586
rect 371382 -2822 406826 -2586
rect 407062 -2822 407146 -2586
rect 407382 -2822 442826 -2586
rect 443062 -2822 443146 -2586
rect 443382 -2822 478826 -2586
rect 479062 -2822 479146 -2586
rect 479382 -2822 514826 -2586
rect 515062 -2822 515146 -2586
rect 515382 -2822 550826 -2586
rect 551062 -2822 551146 -2586
rect 551382 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 15326 -3226
rect 15562 -3462 15646 -3226
rect 15882 -3462 51326 -3226
rect 51562 -3462 51646 -3226
rect 51882 -3462 87326 -3226
rect 87562 -3462 87646 -3226
rect 87882 -3462 123326 -3226
rect 123562 -3462 123646 -3226
rect 123882 -3462 159326 -3226
rect 159562 -3462 159646 -3226
rect 159882 -3462 195326 -3226
rect 195562 -3462 195646 -3226
rect 195882 -3462 231326 -3226
rect 231562 -3462 231646 -3226
rect 231882 -3462 267326 -3226
rect 267562 -3462 267646 -3226
rect 267882 -3462 303326 -3226
rect 303562 -3462 303646 -3226
rect 303882 -3462 339326 -3226
rect 339562 -3462 339646 -3226
rect 339882 -3462 375326 -3226
rect 375562 -3462 375646 -3226
rect 375882 -3462 411326 -3226
rect 411562 -3462 411646 -3226
rect 411882 -3462 447326 -3226
rect 447562 -3462 447646 -3226
rect 447882 -3462 483326 -3226
rect 483562 -3462 483646 -3226
rect 483882 -3462 519326 -3226
rect 519562 -3462 519646 -3226
rect 519882 -3462 555326 -3226
rect 555562 -3462 555646 -3226
rect 555882 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 15326 -3546
rect 15562 -3782 15646 -3546
rect 15882 -3782 51326 -3546
rect 51562 -3782 51646 -3546
rect 51882 -3782 87326 -3546
rect 87562 -3782 87646 -3546
rect 87882 -3782 123326 -3546
rect 123562 -3782 123646 -3546
rect 123882 -3782 159326 -3546
rect 159562 -3782 159646 -3546
rect 159882 -3782 195326 -3546
rect 195562 -3782 195646 -3546
rect 195882 -3782 231326 -3546
rect 231562 -3782 231646 -3546
rect 231882 -3782 267326 -3546
rect 267562 -3782 267646 -3546
rect 267882 -3782 303326 -3546
rect 303562 -3782 303646 -3546
rect 303882 -3782 339326 -3546
rect 339562 -3782 339646 -3546
rect 339882 -3782 375326 -3546
rect 375562 -3782 375646 -3546
rect 375882 -3782 411326 -3546
rect 411562 -3782 411646 -3546
rect 411882 -3782 447326 -3546
rect 447562 -3782 447646 -3546
rect 447882 -3782 483326 -3546
rect 483562 -3782 483646 -3546
rect 483882 -3782 519326 -3546
rect 519562 -3782 519646 -3546
rect 519882 -3782 555326 -3546
rect 555562 -3782 555646 -3546
rect 555882 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 19826 -4186
rect 20062 -4422 20146 -4186
rect 20382 -4422 55826 -4186
rect 56062 -4422 56146 -4186
rect 56382 -4422 91826 -4186
rect 92062 -4422 92146 -4186
rect 92382 -4422 127826 -4186
rect 128062 -4422 128146 -4186
rect 128382 -4422 163826 -4186
rect 164062 -4422 164146 -4186
rect 164382 -4422 199826 -4186
rect 200062 -4422 200146 -4186
rect 200382 -4422 235826 -4186
rect 236062 -4422 236146 -4186
rect 236382 -4422 271826 -4186
rect 272062 -4422 272146 -4186
rect 272382 -4422 307826 -4186
rect 308062 -4422 308146 -4186
rect 308382 -4422 343826 -4186
rect 344062 -4422 344146 -4186
rect 344382 -4422 379826 -4186
rect 380062 -4422 380146 -4186
rect 380382 -4422 415826 -4186
rect 416062 -4422 416146 -4186
rect 416382 -4422 451826 -4186
rect 452062 -4422 452146 -4186
rect 452382 -4422 487826 -4186
rect 488062 -4422 488146 -4186
rect 488382 -4422 523826 -4186
rect 524062 -4422 524146 -4186
rect 524382 -4422 559826 -4186
rect 560062 -4422 560146 -4186
rect 560382 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 19826 -4506
rect 20062 -4742 20146 -4506
rect 20382 -4742 55826 -4506
rect 56062 -4742 56146 -4506
rect 56382 -4742 91826 -4506
rect 92062 -4742 92146 -4506
rect 92382 -4742 127826 -4506
rect 128062 -4742 128146 -4506
rect 128382 -4742 163826 -4506
rect 164062 -4742 164146 -4506
rect 164382 -4742 199826 -4506
rect 200062 -4742 200146 -4506
rect 200382 -4742 235826 -4506
rect 236062 -4742 236146 -4506
rect 236382 -4742 271826 -4506
rect 272062 -4742 272146 -4506
rect 272382 -4742 307826 -4506
rect 308062 -4742 308146 -4506
rect 308382 -4742 343826 -4506
rect 344062 -4742 344146 -4506
rect 344382 -4742 379826 -4506
rect 380062 -4742 380146 -4506
rect 380382 -4742 415826 -4506
rect 416062 -4742 416146 -4506
rect 416382 -4742 451826 -4506
rect 452062 -4742 452146 -4506
rect 452382 -4742 487826 -4506
rect 488062 -4742 488146 -4506
rect 488382 -4742 523826 -4506
rect 524062 -4742 524146 -4506
rect 524382 -4742 559826 -4506
rect 560062 -4742 560146 -4506
rect 560382 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 24326 -5146
rect 24562 -5382 24646 -5146
rect 24882 -5382 60326 -5146
rect 60562 -5382 60646 -5146
rect 60882 -5382 96326 -5146
rect 96562 -5382 96646 -5146
rect 96882 -5382 132326 -5146
rect 132562 -5382 132646 -5146
rect 132882 -5382 168326 -5146
rect 168562 -5382 168646 -5146
rect 168882 -5382 204326 -5146
rect 204562 -5382 204646 -5146
rect 204882 -5382 240326 -5146
rect 240562 -5382 240646 -5146
rect 240882 -5382 276326 -5146
rect 276562 -5382 276646 -5146
rect 276882 -5382 312326 -5146
rect 312562 -5382 312646 -5146
rect 312882 -5382 348326 -5146
rect 348562 -5382 348646 -5146
rect 348882 -5382 384326 -5146
rect 384562 -5382 384646 -5146
rect 384882 -5382 420326 -5146
rect 420562 -5382 420646 -5146
rect 420882 -5382 456326 -5146
rect 456562 -5382 456646 -5146
rect 456882 -5382 492326 -5146
rect 492562 -5382 492646 -5146
rect 492882 -5382 528326 -5146
rect 528562 -5382 528646 -5146
rect 528882 -5382 564326 -5146
rect 564562 -5382 564646 -5146
rect 564882 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 24326 -5466
rect 24562 -5702 24646 -5466
rect 24882 -5702 60326 -5466
rect 60562 -5702 60646 -5466
rect 60882 -5702 96326 -5466
rect 96562 -5702 96646 -5466
rect 96882 -5702 132326 -5466
rect 132562 -5702 132646 -5466
rect 132882 -5702 168326 -5466
rect 168562 -5702 168646 -5466
rect 168882 -5702 204326 -5466
rect 204562 -5702 204646 -5466
rect 204882 -5702 240326 -5466
rect 240562 -5702 240646 -5466
rect 240882 -5702 276326 -5466
rect 276562 -5702 276646 -5466
rect 276882 -5702 312326 -5466
rect 312562 -5702 312646 -5466
rect 312882 -5702 348326 -5466
rect 348562 -5702 348646 -5466
rect 348882 -5702 384326 -5466
rect 384562 -5702 384646 -5466
rect 384882 -5702 420326 -5466
rect 420562 -5702 420646 -5466
rect 420882 -5702 456326 -5466
rect 456562 -5702 456646 -5466
rect 456882 -5702 492326 -5466
rect 492562 -5702 492646 -5466
rect 492882 -5702 528326 -5466
rect 528562 -5702 528646 -5466
rect 528882 -5702 564326 -5466
rect 564562 -5702 564646 -5466
rect 564882 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 28826 -6106
rect 29062 -6342 29146 -6106
rect 29382 -6342 64826 -6106
rect 65062 -6342 65146 -6106
rect 65382 -6342 100826 -6106
rect 101062 -6342 101146 -6106
rect 101382 -6342 136826 -6106
rect 137062 -6342 137146 -6106
rect 137382 -6342 172826 -6106
rect 173062 -6342 173146 -6106
rect 173382 -6342 208826 -6106
rect 209062 -6342 209146 -6106
rect 209382 -6342 244826 -6106
rect 245062 -6342 245146 -6106
rect 245382 -6342 280826 -6106
rect 281062 -6342 281146 -6106
rect 281382 -6342 316826 -6106
rect 317062 -6342 317146 -6106
rect 317382 -6342 352826 -6106
rect 353062 -6342 353146 -6106
rect 353382 -6342 388826 -6106
rect 389062 -6342 389146 -6106
rect 389382 -6342 424826 -6106
rect 425062 -6342 425146 -6106
rect 425382 -6342 460826 -6106
rect 461062 -6342 461146 -6106
rect 461382 -6342 496826 -6106
rect 497062 -6342 497146 -6106
rect 497382 -6342 532826 -6106
rect 533062 -6342 533146 -6106
rect 533382 -6342 568826 -6106
rect 569062 -6342 569146 -6106
rect 569382 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 28826 -6426
rect 29062 -6662 29146 -6426
rect 29382 -6662 64826 -6426
rect 65062 -6662 65146 -6426
rect 65382 -6662 100826 -6426
rect 101062 -6662 101146 -6426
rect 101382 -6662 136826 -6426
rect 137062 -6662 137146 -6426
rect 137382 -6662 172826 -6426
rect 173062 -6662 173146 -6426
rect 173382 -6662 208826 -6426
rect 209062 -6662 209146 -6426
rect 209382 -6662 244826 -6426
rect 245062 -6662 245146 -6426
rect 245382 -6662 280826 -6426
rect 281062 -6662 281146 -6426
rect 281382 -6662 316826 -6426
rect 317062 -6662 317146 -6426
rect 317382 -6662 352826 -6426
rect 353062 -6662 353146 -6426
rect 353382 -6662 388826 -6426
rect 389062 -6662 389146 -6426
rect 389382 -6662 424826 -6426
rect 425062 -6662 425146 -6426
rect 425382 -6662 460826 -6426
rect 461062 -6662 461146 -6426
rect 461382 -6662 496826 -6426
rect 497062 -6662 497146 -6426
rect 497382 -6662 532826 -6426
rect 533062 -6662 533146 -6426
rect 533382 -6662 568826 -6426
rect 569062 -6662 569146 -6426
rect 569382 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 33326 -7066
rect 33562 -7302 33646 -7066
rect 33882 -7302 69326 -7066
rect 69562 -7302 69646 -7066
rect 69882 -7302 105326 -7066
rect 105562 -7302 105646 -7066
rect 105882 -7302 141326 -7066
rect 141562 -7302 141646 -7066
rect 141882 -7302 177326 -7066
rect 177562 -7302 177646 -7066
rect 177882 -7302 213326 -7066
rect 213562 -7302 213646 -7066
rect 213882 -7302 249326 -7066
rect 249562 -7302 249646 -7066
rect 249882 -7302 285326 -7066
rect 285562 -7302 285646 -7066
rect 285882 -7302 321326 -7066
rect 321562 -7302 321646 -7066
rect 321882 -7302 357326 -7066
rect 357562 -7302 357646 -7066
rect 357882 -7302 393326 -7066
rect 393562 -7302 393646 -7066
rect 393882 -7302 429326 -7066
rect 429562 -7302 429646 -7066
rect 429882 -7302 465326 -7066
rect 465562 -7302 465646 -7066
rect 465882 -7302 501326 -7066
rect 501562 -7302 501646 -7066
rect 501882 -7302 537326 -7066
rect 537562 -7302 537646 -7066
rect 537882 -7302 573326 -7066
rect 573562 -7302 573646 -7066
rect 573882 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 33326 -7386
rect 33562 -7622 33646 -7386
rect 33882 -7622 69326 -7386
rect 69562 -7622 69646 -7386
rect 69882 -7622 105326 -7386
rect 105562 -7622 105646 -7386
rect 105882 -7622 141326 -7386
rect 141562 -7622 141646 -7386
rect 141882 -7622 177326 -7386
rect 177562 -7622 177646 -7386
rect 177882 -7622 213326 -7386
rect 213562 -7622 213646 -7386
rect 213882 -7622 249326 -7386
rect 249562 -7622 249646 -7386
rect 249882 -7622 285326 -7386
rect 285562 -7622 285646 -7386
rect 285882 -7622 321326 -7386
rect 321562 -7622 321646 -7386
rect 321882 -7622 357326 -7386
rect 357562 -7622 357646 -7386
rect 357882 -7622 393326 -7386
rect 393562 -7622 393646 -7386
rect 393882 -7622 429326 -7386
rect 429562 -7622 429646 -7386
rect 429882 -7622 465326 -7386
rect 465562 -7622 465646 -7386
rect 465882 -7622 501326 -7386
rect 501562 -7622 501646 -7386
rect 501882 -7622 537326 -7386
rect 537562 -7622 537646 -7386
rect 537882 -7622 573326 -7386
rect 573562 -7622 573646 -7386
rect 573882 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use clk_div  top_cw.clk_div
timestamp 0
transform 1 0 480000 0 1 600000
box 0 0 40000 40000
use top_cw_logic  top_cw.top_cw_logic
timestamp 0
transform 1 0 360000 0 1 500000
box 0 0 40000 50000
use core  top_cw.upc.core
timestamp 0
transform 1 0 300000 0 1 60000
box 0 2048 40000 160000
use dcache  top_cw.upc.dcache
timestamp 0
transform 1 0 52000 0 1 280000
box 0 2128 200000 379760
use icache  top_cw.upc.icache
timestamp 0
transform 1 0 60000 0 1 60000
box 0 2042 160000 157808
use upper_core_logic  top_cw.upc.upper_core_logic
timestamp 0
transform 1 0 300000 0 1 280000
box 0 0 50000 50000
use wishbone_arbiter  top_cw.upc.wb_arbiter
timestamp 0
transform 1 0 280000 0 1 500000
box 1066 0 40000 40000
use wb_compressor  top_cw.wb_compressor
timestamp 0
transform 1 0 280000 0 1 600000
box 0 0 39362 40000
use wb_cross_clk  top_cw.wb_cross_clk
timestamp 0
transform 1 0 360000 0 1 600000
box 1066 0 38862 40000
use uprj_w_const  uprj_w_const
timestamp 0
transform 1 0 480000 0 1 500000
box 0 0 40000 40000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 664000 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 664000 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 664000 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 664000 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 664000 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 278000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 664000 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 542000 290414 598000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 642000 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 58000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 332000 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 642000 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 642000 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 498000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 542000 506414 598000 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 642000 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 10794 -7654 11414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46794 -7654 47414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 -7654 83414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 222000 83414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 82794 664000 83414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 -7654 119414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 222000 119414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 118794 664000 119414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 -7654 155414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 222000 155414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 154794 664000 155414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 -7654 191414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 222000 191414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 190794 664000 191414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 -7654 227414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 226794 664000 227414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 262794 -7654 263414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 -7654 299414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 222000 299414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 332000 299414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 542000 299414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 298794 642000 299414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 -7654 335414 58000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 222000 335414 278000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 334794 332000 335414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 -7654 371414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 552000 371414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 370794 642000 371414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 406794 -7654 407414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 442794 -7654 443414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 -7654 479414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 542000 479414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 478794 642000 479414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 -7654 515414 498000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 542000 515414 598000 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 514794 642000 515414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 550794 -7654 551414 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 19794 -7654 20414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 -7654 56414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 222000 56414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 55794 664000 56414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 -7654 92414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 222000 92414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91794 664000 92414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 -7654 128414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 222000 128414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 127794 664000 128414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 -7654 164414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 222000 164414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 163794 664000 164414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 -7654 200414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 222000 200414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 199794 664000 200414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 -7654 236414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 235794 664000 236414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 271794 -7654 272414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 -7654 308414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 222000 308414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 332000 308414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 542000 308414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 307794 642000 308414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 -7654 344414 58000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 222000 344414 278000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 343794 332000 344414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 -7654 380414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 552000 380414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 379794 642000 380414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 415794 -7654 416414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 451794 -7654 452414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 -7654 488414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 542000 488414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 487794 642000 488414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 -7654 524414 498000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 542000 524414 598000 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 523794 642000 524414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 559794 -7654 560414 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 20866 592650 21486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 56866 592650 57486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 92866 592650 93486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 128866 592650 129486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 164866 592650 165486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 200866 592650 201486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 236866 592650 237486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 272866 592650 273486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 308866 592650 309486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 344866 592650 345486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 380866 592650 381486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 416866 592650 417486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 452866 592650 453486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 488866 592650 489486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 524866 592650 525486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 560866 592650 561486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 596866 592650 597486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 632866 592650 633486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 668866 592650 669486 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 28794 -7654 29414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 -7654 65414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 64794 664000 65414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 -7654 101414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 100794 664000 101414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 -7654 137414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 136794 664000 137414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 -7654 173414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172794 664000 173414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 -7654 209414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 208794 664000 209414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 -7654 245414 278000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 244794 664000 245414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 -7654 281414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 280794 642000 281414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 -7654 317414 58000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 332000 317414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 316794 642000 317414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 -7654 353414 278000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 352794 332000 353414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 -7654 389414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 388794 642000 389414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 424794 -7654 425414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 460794 -7654 461414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 -7654 497414 498000 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 496794 642000 497414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 532794 -7654 533414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 568794 -7654 569414 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 29866 592650 30486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 65866 592650 66486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 101866 592650 102486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 137866 592650 138486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 173866 592650 174486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 209866 592650 210486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 245866 592650 246486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 281866 592650 282486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 317866 592650 318486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 353866 592650 354486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 389866 592650 390486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 425866 592650 426486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 461866 592650 462486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 497866 592650 498486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 533866 592650 534486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 569866 592650 570486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 605866 592650 606486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 641866 592650 642486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 677866 592650 678486 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 24294 -7654 24914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 -7654 60914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 222000 60914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 60294 664000 60914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 -7654 96914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 222000 96914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 96294 664000 96914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 -7654 132914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 222000 132914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 132294 664000 132914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 -7654 168914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 222000 168914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 168294 664000 168914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 -7654 204914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 222000 204914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 204294 664000 204914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 -7654 240914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 240294 664000 240914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 -7654 276914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 276294 642000 276914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 -7654 312914 58000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 222000 312914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 332000 312914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 312294 642000 312914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 -7654 348914 278000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 348294 332000 348914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 -7654 384914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 384294 642000 384914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 420294 -7654 420914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 456294 -7654 456914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 -7654 492914 498000 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 492294 642000 492914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 528294 -7654 528914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 564294 -7654 564914 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 25366 592650 25986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 61366 592650 61986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 97366 592650 97986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 133366 592650 133986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 169366 592650 169986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 205366 592650 205986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 241366 592650 241986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 277366 592650 277986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 313366 592650 313986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 349366 592650 349986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 385366 592650 385986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 421366 592650 421986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 457366 592650 457986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 493366 592650 493986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 529366 592650 529986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 565366 592650 565986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 601366 592650 601986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 637366 592650 637986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 673366 592650 673986 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 33294 -7654 33914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 -7654 69914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 69294 664000 69914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 -7654 105914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 105294 664000 105914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 -7654 141914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 141294 664000 141914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 -7654 177914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 177294 664000 177914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 -7654 213914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213294 664000 213914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 -7654 249914 278000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 249294 664000 249914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 -7654 285914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 285294 642000 285914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 -7654 321914 58000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 332000 321914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 321294 642000 321914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 -7654 357914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 357294 642000 357914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 -7654 393914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 393294 642000 393914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 429294 -7654 429914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 465294 -7654 465914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 -7654 501914 498000 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 501294 642000 501914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 537294 -7654 537914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 573294 -7654 573914 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 34366 592650 34986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 70366 592650 70986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 106366 592650 106986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 142366 592650 142986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 178366 592650 178986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 214366 592650 214986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 250366 592650 250986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 286366 592650 286986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 322366 592650 322986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 358366 592650 358986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 394366 592650 394986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 430366 592650 430986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 466366 592650 466986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 502366 592650 502986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 538366 592650 538986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 574366 592650 574986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 610366 592650 610986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 646366 592650 646986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 682366 592650 682986 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 6294 -7654 6914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42294 -7654 42914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 -7654 78914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 222000 78914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 78294 664000 78914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 -7654 114914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 222000 114914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 114294 664000 114914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 -7654 150914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 222000 150914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 150294 664000 150914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 -7654 186914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 222000 186914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 186294 664000 186914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 -7654 222914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 222000 222914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 222294 664000 222914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 258294 -7654 258914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 -7654 294914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 542000 294914 598000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 294294 642000 294914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 -7654 330914 58000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 222000 330914 278000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 330294 332000 330914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 -7654 366914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 366294 642000 366914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 -7654 402914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 402294 642000 402914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 438294 -7654 438914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 474294 -7654 474914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 -7654 510914 498000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 542000 510914 598000 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 510294 642000 510914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 546294 -7654 546914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 7366 592650 7986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 43366 592650 43986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 79366 592650 79986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 115366 592650 115986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 151366 592650 151986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 187366 592650 187986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 223366 592650 223986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 259366 592650 259986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 295366 592650 295986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 331366 592650 331986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 367366 592650 367986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 403366 592650 403986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 439366 592650 439986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 475366 592650 475986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 511366 592650 511986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 547366 592650 547986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 583366 592650 583986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 619366 592650 619986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 655366 592650 655986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 691366 592650 691986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 15294 -7654 15914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 -7654 51914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 51294 664000 51914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 -7654 87914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 222000 87914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87294 664000 87914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 -7654 123914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 222000 123914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 123294 664000 123914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 -7654 159914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 222000 159914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 159294 664000 159914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 -7654 195914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 222000 195914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 195294 664000 195914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 -7654 231914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 231294 664000 231914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 267294 -7654 267914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 -7654 303914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 222000 303914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 332000 303914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 542000 303914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 303294 642000 303914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 -7654 339914 58000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 222000 339914 278000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 339294 332000 339914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 -7654 375914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 552000 375914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 375294 642000 375914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 411294 -7654 411914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 447294 -7654 447914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 -7654 483914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 542000 483914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 483294 642000 483914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 -7654 519914 498000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 542000 519914 598000 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 519294 642000 519914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 555294 -7654 555914 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
