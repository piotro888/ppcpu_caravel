* NGSPICE file created from core.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt core dbg_in[0] dbg_in[1] dbg_in[2] dbg_in[3] dbg_out[0] dbg_out[10] dbg_out[11]
+ dbg_out[12] dbg_out[13] dbg_out[14] dbg_out[15] dbg_out[16] dbg_out[17] dbg_out[18]
+ dbg_out[19] dbg_out[1] dbg_out[20] dbg_out[21] dbg_out[22] dbg_out[23] dbg_out[24]
+ dbg_out[25] dbg_out[26] dbg_out[27] dbg_out[28] dbg_out[29] dbg_out[2] dbg_out[30]
+ dbg_out[31] dbg_out[32] dbg_out[33] dbg_out[34] dbg_out[35] dbg_out[3] dbg_out[4]
+ dbg_out[5] dbg_out[6] dbg_out[7] dbg_out[8] dbg_out[9] dbg_pc[0] dbg_pc[10] dbg_pc[11]
+ dbg_pc[12] dbg_pc[13] dbg_pc[14] dbg_pc[15] dbg_pc[1] dbg_pc[2] dbg_pc[3] dbg_pc[4]
+ dbg_pc[5] dbg_pc[6] dbg_pc[7] dbg_pc[8] dbg_pc[9] dbg_r0[0] dbg_r0[10] dbg_r0[11]
+ dbg_r0[12] dbg_r0[13] dbg_r0[14] dbg_r0[15] dbg_r0[1] dbg_r0[2] dbg_r0[3] dbg_r0[4]
+ dbg_r0[5] dbg_r0[6] dbg_r0[7] dbg_r0[8] dbg_r0[9] i_clk i_irq i_mem_ack i_mem_data[0]
+ i_mem_data[10] i_mem_data[11] i_mem_data[12] i_mem_data[13] i_mem_data[14] i_mem_data[15]
+ i_mem_data[1] i_mem_data[2] i_mem_data[3] i_mem_data[4] i_mem_data[5] i_mem_data[6]
+ i_mem_data[7] i_mem_data[8] i_mem_data[9] i_mem_exception i_req_data[0] i_req_data[10]
+ i_req_data[11] i_req_data[12] i_req_data[13] i_req_data[14] i_req_data[15] i_req_data[16]
+ i_req_data[17] i_req_data[18] i_req_data[19] i_req_data[1] i_req_data[20] i_req_data[21]
+ i_req_data[22] i_req_data[23] i_req_data[24] i_req_data[25] i_req_data[26] i_req_data[27]
+ i_req_data[28] i_req_data[29] i_req_data[2] i_req_data[30] i_req_data[31] i_req_data[3]
+ i_req_data[4] i_req_data[5] i_req_data[6] i_req_data[7] i_req_data[8] i_req_data[9]
+ i_req_data_valid i_rst o_c_data_page o_c_instr_page o_icache_flush o_mem_addr[0]
+ o_mem_addr[10] o_mem_addr[11] o_mem_addr[12] o_mem_addr[13] o_mem_addr[14] o_mem_addr[15]
+ o_mem_addr[1] o_mem_addr[2] o_mem_addr[3] o_mem_addr[4] o_mem_addr[5] o_mem_addr[6]
+ o_mem_addr[7] o_mem_addr[8] o_mem_addr[9] o_mem_data[0] o_mem_data[10] o_mem_data[11]
+ o_mem_data[12] o_mem_data[13] o_mem_data[14] o_mem_data[15] o_mem_data[1] o_mem_data[2]
+ o_mem_data[3] o_mem_data[4] o_mem_data[5] o_mem_data[6] o_mem_data[7] o_mem_data[8]
+ o_mem_data[9] o_mem_req o_mem_sel[0] o_mem_sel[1] o_mem_we o_req_active o_req_addr[0]
+ o_req_addr[10] o_req_addr[11] o_req_addr[12] o_req_addr[13] o_req_addr[14] o_req_addr[15]
+ o_req_addr[1] o_req_addr[2] o_req_addr[3] o_req_addr[4] o_req_addr[5] o_req_addr[6]
+ o_req_addr[7] o_req_addr[8] o_req_addr[9] o_req_ppl_submit sr_bus_addr[0] sr_bus_addr[10]
+ sr_bus_addr[11] sr_bus_addr[12] sr_bus_addr[13] sr_bus_addr[14] sr_bus_addr[15]
+ sr_bus_addr[1] sr_bus_addr[2] sr_bus_addr[3] sr_bus_addr[4] sr_bus_addr[5] sr_bus_addr[6]
+ sr_bus_addr[7] sr_bus_addr[8] sr_bus_addr[9] sr_bus_data_o[0] sr_bus_data_o[10]
+ sr_bus_data_o[11] sr_bus_data_o[12] sr_bus_data_o[13] sr_bus_data_o[14] sr_bus_data_o[15]
+ sr_bus_data_o[1] sr_bus_data_o[2] sr_bus_data_o[3] sr_bus_data_o[4] sr_bus_data_o[5]
+ sr_bus_data_o[6] sr_bus_data_o[7] sr_bus_data_o[8] sr_bus_data_o[9] sr_bus_we vccd1
+ vssd1
XFILLER_227_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3140__A1 _5660_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3140__B2 _5580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4935__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3155_ _5645_/Q _3147_/X _3149_/X _5565_/Q vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3086_ _2850_/D _3027_/X _3018_/A vssd1 vssd1 vccd1 vccd1 _3086_/X sky130_fd_sc_hd__a21o_1
XFILLER_254_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3979__A0 _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4640__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5766__A _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4928__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4670__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3988_ _5774_/A _5739_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3988_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5727_ _5741_/CLK _5727_/D vssd1 vssd1 vccd1 vccd1 _5727_/Q sky130_fd_sc_hd__dfxtp_1
X_2939_ _3775_/A _2937_/Y _2938_/X vssd1 vssd1 vccd1 vccd1 _2939_/X sky130_fd_sc_hd__a21bo_1
XFILLER_210_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5658_ _5658_/CLK _5658_/D vssd1 vssd1 vccd1 vccd1 _5658_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4609_ _5524_/Q _4619_/B vssd1 vssd1 vccd1 vccd1 _5198_/A sky130_fd_sc_hd__nand2_2
XFILLER_163_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5589_ _5653_/CLK _5589_/D vssd1 vssd1 vccd1 vccd1 _5589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4251__S0 _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2706__A1 _5637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2706__B2 _5669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4459__A1 _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5503__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2890__B1 _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__A1 _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5653__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3198__A1 _5670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3198__B2 _5590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3908__B _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4934__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4698__A1 _5557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5111__A2 _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4755__A _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4663_/X _4949_/Y _4959_/X _4957_/X vssd1 vssd1 vccd1 vccd1 _5663_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3911_ _5508_/Q _3245_/Y _3910_/X vssd1 vssd1 vccd1 vccd1 _5508_/D sky130_fd_sc_hd__a21o_1
XFILLER_251_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4891_ _4679_/X _4874_/Y _4890_/X _4886_/X vssd1 vssd1 vccd1 vccd1 _5634_/D sky130_fd_sc_hd__o211a_1
XFILLER_177_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_199_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4490__A _4600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3842_ _5291_/S _3842_/B vssd1 vssd1 vccd1 vccd1 _5294_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3189__A1 _5604_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3189__B2 _5620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3773_ _5458_/Q _3293_/X _3775_/A _3772_/Y vssd1 vssd1 vccd1 vccd1 _5458_/D sky130_fd_sc_hd__a22o_1
XFILLER_285_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _5741_/CLK _5512_/D vssd1 vssd1 vccd1 vccd1 _5512_/Q sky130_fd_sc_hd__dfxtp_2
X_2724_ _2775_/D _2727_/C _2775_/B _5603_/Q vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__and4b_1
XFILLER_157_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5443_ _5743_/CLK _5443_/D vssd1 vssd1 vccd1 vccd1 _5760_/A sky130_fd_sc_hd__dfxtp_4
X_2655_ _2655_/A vssd1 vssd1 vccd1 vccd1 _2655_/X sky130_fd_sc_hd__buf_4
XFILLER_105_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5374_ _5441_/CLK _5374_/D vssd1 vssd1 vccd1 vccd1 _5374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4325_ _4118_/B _3710_/X _3747_/X _3740_/X _4302_/S _4274_/A vssd1 vssd1 vccd1 vccd1
+ _4326_/B sky130_fd_sc_hd__mux4_1
XANTENNA__5526__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4256_ _4281_/A _4280_/B _4080_/X vssd1 vssd1 vccd1 vccd1 _4259_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5102__A2 _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4310__B1 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3207_ _5559_/Q _3131_/A _3204_/X _3206_/X vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__o22a_1
XFILLER_274_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5260__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4187_ _4372_/B _4175_/Y _4181_/X _4182_/X _4186_/Y vssd1 vssd1 vccd1 vccd1 _4187_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5676__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3138_ input3/X input1/X input2/X vssd1 vssd1 vccd1 vccd1 _3139_/A sky130_fd_sc_hd__nor3b_4
XFILLER_227_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _5401_/Q _5400_/Q _3069_/C vssd1 vssd1 vccd1 vccd1 _3075_/B sky130_fd_sc_hd__and3_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2913__A _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4916__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5326__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_30_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3655__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_364 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__C1 _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__A2 _4079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3919__A _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_392 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_169_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5549__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4469__B _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4386_/A _4386_/B _4368_/A _4368_/B _4386_/C vssd1 vssd1 vccd1 vccd1 _4110_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5699__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _4522_/B _5156_/B _5089_/X vssd1 vssd1 vccd1 vccd1 _5090_/Y sky130_fd_sc_hd__a21oi_1
X_4041_ _4025_/Y _4036_/Y _4038_/Y _4040_/X vssd1 vssd1 vccd1 vccd1 _4041_/X sky130_fd_sc_hd__a211o_2
XANTENNA__4485__A _4485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4843__A1 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _4981_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4943_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4932__B _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2733__A _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4874_ _5685_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4874_/Y sky130_fd_sc_hd__nand2_8
XFILLER_220_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4359__B1 _4355_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3825_ _3825_/A vssd1 vssd1 vccd1 vccd1 _5479_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5020__A1 _4537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3756_ _5461_/Q vssd1 vssd1 vccd1 vccd1 _4550_/S sky130_fd_sc_hd__inv_2
XANTENNA__3582__A1 _5477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2707_ _2757_/D vssd1 vssd1 vccd1 vccd1 _2775_/D sky130_fd_sc_hd__buf_4
XANTENNA__5308__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3687_ _4272_/S vssd1 vssd1 vccd1 vccd1 _4447_/S sky130_fd_sc_hd__buf_4
XFILLER_145_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5426_ _5441_/CLK _5426_/D vssd1 vssd1 vccd1 vccd1 _5426_/Q sky130_fd_sc_hd__dfxtp_1
X_2638_ _2682_/A _2747_/B _5627_/Q _2681_/A vssd1 vssd1 vccd1 vccd1 _2638_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__4379__B _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3334__B2 _5365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4531__B1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5357_ _5441_/CLK _5357_/D vssd1 vssd1 vccd1 vccd1 _5357_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4308_ _4271_/A _4307_/X _4116_/A vssd1 vssd1 vccd1 vccd1 _4308_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _5739_/Q _5774_/A _5291_/S vssd1 vssd1 vccd1 vccd1 _5289_/B sky130_fd_sc_hd__mux2_1
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4239_/X sky130_fd_sc_hd__xor2_1
XFILLER_261_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3637__A2 _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3503__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_261_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4598__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4842__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3739__A _4363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3458__B _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3573__A1 _5325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4289__B _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input55_A i_req_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2818__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__A1 _5606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3628__A2 _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3413__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output211_A _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5250__A1 _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5371__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3610_ _5643_/Q _3605_/X _3606_/X _3609_/X vssd1 vssd1 vccd1 vccd1 _3610_/X sky130_fd_sc_hd__a211o_1
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3013__B1 _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4590_ _5770_/A _4590_/B _4590_/C vssd1 vssd1 vccd1 vccd1 _4613_/C sky130_fd_sc_hd__and3_1
XFILLER_196_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3564__A1 _5628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3541_ _4229_/A _4301_/S vssd1 vssd1 vccd1 vccd1 _4124_/B sky130_fd_sc_hd__nor2_2
XANTENNA__3564__B2 _5596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3472_ _3472_/A vssd1 vssd1 vccd1 vccd1 _5416_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4199__B _4199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4513__A0 _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3316__A1 _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5211_ _5210_/X _5323_/A _5464_/Q vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5142_ _5155_/B _5142_/B vssd1 vssd1 vccd1 vccd1 _5142_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4927__B _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5069__A1 _5068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5073_ _5529_/Q _5051_/B _5055_/X _5489_/Q vssd1 vssd1 vccd1 vccd1 _5073_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4277__C1 _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4816__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4024_ _4024_/A _4024_/B vssd1 vssd1 vccd1 vccd1 _4084_/B sky130_fd_sc_hd__or2_2
XFILLER_244_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4943__A _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4044__A2 _4041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5714__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4926_ _4674_/X _4912_/Y _4925_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5649_/D sky130_fd_sc_hd__o211a_1
XFILLER_52_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4857_ _4970_/A _4859_/B vssd1 vssd1 vccd1 vccd1 _4857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5774__A _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3808_ _3808_/A vssd1 vssd1 vccd1 vccd1 _5471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4788_ _4976_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4788_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3739_ _4363_/B vssd1 vssd1 vccd1 vccd1 _4105_/B sky130_fd_sc_hd__clkinv_2
XFILLER_180_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5409_ _5743_/CLK _5409_/D vssd1 vssd1 vccd1 vccd1 _5409_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3858__A2 _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4837__B _4950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4268__C1 _4454_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4807__A1 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4283__A2 _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5394__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5232__A1 _2650_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4999__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output161_A _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3932__A _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4510__A3 _3761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4747__B _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_343 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5737__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4482__B _4482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5760_ _5760_/A vssd1 vssd1 vccd1 vccd1 _5760_/X sky130_fd_sc_hd__clkbuf_1
X_2972_ _2970_/Y _2850_/A _2968_/X _2971_/Y vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__o211a_1
XFILLER_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4711_ _5717_/Q vssd1 vssd1 vccd1 vccd1 _4711_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5724_/CLK _5691_/D vssd1 vssd1 vccd1 vccd1 _5691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4642_ _5680_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4642_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__3537__A1 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4573_ _4532_/X _4567_/Y _4568_/X _4572_/Y _4529_/X vssd1 vssd1 vccd1 vccd1 _4573_/X
+ sky130_fd_sc_hd__a311o_1
X_3524_ _3524_/A vssd1 vssd1 vccd1 vccd1 _5441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3455_ _5407_/Q _5408_/D _3475_/S vssd1 vssd1 vccd1 vccd1 _3456_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3842__A _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3386_ _3385_/X _5373_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3387_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5125_ _5125_/A vssd1 vssd1 vccd1 vccd1 _5193_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5056_ _5743_/Q _3840_/A _5055_/X _5488_/Q vssd1 vssd1 vccd1 vccd1 _5056_/X sky130_fd_sc_hd__a22o_1
XFILLER_284_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3988__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5769__A _5769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4007_ _4096_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__and2_1
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2905__B _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3225__B1 _3149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _5642_/Q _4897_/B _4907_/Y _4908_/X vssd1 vssd1 vccd1 vccd1 _5642_/D sky130_fd_sc_hd__o211a_1
XFILLER_112_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3752__A _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3700__A1 _5641_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input18_A i_mem_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_216_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5205__B2 _5505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3216__B1 _3145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4712__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4716__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2990__A2 _2850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output86_A _2863_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2742__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3240_ _5475_/Q _5474_/Q _5477_/Q _5476_/Q vssd1 vssd1 vccd1 vccd1 _3860_/B sky130_fd_sc_hd__nor4_1
XFILLER_3_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_239_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3171_ _5632_/Q _3143_/X _3145_/X _3170_/X vssd1 vssd1 vccd1 vccd1 _3171_/X sky130_fd_sc_hd__a211o_1
XANTENNA__2709__C _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5743_ _5743_/CLK _5743_/D vssd1 vssd1 vccd1 vccd1 _5743_/Q sky130_fd_sc_hd__dfxtp_1
X_2955_ _3308_/A _2943_/C _3283_/B _3307_/A _3293_/A vssd1 vssd1 vccd1 vccd1 _2955_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_194_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5674_ _5674_/CLK _5674_/D vssd1 vssd1 vccd1 vccd1 _5674_/Q sky130_fd_sc_hd__dfxtp_2
X_2886_ _5361_/Q _5360_/Q vssd1 vssd1 vccd1 vccd1 _2922_/A sky130_fd_sc_hd__nand2b_2
XFILLER_175_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4625_ _5773_/A _4511_/X _3919_/A _4624_/X vssd1 vssd1 vccd1 vccd1 _5545_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2981__A2 _2840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4556_ _5765_/A _4581_/B vssd1 vssd1 vccd1 vccd1 _4556_/X sky130_fd_sc_hd__or2_1
XFILLER_190_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3507_ _5433_/Q input39/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3508_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4668__A _4668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4487_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4487_/X sky130_fd_sc_hd__buf_4
X_3438_ _3438_/A vssd1 vssd1 vccd1 vccd1 _5398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4486__A2 _4485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3369_/A vssd1 vssd1 vccd1 vccd1 _5367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4891__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5109_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5108_/Y sky130_fd_sc_hd__nand2_1
XFILLER_245_302 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_257_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5039_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5039_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2916__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3511__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4850__B _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5432__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2972__A2 _2850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4174__A1 _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5582__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5123__A0 _5709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 _3227_/X vssd1 vssd1 vccd1 vccd1 dbg_out[15] sky130_fd_sc_hd__buf_2
Xoutput75 _5769_/A vssd1 vssd1 vccd1 vccd1 dbg_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__4477__A2 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 _2863_/Y vssd1 vssd1 vccd1 vccd1 dbg_out[35] sky130_fd_sc_hd__buf_2
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput97 _5772_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[12] sky130_fd_sc_hd__buf_2
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_381 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3685__B1 _3690_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2826__A _2826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output124_A _5556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3421__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_187 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_25_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4252__S _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2740_ _2727_/C _2789_/C _5650_/Q _2774_/C vssd1 vssd1 vccd1 vccd1 _2740_/X sky130_fd_sc_hd__and4b_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2671_ _2671_/A vssd1 vssd1 vccd1 vccd1 _5323_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__4165__A1 _4454_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4410_ _4410_/A _4410_/B vssd1 vssd1 vccd1 vccd1 _4483_/B sky130_fd_sc_hd__nand2_2
XFILLER_117_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5390_ _5404_/CLK _5390_/D vssd1 vssd1 vccd1 vccd1 _5390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4341_ _4454_/A _3749_/X _3555_/C _3650_/B _4116_/A vssd1 vssd1 vccd1 vccd1 _4341_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2715__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_220 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4272_ _4281_/A _4083_/B _4272_/S vssd1 vssd1 vccd1 vccd1 _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3223_ _5675_/Q _3137_/A _3139_/A _5595_/Q vssd1 vssd1 vccd1 vccd1 _3223_/X sky130_fd_sc_hd__a22o_1
XFILLER_100_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4873__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3140__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ _5597_/Q _3133_/X _3135_/X _5613_/Q _3153_/X vssd1 vssd1 vccd1 vccd1 _3154_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_254_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4935__B _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3085_ _3085_/A _3088_/B _3085_/C vssd1 vssd1 vccd1 vccd1 _3085_/Y sky130_fd_sc_hd__nor3_1
XFILLER_227_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5455__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3987_ _5525_/Q _3923_/A _3985_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5525_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3567__A _5660_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2938_ _3317_/A _2938_/B vssd1 vssd1 vccd1 vccd1 _2938_/X sky130_fd_sc_hd__or2_1
X_5726_ _5741_/CLK _5726_/D vssd1 vssd1 vccd1 vccd1 _5726_/Q sky130_fd_sc_hd__dfxtp_1
X_2869_ _5242_/S vssd1 vssd1 vccd1 vccd1 _3337_/B sky130_fd_sc_hd__buf_4
X_5657_ _5658_/CLK _5657_/D vssd1 vssd1 vccd1 vccd1 _5657_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4608_ _5771_/A _4581_/B _4602_/Y _4607_/X _3919_/X vssd1 vssd1 vccd1 vccd1 _5543_/D
+ sky130_fd_sc_hd__o221a_1
X_5588_ _5653_/CLK _5588_/D vssd1 vssd1 vccd1 vccd1 _5588_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_163_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4251__S1 _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2706__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4539_ _4536_/Y _4538_/X _4634_/A vssd1 vssd1 vccd1 vccd1 _4539_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5105__B1 _5051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4459__A2 _4289_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3667__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_346 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_245_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3419__A0 _2850_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2890__A1 _2928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4616__C1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4861__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2642__A1 _5595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3477__A _3523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3198__A2 _3137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4147__A1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_268_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_174_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_268_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3658__B1 _3608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4855__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4755__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4247__S _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5478__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4771__A _5583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3910_ _5510_/Q _3843_/B _3245_/B _4987_/A vssd1 vssd1 vccd1 vccd1 _3910_/X sky130_fd_sc_hd__a31o_1
X_4890_ _5634_/Q _4894_/A vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__or2_1
XANTENNA__3830__A0 _5482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _5743_/Q _4635_/A _3840_/X _4619_/B vssd1 vssd1 vccd1 vccd1 _3842_/B sky130_fd_sc_hd__a31o_1
XANTENNA__4490__B _4490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3189__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3772_ _3795_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _3772_/Y sky130_fd_sc_hd__nor2_1
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2723_ _2775_/B _2727_/C _2775_/D _5635_/Q vssd1 vssd1 vccd1 vccd1 _2723_/X sky130_fd_sc_hd__and4b_1
X_5511_ _5741_/CLK _5511_/D vssd1 vssd1 vccd1 vccd1 _5511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5442_ _5743_/CLK _5442_/D vssd1 vssd1 vccd1 vccd1 _5442_/Q sky130_fd_sc_hd__dfxtp_1
X_2654_ _5345_/Q _5346_/Q _5344_/Q vssd1 vssd1 vccd1 vccd1 _2655_/A sky130_fd_sc_hd__and3b_1
XFILLER_145_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5373_ _5757_/CLK _5373_/D vssd1 vssd1 vccd1 vccd1 _5373_/Q sky130_fd_sc_hd__dfxtp_1
X_4324_ _5453_/Q _4324_/B vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4011__A _4306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4255_ _4355_/A _4271_/A _4255_/C vssd1 vssd1 vccd1 vccd1 _4255_/X sky130_fd_sc_hd__and3_1
XANTENNA__3850__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4310__A1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3206_ _5639_/Q _3143_/A _3145_/A _3205_/X vssd1 vssd1 vccd1 vccd1 _3206_/X sky130_fd_sc_hd__a211o_1
X_4186_ _2954_/X _4046_/Y _4185_/X vssd1 vssd1 vccd1 vccd1 _4186_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_267_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_227_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3137_ _3137_/A vssd1 vssd1 vccd1 vccd1 _3137_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_227_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4384__C _4384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3068_ _5770_/A _3063_/B _3066_/Y _3067_/X _3016_/A vssd1 vssd1 vccd1 vccd1 _3068_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5709_ _5716_/CLK _5709_/D vssd1 vssd1 vccd1 vccd1 _5709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4856__A _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4301__A1 _3717_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2918__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output191_A _5474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3935__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4540__A1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4766__A _5581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4040_ _4192_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4040_/X sky130_fd_sc_hd__or2b_1
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4843__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2717__C _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _5656_/Q _4935_/B _4941_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5656_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3803__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4873_ _5627_/Q _4859_/B _4872_/Y _4862_/X vssd1 vssd1 vccd1 vccd1 _5627_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4359__A1 _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3824_ _5479_/Q _5383_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3825_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3755_ _4500_/A vssd1 vssd1 vccd1 vccd1 _3755_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_192_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2706_ _5637_/Q _2655_/X _2657_/X _5669_/Q vssd1 vssd1 vccd1 vccd1 _2706_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3582__A2 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3686_ _4278_/B _3686_/B vssd1 vssd1 vccd1 vccd1 _3686_/Y sky130_fd_sc_hd__nor2_1
Xoutput210 _5311_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[7] sky130_fd_sc_hd__buf_2
X_5425_ _5757_/CLK _5425_/D vssd1 vssd1 vccd1 vccd1 _5425_/Q sky130_fd_sc_hd__dfxtp_1
X_2637_ _5345_/Q vssd1 vssd1 vccd1 vccd1 _2747_/B sky130_fd_sc_hd__buf_2
XFILLER_279_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3056__S _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__C _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3334__A2 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4531__A1 _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5356_ _5743_/CLK _5356_/D vssd1 vssd1 vccd1 vccd1 _5356_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5643__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4307_ _4307_/A _4307_/B vssd1 vssd1 vccd1 vccd1 _4307_/X sky130_fd_sc_hd__or2_1
XFILLER_181_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5287_ _5287_/A vssd1 vssd1 vccd1 vccd1 _5738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3580__A _5476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5087__A2 _5086_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4238_ _4016_/X _4239_/A _4237_/Y vssd1 vssd1 vccd1 vccd1 _4238_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2908__B _5363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _4167_/Y _4168_/Y _4112_/C vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4598__A1 _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2924__A _5361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2697__A_N _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5300__A _5300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3458__C _3458_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3755__A _4500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4770__A1 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4289__C _4289_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input48_A i_req_data[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4586__A _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_238_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5078__A2 _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4825__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4589__A1 _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output204_A _2785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3261__A1 _5528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5516__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3013__A1 _2840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4210__B1 _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3564__A2 _3605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3540_ _3673_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _4301_/S sky130_fd_sc_hd__nand2_4
XFILLER_196_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5666__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3471_ _5416_/Q input52/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3472_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5210_ _4617_/Y _5209_/Y _5231_/S vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4513__A1 _5015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3316__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5141_ _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5142_/B sky130_fd_sc_hd__and2_1
XFILLER_269_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4496__A _4496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5072_ _5509_/Q _5094_/C _3996_/B _5082_/B _5493_/Q vssd1 vssd1 vccd1 vccd1 _5072_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_107 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2728__B _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4816__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4023_ _4348_/A _4087_/A _4071_/C _4069_/C vssd1 vssd1 vccd1 vccd1 _4023_/X sky130_fd_sc_hd__and4_1
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4943__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3559__B _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4925_ _5649_/Q _4931_/A vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__or2_1
X_4856_ _4856_/A vssd1 vssd1 vccd1 vccd1 _4859_/B sky130_fd_sc_hd__buf_4
XFILLER_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3807_ _5471_/Q _5375_/Q _3813_/S vssd1 vssd1 vccd1 vccd1 _3808_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4787_ _5590_/Q _4784_/B _4786_/Y _4769_/X vssd1 vssd1 vccd1 vccd1 _5590_/D sky130_fd_sc_hd__o211a_1
XFILLER_118_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4752__A1 _5575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3738_ _5558_/Q _3596_/X _3735_/X _3737_/X vssd1 vssd1 vccd1 vccd1 _4363_/B sky130_fd_sc_hd__o22a_4
XFILLER_109_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2763__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3669_ _5549_/Q _3596_/X _3666_/X _3668_/X vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__o22a_4
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_256_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5408_ _5722_/CLK _5408_/D vssd1 vssd1 vccd1 vccd1 _5408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2919__A _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5339_ _5686_/CLK _5339_/D vssd1 vssd1 vccd1 vccd1 _5339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4807__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5539__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5689__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_19_i_clk clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5659_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_109_131 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2829__A _2829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_219_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2971_ _5400_/Q _2966_/Y _2969_/X vssd1 vssd1 vccd1 vccd1 _2971_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4431__B1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _5560_/Q _4697_/A _4709_/Y _4670_/X vssd1 vssd1 vccd1 vccd1 _5560_/D sky130_fd_sc_hd__o211a_1
XFILLER_277_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4982__A1 _5673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5690_ _5724_/CLK _5690_/D vssd1 vssd1 vccd1 vccd1 _5690_/Q sky130_fd_sc_hd__dfxtp_1
X_4641_ _4950_/B vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__buf_12
XFILLER_147_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3537__A2 _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4734__A1 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4572_ _5154_/A _4571_/X _4634_/A vssd1 vssd1 vccd1 vccd1 _4572_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2745__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3523_ _5441_/Q input48/X _3523_/S vssd1 vssd1 vccd1 vccd1 _3524_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3454_ _3523_/S vssd1 vssd1 vccd1 vccd1 _3475_/S sky130_fd_sc_hd__buf_4
XFILLER_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3385_ input30/X _5425_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3385_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2739__A _5666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3170__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5124_ _5124_/A vssd1 vssd1 vccd1 vccd1 _5709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _5055_/A _5094_/B _5055_/C vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__and3_1
XANTENNA__4954__A _5661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4006_ _4006_/A _4006_/B vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__or2_4
XFILLER_84_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3225__A1 _5659_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3225__B2 _5579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4908_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4908_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__4973__A1 _5669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2984__B1 _2840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2735__A_N _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4839_ _5612_/Q _4872_/B vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__or2_1
XANTENNA__3509__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4489__B1 _5200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4848__B _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3161__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3700__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5361__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4864__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4661__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_231_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3216__A1 _5641_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4964__A1 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3419__S _3419_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3943__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output79_A _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5704__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3170_ _5648_/Q _3147_/X _3149_/X _5568_/Q vssd1 vssd1 vccd1 vccd1 _3170_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_21_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4652__A0 _5705_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3455__A1 _5408_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__C _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3207__A1 _5559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5742_ _5756_/CLK _5742_/D vssd1 vssd1 vccd1 vccd1 _5742_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4955__A1 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2954_ _5449_/Q vssd1 vssd1 vccd1 vccd1 _2954_/X sky130_fd_sc_hd__buf_4
XFILLER_187_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5673_ _5675_/CLK _5673_/D vssd1 vssd1 vccd1 vccd1 _5673_/Q sky130_fd_sc_hd__dfxtp_1
X_2885_ _4132_/A vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__buf_4
X_4624_ _4585_/A _4620_/X _4629_/B _4623_/X _4529_/X vssd1 vssd1 vccd1 vccd1 _4624_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4949__A _5687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4555_ _4551_/X _4554_/Y _4634_/A vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__mux2_1
X_3506_ _3506_/A vssd1 vssd1 vccd1 vccd1 _5432_/D sky130_fd_sc_hd__clkbuf_1
X_4486_ _3943_/A _4485_/A _4458_/A vssd1 vssd1 vccd1 vccd1 _4486_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5384__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3437_ _5398_/Q _3058_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3438_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3001_/C _5367_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3369_/A sky130_fd_sc_hd__mux2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3694__A1 _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3694__B2 _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5219_/S _5106_/X _4542_/Y vssd1 vssd1 vccd1 vccd1 _5109_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__4684__A _4684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3299_ _5365_/Q _5366_/Q _3297_/X _3795_/A _5337_/Q vssd1 vssd1 vccd1 vccd1 _5337_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_245_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5038_ _5038_/A vssd1 vssd1 vccd1 vccd1 _5699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2916__B _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4643__A0 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5199__A1 _5198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2932__A _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4946__A1 _5658_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_170 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2651__B _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4159__C1 _4372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4859__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2804__S0 _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5727__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5123__A1 _5122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput65 _5760_/A vssd1 vssd1 vccd1 vccd1 dbg_out[16] sky130_fd_sc_hd__buf_2
Xoutput76 _5770_/A vssd1 vssd1 vccd1 vccd1 dbg_out[26] sky130_fd_sc_hd__buf_2
Xoutput87 _3167_/X vssd1 vssd1 vccd1 vccd1 dbg_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput98 _5773_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[13] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A i_req_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output117_A _5549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3003__A _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2670_ _2665_/X _2666_/X _2669_/X _2791_/B _5561_/Q vssd1 vssd1 vccd1 vccd1 _2671_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_157_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4769__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4340_ _4454_/A _4182_/B _4271_/A vssd1 vssd1 vccd1 vccd1 _4340_/X sky130_fd_sc_hd__o21a_1
XFILLER_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4271_ _4271_/A _4271_/B vssd1 vssd1 vccd1 vccd1 _4271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3125__A0 _5710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_168 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3222_ _5562_/Q _3131_/A _3219_/X _3221_/X vssd1 vssd1 vccd1 vccd1 _3222_/X sky130_fd_sc_hd__o22a_2
XFILLER_86_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_239_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3153_ _5661_/Q _3137_/X _3139_/X _5581_/Q vssd1 vssd1 vccd1 vccd1 _3153_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _3084_/A _3084_/B vssd1 vssd1 vccd1 vccd1 _3085_/C sky130_fd_sc_hd__and2_1
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4625__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3848__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4928__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3986_ _5331_/A vssd1 vssd1 vccd1 vccd1 _3986_/X sky130_fd_sc_hd__buf_6
XFILLER_148_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5725_ _5740_/CLK _5725_/D vssd1 vssd1 vccd1 vccd1 _5725_/Q sky130_fd_sc_hd__dfxtp_1
X_2937_ _2949_/B _3304_/A _3799_/B vssd1 vssd1 vccd1 vccd1 _2937_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5656_ _5658_/CLK _5656_/D vssd1 vssd1 vccd1 vccd1 _5656_/Q sky130_fd_sc_hd__dfxtp_2
X_2868_ _3791_/A vssd1 vssd1 vccd1 vccd1 _5242_/S sky130_fd_sc_hd__clkinv_4
X_4607_ _4532_/X _4605_/Y _4606_/X _4529_/A vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4679__A _4679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5587_ _5667_/CLK _5587_/D vssd1 vssd1 vccd1 vccd1 _5587_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_190_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2799_ _3854_/A _5723_/Q _5722_/Q _3856_/C vssd1 vssd1 vccd1 vccd1 _2800_/A sky130_fd_sc_hd__or4_1
XFILLER_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4538_ _4600_/A _3943_/A _4537_/Y _5294_/A vssd1 vssd1 vccd1 vccd1 _4538_/X sky130_fd_sc_hd__a211o_1
XFILLER_116_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5105__B2 _5532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4469_ _4484_/A _4469_/B _4469_/C _4469_/D vssd1 vssd1 vccd1 vccd1 _4469_/Y sky130_fd_sc_hd__nand4_1
XFILLER_264_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3667__A1 _5565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3667__B2 _5581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4618__S _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2890__A2 _3799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4861__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2642__A2 _2635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3052__C1 _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3658__A1 _5567_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3658__B2 _5583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4607__B1 _4529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4771__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _3840_/A vssd1 vssd1 vccd1 vccd1 _3840_/X sky130_fd_sc_hd__buf_2
XFILLER_149_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3771_ _4987_/B _3771_/B vssd1 vssd1 vccd1 vccd1 _5457_/D sky130_fd_sc_hd__nor2_1
XANTENNA__3043__C1 _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3594__B1 _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5510_ _5741_/CLK _5510_/D vssd1 vssd1 vccd1 vccd1 _5510_/Q sky130_fd_sc_hd__dfxtp_1
X_2722_ _2722_/A vssd1 vssd1 vccd1 vccd1 _5313_/A sky130_fd_sc_hd__buf_4
XFILLER_285_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5441_ _5441_/CLK _5441_/D vssd1 vssd1 vccd1 vccd1 _5441_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4499__A _4543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2653_ _5594_/Q _2635_/Y _2652_/X _5626_/Q vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__a22o_2
XFILLER_160_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5372_ _5721_/CLK _5372_/D vssd1 vssd1 vccd1 vccd1 _5372_/Q sky130_fd_sc_hd__dfxtp_1
X_4323_ _4323_/A _4323_/B vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4011__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4254_ _4276_/A _4251_/X _4253_/X vssd1 vssd1 vccd1 vccd1 _4255_/C sky130_fd_sc_hd__a21oi_1
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3205_ _5655_/Q _3147_/A _3149_/A _5575_/Q vssd1 vssd1 vccd1 vccd1 _3205_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4310__A2 _4034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4185_ _2936_/X _4403_/A _4183_/Y _2904_/X _4184_/X vssd1 vssd1 vccd1 vccd1 _4185_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5422__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3136_ input3/X input2/X input1/X vssd1 vssd1 vccd1 vccd1 _3137_/A sky130_fd_sc_hd__and3_4
XFILLER_82_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3067_ _2966_/A _3027_/X _3018_/A vssd1 vssd1 vccd1 vccd1 _3067_/X sky130_fd_sc_hd__a21o_1
XFILLER_215_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_242_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5572__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3034__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3969_ _3990_/A _3969_/B vssd1 vssd1 vccd1 vccd1 _3969_/X sky130_fd_sc_hd__or2_1
XFILLER_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5708_ _5721_/CLK _5708_/D vssd1 vssd1 vccd1 vccd1 _5708_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2927__A3 _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5639_ _5658_/CLK _5639_/D vssd1 vssd1 vccd1 vccd1 _5639_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3517__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__A _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__A1 _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_233_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5179__S _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output184_A _5482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3427__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4112__A _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4469__D _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5445__CLK _5528_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_382 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4766__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output61_A _3212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2717__D _5588_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5595__CLK _5659_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4782__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _4978_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4941_/Y sky130_fd_sc_hd__nand2_1
XFILLER_224_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3803__A1 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3803__B2 _3802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5005__A0 _5685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4872_ _4985_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4872_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4359__A2 _4352_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3823_ _3823_/A vssd1 vssd1 vccd1 vccd1 _5478_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4006__B _4006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3754_ _4347_/A _3615_/X _3696_/X _3753_/X vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__a211oi_4
XFILLER_192_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_229_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2705_ _5573_/Q _2644_/X _2664_/X _5605_/Q vssd1 vssd1 vccd1 vccd1 _2705_/X sky130_fd_sc_hd__a22o_1
X_3685_ _3683_/X _4076_/B _3690_/C vssd1 vssd1 vccd1 vccd1 _3686_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2790__A1 _5612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4022__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5424_ _5441_/CLK _5424_/D vssd1 vssd1 vccd1 vccd1 _5424_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput200 _5321_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[12] sky130_fd_sc_hd__buf_2
X_2636_ _2761_/B _2682_/A _2681_/A _5643_/Q vssd1 vssd1 vccd1 vccd1 _2636_/X sky130_fd_sc_hd__and4b_1
Xoutput211 _5313_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4531__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4957__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5355_ _5404_/CLK _5355_/D vssd1 vssd1 vccd1 vccd1 _5355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3861__A _5471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4306_ _4306_/A _4326_/A vssd1 vssd1 vccd1 vccd1 _4306_/X sky130_fd_sc_hd__or2_1
X_5286_ _5292_/A _5286_/B vssd1 vssd1 vccd1 vccd1 _5287_/A sky130_fd_sc_hd__and2_1
X_4237_ _4016_/X _4239_/A _4350_/A vssd1 vssd1 vccd1 vccd1 _4237_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4168_ _4168_/A _4389_/A vssd1 vssd1 vccd1 vccd1 _4168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_255_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3119_ _5707_/Q _5715_/Q _4651_/S vssd1 vssd1 vccd1 vccd1 _3120_/A sky130_fd_sc_hd__mux2_1
X_4099_ _4102_/A _4101_/A vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__or2_1
XFILLER_215_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4598__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2924__B _5360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3101__A _5706_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4770__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5468__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3771__A _4987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3730__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4286__A1 _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4589__A2 _4581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4746__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2850__A _2850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3013__A2 _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3470_ _3470_/A vssd1 vssd1 vccd1 vccd1 _5415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4777__A _5586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3681__A _5529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3721__B1 _3602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _5219_/S _5140_/B vssd1 vssd1 vccd1 vccd1 _5154_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4496__B _5132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _5761_/A _5071_/B vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__or2_1
XANTENNA__4277__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2728__C _5651_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4022_ _4071_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4069_/C sky130_fd_sc_hd__xnor2_2
XFILLER_284_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2878__C_N _5363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4017__A _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4924_ _4668_/X _4912_/Y _4923_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5648_/D sky130_fd_sc_hd__o211a_1
XFILLER_212_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855_ _4684_/X _4836_/Y _4854_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5619_/D sky130_fd_sc_hd__o211a_1
XFILLER_220_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3856__A _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_i_clk_A clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3806_ _3806_/A vssd1 vssd1 vccd1 vccd1 _5470_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2760__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4786_ _4974_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5610__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2748__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3737_ _5638_/Q _3605_/X _3606_/X _3736_/X vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4752__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2763__A1 _5583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2763__B2 _5663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3668_ _5629_/Q _3605_/X _3606_/X _3667_/X vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__a211o_1
XFILLER_279_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5407_ _5743_/CLK _5407_/D vssd1 vssd1 vccd1 vccd1 _5407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5282__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3591__A _4128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3599_ _3601_/C _3599_/B _3601_/B vssd1 vssd1 vccd1 vccd1 _3600_/A sky130_fd_sc_hd__and3_4
XANTENNA__3712__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5338_ _5686_/CLK _5338_/D vssd1 vssd1 vccd1 vccd1 _5338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5269_ _5269_/A vssd1 vssd1 vccd1 vccd1 _5732_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4268__A1 _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2638__C _5627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4626__S _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5311__A _5311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4728__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_194 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_143 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3951__A0 _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_168 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4900__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2829__B _2829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_219_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5208__B1 _4619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2970_ _5399_/Q vssd1 vssd1 vccd1 vccd1 _2970_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4431__A1 _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5633__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4982__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3676__A _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ _5720_/Q input6/X _5679_/Q vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__mux2_4
XANTENNA__4719__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4571_ _4626_/S _4496_/A _4570_/Y _4619_/B vssd1 vssd1 vccd1 vccd1 _4571_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4734__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2745__A1 _5633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3942__A0 _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3522_ _3522_/A vssd1 vssd1 vccd1 vccd1 _5440_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2745__B2 _5665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3453_ _5457_/Q _3228_/A _3345_/A _5263_/A _3346_/B vssd1 vssd1 vccd1 vccd1 _3523_/S
+ sky130_fd_sc_hd__o2111a_2
XFILLER_115_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2739__B _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3384_ _3384_/A vssd1 vssd1 vccd1 vccd1 _5372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3170__A1 _5648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5123_ _5709_/Q _5122_/X _5135_/S vssd1 vssd1 vccd1 vccd1 _5124_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3170__B2 _5568_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5512_/Q _3931_/A _5053_/X vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__a21o_1
XFILLER_242_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4954__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4005_ _4108_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__and2_1
XFILLER_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3350__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4958__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4970__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3225__A2 _3147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4907_ _4983_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4907_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4973__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4838_ _4856_/A vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__buf_4
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4769_ _5331_/A vssd1 vssd1 vccd1 vccd1 _4769_/X sky130_fd_sc_hd__buf_4
XFILLER_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3161__A1 _5630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5506__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_275_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4864__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_263_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4661__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5656__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2672__B1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3216__A2 _3143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4964__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_96 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3924__B1 _3851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3435__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3152__A1 _5548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__D _5571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4790__A _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3207__A2 _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5741_ _5741_/CLK _5741_/D vssd1 vssd1 vccd1 vccd1 _5741_/Q sky130_fd_sc_hd__dfxtp_1
X_2953_ _2953_/A vssd1 vssd1 vccd1 vccd1 _5447_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4955__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5672_ _5675_/CLK _5672_/D vssd1 vssd1 vccd1 vccd1 _5672_/Q sky130_fd_sc_hd__dfxtp_2
X_2884_ _5454_/Q vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_187_193 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4623_ _5773_/A _4621_/B _4528_/A vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__o21a_1
XFILLER_135_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4554_ _4560_/B _4554_/B vssd1 vssd1 vccd1 vccd1 _4554_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4949__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3505_ _5432_/Q input38/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3506_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5529__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4485_ _4485_/A _4485_/B _4485_/C _4485_/D vssd1 vssd1 vccd1 vccd1 _4485_/X sky130_fd_sc_hd__and4_1
XANTENNA__4030__A _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3436_ _3436_/A vssd1 vssd1 vccd1 vccd1 _5397_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5117__A2_N _5125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4340__B1 _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3367_ _3367_/A vssd1 vssd1 vccd1 vccd1 _5366_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4965__A _5666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4891__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3694__A2 _3683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5679__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5106_ _4552_/B _5125_/A _5105_/X _5071_/B vssd1 vssd1 vccd1 vccd1 _5106_/X sky130_fd_sc_hd__a22o_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3298_ _3295_/Y _5366_/Q _3297_/X _3795_/A _5336_/Q vssd1 vssd1 vccd1 vccd1 _5336_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_245_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_186 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5037_ _5699_/Q _4600_/B _5135_/S vssd1 vssd1 vccd1 vccd1 _5038_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_i_clk clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5675_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4643__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_213_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4946__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4859__B _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2804__S1 _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 _5761_/A vssd1 vssd1 vccd1 vccd1 dbg_out[17] sky130_fd_sc_hd__buf_2
Xoutput77 _5771_/A vssd1 vssd1 vccd1 vccd1 dbg_out[27] sky130_fd_sc_hd__buf_2
Xoutput88 _3172_/X vssd1 vssd1 vccd1 vccd1 dbg_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__4875__A _5685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput99 _5774_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[14] sky130_fd_sc_hd__buf_2
XFILLER_248_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4882__A1 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A i_mem_exception vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2948__A1 _3799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3673__B _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4270_ _4347_/A _4250_/Y _4255_/X _4269_/Y vssd1 vssd1 vccd1 vccd1 _4522_/B sky130_fd_sc_hd__a211o_4
XFILLER_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3221_ _5642_/Q _3143_/A _3145_/A _3220_/X vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__a211o_1
XFILLER_79_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4873__A1 _5627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3152_ _5548_/Q _3131_/X _3141_/X _3151_/X vssd1 vssd1 vccd1 vccd1 _3152_/X sky130_fd_sc_hd__o22a_2
XFILLER_239_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__A_N _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _3084_/A _3084_/B vssd1 vssd1 vccd1 vccd1 _3088_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4625__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2736__C _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2875__A_N _5360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4928__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2752__B _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3985_ _3990_/A _3985_/B vssd1 vssd1 vccd1 vccd1 _3985_/X sky130_fd_sc_hd__or2_1
XANTENNA__5050__A1 _5760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2939__A1 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5724_ _5724_/CLK _5724_/D vssd1 vssd1 vccd1 vccd1 _5724_/Q sky130_fd_sc_hd__dfxtp_1
X_2936_ _5445_/Q vssd1 vssd1 vccd1 vccd1 _2936_/X sky130_fd_sc_hd__buf_4
XFILLER_210_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5655_ _5658_/CLK _5655_/D vssd1 vssd1 vccd1 vccd1 _5655_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5351__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2867_ _2867_/A vssd1 vssd1 vccd1 vccd1 _3791_/A sky130_fd_sc_hd__buf_2
XANTENNA__3864__A _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4606_ _5771_/A _4613_/C vssd1 vssd1 vccd1 vccd1 _4606_/X sky130_fd_sc_hd__or2_1
XFILLER_175_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5586_ _5680_/CLK _5586_/D vssd1 vssd1 vccd1 vccd1 _5586_/Q sky130_fd_sc_hd__dfxtp_4
X_2798_ _5487_/Q input5/X vssd1 vssd1 vccd1 vccd1 _3856_/C sky130_fd_sc_hd__and2_1
XANTENNA__3364__A1 _5365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4537_ _4635_/A _4537_/B vssd1 vssd1 vccd1 vccd1 _4537_/Y sky130_fd_sc_hd__nor2_1
XFILLER_190_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4468_ _4468_/A _4468_/B vssd1 vssd1 vccd1 vccd1 _4468_/X sky130_fd_sc_hd__or2_1
XANTENNA__4313__B1 _4305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3419_ _2850_/C _5389_/Q _3419_/S vssd1 vssd1 vccd1 vccd1 _3420_/A sky130_fd_sc_hd__mux2_1
X_4399_ _4399_/A _4399_/B _4399_/C vssd1 vssd1 vccd1 vccd1 _4399_/X sky130_fd_sc_hd__or3_1
XANTENNA__3667__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4616__A1 _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_245_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4395__A3 _4141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3774__A _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_268_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4855__A1 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3658__A2 _3607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4607__A1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3014__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3291__B1 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5374__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3770_ _3770_/A vssd1 vssd1 vccd1 vccd1 _5456_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2999__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2721_ _2715_/X _2716_/X _2719_/X _2720_/X vssd1 vssd1 vccd1 vccd1 _2722_/A sky130_fd_sc_hd__o31a_1
XFILLER_285_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3684__A _5453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5440_ _5722_/CLK _5440_/D vssd1 vssd1 vccd1 vccd1 _5440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2652_ _2652_/A vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__buf_8
XANTENNA__4499__B _4499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5371_ _5721_/CLK _5371_/D vssd1 vssd1 vccd1 vccd1 _5371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4322_ _4322_/A _4322_/B _4321_/X vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__or3b_1
XFILLER_172_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5099__A1 _4536_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4253_ _4454_/B _4252_/X _3617_/A vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__o21a_1
X_3204_ _5607_/Q _3133_/A _3135_/A _5623_/Q _3203_/X vssd1 vssd1 vccd1 vccd1 _3204_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_234_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4184_ _2919_/X _4045_/A _4059_/B _4333_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4184_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_274_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2747__B _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3135_ _3135_/A vssd1 vssd1 vccd1 vccd1 _3135_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_67_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3066_ _3085_/A _3066_/B vssd1 vssd1 vccd1 vccd1 _3066_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5717__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_250_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3968_ _3967_/X _5315_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3969_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2919_ _5450_/Q vssd1 vssd1 vccd1 vccd1 _2919_/X sky130_fd_sc_hd__buf_4
X_5707_ _5707_/CLK _5707_/D vssd1 vssd1 vccd1 vccd1 _5707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5285__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3899_ _5504_/Q _5321_/A _3905_/S vssd1 vssd1 vccd1 vccd1 _3900_/B sky130_fd_sc_hd__mux2_1
X_5638_ _5654_/CLK _5638_/D vssd1 vssd1 vccd1 vccd1 _5638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5569_ _5747_/CLK _5569_/D vssd1 vssd1 vccd1 vccd1 _5569_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2938__A _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2848__A0 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3328__A1 _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3009__A _5355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3443__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_394 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4782__B _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5253__A1 _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3679__A _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3264__A0 _5531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4940_ _5655_/Q _4935_/B _4939_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5655_/D sky130_fd_sc_hd__o211a_1
XFILLER_220_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3803__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_220_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4871_ _5626_/Q _4859_/B _4870_/Y _4862_/X vssd1 vssd1 vccd1 vccd1 _5626_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3822_ _5478_/Q _5382_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3823_/A sky130_fd_sc_hd__mux2_1
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _3750_/X _4355_/A _4271_/A vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__and3b_1
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2704_ _2704_/A vssd1 vssd1 vccd1 vccd1 _5317_/A sky130_fd_sc_hd__buf_4
XANTENNA__4303__A _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3684_ _5453_/Q _5447_/Q vssd1 vssd1 vccd1 vccd1 _3690_/C sky130_fd_sc_hd__or2_2
XFILLER_145_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5423_ _5757_/CLK _5423_/D vssd1 vssd1 vccd1 vccd1 _5423_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2790__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2635_ _2681_/A _2682_/A _5345_/Q vssd1 vssd1 vccd1 vccd1 _2635_/Y sky130_fd_sc_hd__nor3b_4
Xoutput201 _5323_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[13] sky130_fd_sc_hd__buf_2
XANTENNA__4022__B _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput212 _5315_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_145_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5354_ _5441_/CLK _5354_/D vssd1 vssd1 vccd1 vccd1 _5354_/Q sky130_fd_sc_hd__dfxtp_1
X_4305_ _4454_/A _4305_/B vssd1 vssd1 vccd1 vccd1 _4305_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4449__S _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5285_ _5738_/Q _5773_/A _5285_/S vssd1 vssd1 vccd1 vccd1 _5286_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _3617_/A _4230_/Y _4235_/X _4271_/A vssd1 vssd1 vccd1 vccd1 _4236_/X sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_12_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4167_ _4379_/B _4379_/C vssd1 vssd1 vccd1 vccd1 _4167_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3118_ _3118_/A vssd1 vssd1 vccd1 vccd1 _3118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_255_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4098_ _4097_/A _4132_/B _4192_/C vssd1 vssd1 vccd1 vccd1 _4101_/A sky130_fd_sc_hd__o21a_1
XANTENNA__5244__A1 _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3255__A0 _5528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3049_ _5397_/Q _3053_/C vssd1 vssd1 vccd1 vccd1 _3050_/B sky130_fd_sc_hd__xnor2_1
XFILLER_215_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3101__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3730__A1 _5620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4883__A _5631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3797__A1 _3310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_387 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2850__B _2850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5412__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3681__B _5466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3721__A1 _5669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5562__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5070_ _5070_/A vssd1 vssd1 vccd1 vccd1 _5704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4277__A2 _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4021_ _4027_/A _4027_/B vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__nor2_4
XANTENNA__2728__D _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4793__A _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5226__A1 _5527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3788__A1 _3791_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4923_ _5648_/Q _4931_/A vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__or2_1
XANTENNA__4017__B _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4854_ _5619_/Q _4856_/A vssd1 vssd1 vccd1 vccd1 _4854_/X sky130_fd_sc_hd__or2_1
X_3805_ _5470_/Q _5374_/Q _3813_/S vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__mux2_1
X_4785_ _5589_/Q _4784_/B _4784_/Y _4769_/X vssd1 vssd1 vccd1 vccd1 _5589_/D sky130_fd_sc_hd__o211a_1
XFILLER_165_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3736_ _5574_/Q _3607_/X _3608_/X _5590_/Q vssd1 vssd1 vccd1 vccd1 _3736_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4033__A _4033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2763__A2 _2635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3960__A1 _5311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3667_ _5565_/Q _3607_/X _3608_/X _5581_/Q vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3872__A _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5406_ _5743_/CLK _5406_/D vssd1 vssd1 vccd1 vccd1 _5406_/Q sky130_fd_sc_hd__dfxtp_1
X_3598_ _3598_/A vssd1 vssd1 vccd1 vccd1 _3598_/X sky130_fd_sc_hd__buf_6
XANTENNA__3712__A1 _5674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3241__A_N _5472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5337_ _5707_/CLK _5337_/D vssd1 vssd1 vccd1 vccd1 _5337_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3712__B2 _5658_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _5292_/A _5268_/B vssd1 vssd1 vccd1 vccd1 _5269_/A sky130_fd_sc_hd__and2_1
XFILLER_275_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4219_ _4192_/B _4210_/X _4218_/X vssd1 vssd1 vccd1 vccd1 _5156_/A sky130_fd_sc_hd__o21bai_4
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5199_ _5198_/A _5198_/C _5198_/B vssd1 vssd1 vccd1 vccd1 _5225_/B sky130_fd_sc_hd__a21o_1
XANTENNA__3811__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5435__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2939__B1_N _2938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5039__A _5200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5585__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3782__A _5461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input53_A i_req_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5208__A1 _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2845__B _2845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4118__A _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3219__B1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3022__A _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4431__A2 _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2861__A _5300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2993__A2 _2835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4570_ _4626_/S _5311_/A vssd1 vssd1 vccd1 vccd1 _4570_/Y sky130_fd_sc_hd__nor2_1
X_3521_ _5440_/Q input47/X _3523_/S vssd1 vssd1 vccd1 vccd1 _3522_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2745__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4788__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3452_ _3452_/A vssd1 vssd1 vccd1 vccd1 _5405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3383_ _3382_/X _5372_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3384_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2739__C _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5122_ _5121_/X _5307_/A _5179_/S vssd1 vssd1 vccd1 vccd1 _5122_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3170__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5053_ _5471_/Q _5094_/B _5055_/C vssd1 vssd1 vccd1 vccd1 _5053_/X sky130_fd_sc_hd__and3_2
XFILLER_284_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4655__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ _5479_/Q _3532_/X _3584_/X vssd1 vssd1 vccd1 vccd1 _4108_/A sky130_fd_sc_hd__a21o_2
XFILLER_272_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_225_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4028__A _4033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5458__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4970__B _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3867__A _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2771__A _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4906_ _5641_/Q _4897_/B _4905_/Y _4886_/X vssd1 vssd1 vccd1 vccd1 _5641_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3630__B1 _3606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2984__A2 _2845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4837_ _5684_/Q _4950_/B vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__and2_4
XFILLER_193_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4186__A1 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4768_ _5582_/Q _4797_/B vssd1 vssd1 vccd1 vccd1 _4768_/X sky130_fd_sc_hd__or2_1
XFILLER_267_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3719_ _3717_/Y _4307_/A _4272_/S vssd1 vssd1 vccd1 vccd1 _4454_/C sky130_fd_sc_hd__mux2_1
X_4699_ _5714_/Q vssd1 vssd1 vccd1 vccd1 _4699_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5135__A0 _5710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3697__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3107__A _5709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3161__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2781__A_N _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4110__A1 _4386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2672__A1 _5576_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2672__B2 _5608_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3924__A1 _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3152__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3451__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5600__CLK _5680_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4790__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3687__A _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5750__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2952_ _4350_/A _2951_/X _3337_/B vssd1 vssd1 vccd1 vccd1 _2953_/A sky130_fd_sc_hd__mux2_1
X_5740_ _5740_/CLK _5740_/D vssd1 vssd1 vccd1 vccd1 _5740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4696__A1_N input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2883_ _5455_/Q _5486_/D _2882_/Y vssd1 vssd1 vccd1 vccd1 _5455_/D sky130_fd_sc_hd__o21a_1
XANTENNA__2820__D1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5671_ _5675_/CLK _5671_/D vssd1 vssd1 vccd1 vccd1 _5671_/Q sky130_fd_sc_hd__dfxtp_2
X_4622_ _4622_/A vssd1 vssd1 vccd1 vccd1 _4629_/B sky130_fd_sc_hd__inv_2
XANTENNA__2654__A_N _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4553_ _4552_/B _4552_/C _5765_/A vssd1 vssd1 vccd1 vccd1 _4554_/B sky130_fd_sc_hd__a21oi_1
XFILLER_190_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3504_ _3504_/A vssd1 vssd1 vccd1 vccd1 _5431_/D sky130_fd_sc_hd__clkbuf_1
X_4484_ _4484_/A _4484_/B _4484_/C vssd1 vssd1 vccd1 vccd1 _4485_/D sky130_fd_sc_hd__or3_1
XFILLER_143_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3435_ _5397_/Q _3052_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3436_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4030__B _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4340__A1 _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3366_ _3001_/A _5366_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3367_/A sky130_fd_sc_hd__mux2_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4891__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5745_/Q _3840_/A _5051_/B _5532_/Q _5104_/X vssd1 vssd1 vccd1 vccd1 _5105_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_1_i_clk clkbuf_1_0_1_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_97_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3297_ _5367_/Q _3297_/B vssd1 vssd1 vccd1 vccd1 _3297_/X sky130_fd_sc_hd__and2b_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5036_ _5036_/A vssd1 vssd1 vccd1 vccd1 _5698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_257_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4981__A _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5288__S _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3597__A _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3603__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5317__A _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4867__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput67 _5762_/A vssd1 vssd1 vccd1 vccd1 dbg_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__4331__A1 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 _5772_/A vssd1 vssd1 vccd1 vccd1 dbg_out[28] sky130_fd_sc_hd__buf_2
Xoutput89 _3177_/X vssd1 vssd1 vccd1 vccd1 dbg_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__4875__B _4950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4882__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input16_A i_mem_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3300__A _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2948__A2 _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_172_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4131__A _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3673__C _4076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output84_A _5357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4858__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3220_ _5658_/Q _3147_/A _3149_/A _5578_/Q vssd1 vssd1 vccd1 vccd1 _3220_/X sky130_fd_sc_hd__a22o_1
XFILLER_97_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4873__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3151_ _5628_/Q _3143_/X _3145_/X _3150_/X vssd1 vssd1 vccd1 vccd1 _3151_/X sky130_fd_sc_hd__a211o_1
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3082_ _5773_/A _3010_/X _3081_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3082_/X sky130_fd_sc_hd__o211a_1
XFILLER_94_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2736__D _5570_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4625__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_254_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_235_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4306__A _4306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2752__C _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3984_ _3983_/X _5323_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3985_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5050__A2 _5125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2939__A2 _2937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5723_ _5741_/CLK _5723_/D vssd1 vssd1 vccd1 vccd1 _5723_/Q sky130_fd_sc_hd__dfxtp_1
X_2935_ _2919_/X _3780_/A _2931_/X _2934_/X vssd1 vssd1 vccd1 vccd1 _5450_/D sky130_fd_sc_hd__o22a_1
XFILLER_175_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5654_ _5654_/CLK _5654_/D vssd1 vssd1 vccd1 vccd1 _5654_/Q sky130_fd_sc_hd__dfxtp_1
X_2866_ _3228_/A _3771_/B vssd1 vssd1 vccd1 vccd1 _2867_/A sky130_fd_sc_hd__or2_1
XFILLER_108_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3864__B _4988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _4605_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3356__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2797_ _3000_/S vssd1 vssd1 vccd1 vccd1 _3768_/S sky130_fd_sc_hd__buf_4
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5585_ _5667_/CLK _5585_/D vssd1 vssd1 vccd1 vccd1 _5585_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_163_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5646__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4536_ _5515_/Q _4599_/B vssd1 vssd1 vccd1 vccd1 _4536_/Y sky130_fd_sc_hd__nand2_2
XFILLER_190_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4976__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4467_ _4467_/A _4467_/B vssd1 vssd1 vccd1 vccd1 _4474_/B sky130_fd_sc_hd__xnor2_1
XFILLER_117_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4849__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4313__A1 _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4313__B2 _4309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3418_ _3418_/A vssd1 vssd1 vccd1 vccd1 _5388_/D sky130_fd_sc_hd__clkbuf_1
X_4398_ _4468_/A _4250_/Y _4397_/X vssd1 vssd1 vccd1 vccd1 _4399_/C sky130_fd_sc_hd__o21ba_1
XFILLER_277_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input8_A i_mem_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ _3419_/S vssd1 vssd1 vccd1 vccd1 _3368_/S sky130_fd_sc_hd__buf_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4616__A2 _4581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5019_ _5019_/A vssd1 vssd1 vccd1 vccd1 _5690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3824__A0 _5479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3052__A1 _5539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4886__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4855__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output122_A _5554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_251_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3291__A1 _5365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5519__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3579__C1 _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3043__A1 _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3594__A2 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2720_ _5556_/Q _2720_/B vssd1 vssd1 vccd1 vccd1 _2720_/X sky130_fd_sc_hd__or2_1
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5669__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2651_ _5346_/Q _5345_/Q _5344_/Q vssd1 vssd1 vccd1 vccd1 _2652_/A sky130_fd_sc_hd__nor3b_4
XFILLER_200_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_i_clk clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5674_/CLK sky130_fd_sc_hd__clkbuf_16
X_5370_ _5757_/CLK _5370_/D vssd1 vssd1 vccd1 vccd1 _5370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4321_ _4348_/A _4348_/C _4032_/X _4069_/C vssd1 vssd1 vccd1 vccd1 _4321_/X sky130_fd_sc_hd__a211o_1
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4252_ _3717_/Y _4307_/A _4447_/S vssd1 vssd1 vccd1 vccd1 _4252_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3203_ _5671_/Q _3137_/A _3139_/A _5591_/Q vssd1 vssd1 vccd1 vccd1 _3203_/X sky130_fd_sc_hd__a22o_1
XFILLER_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4183_ _4183_/A vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2747__C _5649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3134_ input2/X input1/X input3/X vssd1 vssd1 vccd1 vccd1 _3135_/A sky130_fd_sc_hd__nor3b_4
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3065_ _5400_/Q _3069_/C vssd1 vssd1 vccd1 vccd1 _3066_/B sky130_fd_sc_hd__xnor2_1
XFILLER_242_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4231__A0 _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3034__A1 _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3967_ _4590_/B _5734_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3967_/X sky130_fd_sc_hd__mux2_1
XFILLER_259_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5706_ _5743_/CLK _5706_/D vssd1 vssd1 vccd1 vccd1 _5706_/Q sky130_fd_sc_hd__dfxtp_2
X_2918_ _5448_/Q _5486_/D _2917_/X vssd1 vssd1 vccd1 vccd1 _5448_/D sky130_fd_sc_hd__o21a_1
X_3898_ _5263_/A vssd1 vssd1 vccd1 vccd1 _5261_/A sky130_fd_sc_hd__buf_2
X_5637_ _5654_/CLK _5637_/D vssd1 vssd1 vccd1 vccd1 _5637_/Q sky130_fd_sc_hd__dfxtp_4
X_2849_ input47/X _5440_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2850_/D sky130_fd_sc_hd__mux2_2
XFILLER_275_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5568_ _5667_/CLK _5568_/D vssd1 vssd1 vccd1 vccd1 _5568_/Q sky130_fd_sc_hd__dfxtp_2
X_4519_ _4634_/A _4517_/Y _4518_/X _4529_/A vssd1 vssd1 vccd1 vccd1 _4519_/X sky130_fd_sc_hd__a31o_1
X_5499_ _5740_/CLK _5499_/D vssd1 vssd1 vccd1 vccd1 _5499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2938__B _2938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2954__A _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4645__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2784__B1 _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3328__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4525__A1 _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3009__B _5678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5341__CLK _5680_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4555__S _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3679__B _4076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3264__A1 _5532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4870_ _4983_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4870_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5491__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3821_ _3821_/A vssd1 vssd1 vccd1 vccd1 _5477_/D sky130_fd_sc_hd__clkbuf_1
X_3752_ _4326_/A vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__buf_2
X_2703_ _5558_/Q _2720_/B _2699_/X _2702_/X vssd1 vssd1 vccd1 vccd1 _2704_/A sky130_fd_sc_hd__o22a_1
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _3683_/A _3683_/B vssd1 vssd1 vccd1 vccd1 _3683_/X sky130_fd_sc_hd__and2_1
X_5422_ _5757_/CLK _5422_/D vssd1 vssd1 vccd1 vccd1 _5422_/Q sky130_fd_sc_hd__dfxtp_1
X_2634_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2791_/B sky130_fd_sc_hd__buf_6
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput202 _5325_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput213 _3250_/A vssd1 vssd1 vccd1 vccd1 sr_bus_we sky130_fd_sc_hd__buf_2
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5353_ _5692_/CLK _5353_/D vssd1 vssd1 vccd1 vccd1 _5353_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3634__S _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4304_ _4301_/X _4303_/Y _4304_/S vssd1 vssd1 vccd1 vccd1 _4305_/B sky130_fd_sc_hd__mux2_2
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5284_ _5284_/A vssd1 vssd1 vccd1 vccd1 _5737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4235_ _4454_/B _4231_/X _4303_/A _4276_/A _4234_/Y vssd1 vssd1 vccd1 vccd1 _4235_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_141_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4166_ _4171_/A _4114_/Y _4115_/X _4165_/X vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__o31a_1
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3117_ _5706_/Q _5714_/Q _4651_/S vssd1 vssd1 vccd1 vccd1 _3118_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4097_ _4097_/A _4132_/B _4192_/C vssd1 vssd1 vccd1 vccd1 _4102_/A sky130_fd_sc_hd__nor3_1
XFILLER_255_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3048_ _5766_/A _3010_/X _3046_/Y _3047_/X _3016_/A vssd1 vssd1 vccd1 vccd1 _3048_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3255__A1 _5530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4204__A0 _4121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4999_ _5682_/Q _5336_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _5000_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3809__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5180__A1 _5179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_278_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5325__A _5325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3191__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3730__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2668__B _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5364__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_278_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4883__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5060__A _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2756__B_N _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3719__S _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4404__A _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4746__A1 _5572_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2850__C _2850_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5707__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3721__A2 _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4020_ _4034_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4071_/C sky130_fd_sc_hd__xor2_2
XFILLER_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4682__A0 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4793__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4922_ _4663_/X _4912_/Y _4921_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5647_/D sky130_fd_sc_hd__o211a_1
XFILLER_252_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2996__B1 _2850_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4853_ _4679_/X _4836_/Y _4852_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5618_/D sky130_fd_sc_hd__o211a_1
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3804_ _3775_/X _2934_/X _3293_/X _5469_/Q vssd1 vssd1 vccd1 vccd1 _5469_/D sky130_fd_sc_hd__a2bb2o_1
X_4784_ _4972_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3735_ _5622_/Q _3597_/X _3598_/X _5606_/Q _3734_/X vssd1 vssd1 vccd1 vccd1 _3735_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4033__B _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3666_ _5613_/Q _3597_/X _3598_/X _5597_/Q _3665_/X vssd1 vssd1 vccd1 vccd1 _3666_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_256_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5405_ _5722_/CLK _5405_/D vssd1 vssd1 vccd1 vccd1 _5405_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5162__A1 _5521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5387__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2769__A _5662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3597_ _3597_/A vssd1 vssd1 vccd1 vccd1 _3597_/X sky130_fd_sc_hd__buf_6
XANTENNA__3364__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3173__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5336_ _5686_/CLK _5336_/D vssd1 vssd1 vccd1 vccd1 _5336_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3712__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_303 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5267_ _5732_/Q _5539_/Q _5285_/S vssd1 vssd1 vccd1 vccd1 _5268_/B sky130_fd_sc_hd__mux2_1
X_4218_ _4132_/B _4333_/A _4212_/X _4201_/Y _4217_/X vssd1 vssd1 vccd1 vccd1 _4218_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4673__A0 _5709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5198_ _5198_/A _5198_/B _5198_/C vssd1 vssd1 vccd1 vccd1 _5198_/Y sky130_fd_sc_hd__nand3_1
XFILLER_205_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4149_ _4132_/A _4063_/A _3613_/X _4469_/C _4469_/B vssd1 vssd1 vccd1 vccd1 _4149_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_28_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4208__B _4208_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2987__B1 _2852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4728__A1 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4224__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3164__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4900__A1 _5638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2911__A0 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input46_A i_req_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4894__A _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2845__C _2845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3219__A1 _5610_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3219__B2 _5626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3022__B _3063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output202_A _5325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2861__B _3343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4134__A _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4719__A1 _5562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _3520_/A vssd1 vssd1 vccd1 vccd1 _5439_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4788__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3451_ _5405_/Q _3091_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3452_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3155__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3382_ input29/X _5424_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3382_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2902__A0 _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2739__D _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5121_ _5119_/Y _5120_/X _4499_/B _5156_/B vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_111_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _5508_/Q _5094_/C _3996_/B _5082_/B _5492_/Q vssd1 vssd1 vccd1 vccd1 _5052_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_111_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_284_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4003_ _4043_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__nand2_1
XFILLER_242_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5131__C _5131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4028__B _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4958__A1 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4905_ _4981_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4905_/Y sky130_fd_sc_hd__nand2_1
XFILLER_240_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2771__B _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3630__A1 _5632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3091__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4836_ _5684_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4836_/Y sky130_fd_sc_hd__nand2_8
XFILLER_138_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_267_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4979__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4767_ _4653_/X _4761_/Y _4766_/X _4745_/X vssd1 vssd1 vccd1 vccd1 _5581_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3394__A0 _2845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3718_ _3732_/A _4484_/A vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__nand2_2
XFILLER_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4698_ _5557_/Q _4697_/A _4697_/Y _4670_/X vssd1 vssd1 vccd1 vccd1 _5557_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5135__A1 _5134_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3649_ _3635_/Y _3647_/Y _4454_/B vssd1 vssd1 vccd1 vccd1 _3650_/B sky130_fd_sc_hd__mux2_1
XFILLER_283_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3697__A1 _5673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3697__B2 _5657_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3107__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5319_ _5319_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5319_/X sky130_fd_sc_hd__or2_1
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3822__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3449__A1 _3087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4110__A2 _4386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2672__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3082__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5552__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_i_clk clkbuf_2_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_i_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_129_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3909__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__S0 _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4582__C1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5126__A1 _5518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4637__B1 _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_254_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_266_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _3791_/C _2951_/B _3318_/C _3308_/D vssd1 vssd1 vccd1 vccd1 _2951_/X sky130_fd_sc_hd__or4_1
XANTENNA__3073__C1 _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ _5675_/CLK _5670_/D vssd1 vssd1 vccd1 vccd1 _5670_/Q sky130_fd_sc_hd__dfxtp_2
X_2882_ _2949_/A _2877_/Y _3799_/A _2938_/B _3337_/B vssd1 vssd1 vccd1 vccd1 _2882_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4621_ _5773_/A _4621_/B vssd1 vssd1 vccd1 vccd1 _4622_/A sky130_fd_sc_hd__and2_1
XANTENNA__4799__A _5683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4573__C1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552_ _5765_/A _4552_/B _4552_/C vssd1 vssd1 vccd1 vccd1 _4560_/B sky130_fd_sc_hd__and3_1
XFILLER_128_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3503_ _5431_/Q input37/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3504_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5117__B2 _5460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4483_ _4483_/A _4483_/B vssd1 vssd1 vccd1 vccd1 _4485_/C sky130_fd_sc_hd__xnor2_1
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3434_ _3434_/A vssd1 vssd1 vccd1 vccd1 _5396_/D sky130_fd_sc_hd__clkbuf_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _3365_/A vssd1 vssd1 vccd1 vccd1 _5365_/D sky130_fd_sc_hd__clkbuf_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5425__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5104_ _5516_/Q _3931_/A _5082_/B _5496_/Q _5053_/X vssd1 vssd1 vccd1 vccd1 _5104_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_253_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3295_/Y _3292_/X _3293_/X _5335_/Q vssd1 vssd1 vccd1 vccd1 _5335_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_253_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5035_ _5698_/Q _4490_/B _5135_/S vssd1 vssd1 vccd1 vccd1 _5036_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4039__A _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4981__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5575__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3064__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3603__A1 _5675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3603__B2 _5659_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4819_ _4819_/A vssd1 vssd1 vccd1 vccd1 _4822_/B sky130_fd_sc_hd__buf_6
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3119__A0 _5707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput68 _5763_/A vssd1 vssd1 vccd1 vccd1 dbg_out[19] sky130_fd_sc_hd__buf_2
Xoutput79 _5773_/A vssd1 vssd1 vccd1 vccd1 dbg_out[29] sky130_fd_sc_hd__buf_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4095__A1 _4034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2692__A _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5448__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output77_A _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2867__A _2867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _5644_/Q _3147_/X _3149_/X _5564_/Q vssd1 vssd1 vccd1 vccd1 _3150_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3081_ _2845_/A _3089_/A _3084_/B _3080_/X _3018_/A vssd1 vssd1 vccd1 vccd1 _3081_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4086__A1 _4240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_242_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_250_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4306__B _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3983_ _5773_/A _5738_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3983_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2752__D _5600_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5722_ _5722_/CLK _5722_/D vssd1 vssd1 vccd1 vccd1 _5722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2934_ _3293_/A _2934_/B vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__or2_1
XANTENNA__4794__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5653_ _5653_/CLK _5653_/D vssd1 vssd1 vccd1 vccd1 _5653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2865_ _5678_/Q _5300_/A _2865_/C vssd1 vssd1 vccd1 vccd1 _3771_/B sky130_fd_sc_hd__or3_1
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4604_ _4604_/A _4604_/B vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4322__A _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5584_ _5667_/CLK _5584_/D vssd1 vssd1 vccd1 vccd1 _5584_/Q sky130_fd_sc_hd__dfxtp_1
X_2796_ _2849_/S vssd1 vssd1 vccd1 vccd1 _3000_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_7_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4535_ _5081_/A _4533_/C _4527_/C _5763_/A vssd1 vssd1 vccd1 vccd1 _4535_/X sky130_fd_sc_hd__a31o_1
XFILLER_264_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4466_ _4466_/A _4466_/B vssd1 vssd1 vccd1 vccd1 _4467_/B sky130_fd_sc_hd__and2_1
XFILLER_89_116 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4976__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3417_ _2850_/D _5388_/Q _3419_/S vssd1 vssd1 vccd1 vccd1 _3418_/A sky130_fd_sc_hd__mux2_1
X_4397_ _4372_/A _4396_/A _4395_/X _4396_/Y _4372_/B vssd1 vssd1 vccd1 vccd1 _4397_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3348_ _5357_/Q _3346_/Y _3435_/S vssd1 vssd1 vccd1 vccd1 _5357_/D sky130_fd_sc_hd__a21o_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3308_/C _3308_/D _3278_/Y vssd1 vssd1 vccd1 vccd1 _3287_/C sky130_fd_sc_hd__or3b_1
XFILLER_93_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _5690_/Q _4522_/B _5030_/S vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__mux2_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3285__C1 _2938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2943__C _2943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3588__A0 _5481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4785__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4232__A _4301_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5740__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5063__A _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4068__A1 _4467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_i_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_91_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output115_A _5562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4407__A _4408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3291__A2 _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3579__B1 _2726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4776__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3594__A3 _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_i_clk/A
+ sky130_fd_sc_hd__clkbuf_8
X_2650_ _4635_/B vssd1 vssd1 vccd1 vccd1 _2650_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_145_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4320_ _4347_/A _4320_/B vssd1 vssd1 vccd1 vccd1 _4320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4251_ _4118_/B _3710_/X _3747_/X _3740_/X _4231_/S _4304_/S vssd1 vssd1 vccd1 vccd1
+ _4251_/X sky130_fd_sc_hd__mux4_2
X_3202_ _5558_/Q _3131_/A _3199_/X _3201_/X vssd1 vssd1 vccd1 vccd1 _3202_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4182_ _4454_/A _4182_/B _4454_/D vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__or3_1
XFILLER_274_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2711__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2747__D _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3133_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3133_/X sky130_fd_sc_hd__buf_4
XFILLER_227_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3064_ _3343_/C _3062_/X _3063_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3064_/X sky130_fd_sc_hd__o211a_1
XFILLER_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_241 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4767__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4231__A1 _4024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ _5520_/Q _3923_/X _3965_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5520_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5613__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5705_ _5721_/CLK _5705_/D vssd1 vssd1 vccd1 vccd1 _5705_/Q sky130_fd_sc_hd__dfxtp_1
X_2917_ _3307_/A _3775_/A _3775_/C _3795_/A vssd1 vssd1 vccd1 vccd1 _2917_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3897_ _3895_/Y _3874_/B _3896_/Y vssd1 vssd1 vccd1 vccd1 _5503_/D sky130_fd_sc_hd__a21oi_1
XFILLER_12_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5148__A _5520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5636_ _5654_/CLK _5636_/D vssd1 vssd1 vccd1 vccd1 _5636_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2848_ input48/X _5441_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2850_/C sky130_fd_sc_hd__mux2_2
XANTENNA__4987__A _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5567_ _5738_/CLK _5567_/D vssd1 vssd1 vccd1 vccd1 _5567_/Q sky130_fd_sc_hd__dfxtp_2
X_2779_ _5629_/Q _2655_/X _2761_/X _5645_/Q vssd1 vssd1 vccd1 vccd1 _2779_/X sky130_fd_sc_hd__a22o_1
XFILLER_275_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3742__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4518_ _4533_/C _4527_/C vssd1 vssd1 vccd1 vccd1 _4518_/X sky130_fd_sc_hd__or2_1
X_5498_ _5741_/CLK _5498_/D vssd1 vssd1 vccd1 vccd1 _5498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4449_ _4448_/Y _4424_/B _4449_/S vssd1 vssd1 vccd1 vccd1 _4449_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2667__A_N _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2702__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3830__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4470__A1 _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3131__A _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4470__B2 _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_214_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4758__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2784__B2 _5549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4897__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4930__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3041__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3820_ _5477_/Q _5381_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3821_/A sky130_fd_sc_hd__mux2_1
XFILLER_177_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3751_ _4030_/A _3751_/B vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__nor2_2
XFILLER_229_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2702_ _5622_/Q _2652_/X _2700_/X _2701_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2702_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_229_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3682_ _3683_/A _3683_/B _4076_/B vssd1 vssd1 vccd1 vccd1 _4278_/B sky130_fd_sc_hd__and3_2
X_5421_ _5441_/CLK _5421_/D vssd1 vssd1 vccd1 vccd1 _5421_/Q sky130_fd_sc_hd__dfxtp_1
X_2633_ _2681_/A _2682_/A _2761_/B vssd1 vssd1 vccd1 vccd1 _2634_/A sky130_fd_sc_hd__or3_1
Xoutput203 _2650_/Y vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[15] sky130_fd_sc_hd__buf_2
XANTENNA__3724__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5352_ _5721_/CLK _5352_/D vssd1 vssd1 vccd1 vccd1 _5352_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4600__A _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4303_ _4303_/A _4303_/B vssd1 vssd1 vccd1 vccd1 _4303_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5283_ _5292_/A _5283_/B vssd1 vssd1 vccd1 vccd1 _5284_/A sky130_fd_sc_hd__and2_1
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4234_ _4454_/B _4234_/B vssd1 vssd1 vccd1 vccd1 _4234_/Y sky130_fd_sc_hd__nand2_1
X_4165_ _4454_/D _4121_/X _4159_/X _4164_/Y vssd1 vssd1 vccd1 vccd1 _4165_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5229__A0 _5527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3116_ _3116_/A vssd1 vssd1 vccd1 vccd1 _3116_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2774__B _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4096_ _4096_/A vssd1 vssd1 vccd1 vccd1 _4097_/A sky130_fd_sc_hd__inv_2
XANTENNA__4047__A _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3047_ _2852_/A _3027_/X _3343_/C vssd1 vssd1 vccd1 vccd1 _3047_/X sky130_fd_sc_hd__a21o_1
XFILLER_270_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4452__A1 _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4204__A1 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4998_ _4998_/A vssd1 vssd1 vccd1 vccd1 _5681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_210_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3949_ _3948_/B _3947_/X _3948_/Y _3965_/A vssd1 vssd1 vccd1 vccd1 _3949_/X sky130_fd_sc_hd__a211o_1
XFILLER_23_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2766__A1 _5615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3963__A0 _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5619_ _5653_/CLK _5619_/D vssd1 vssd1 vccd1 vccd1 _5619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3715__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3191__A1 _5636_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5509__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2668__C _5657_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_278_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4140__B1 _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5659__CLK _5659_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5060__B _5060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_i_clk clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5738_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4746__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4404__B _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2850__D _2850_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output182_A _5480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3706__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3182__A1 _5554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3036__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4682__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5251__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4434__A1 _4454_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4921_ _5647_/Q _4947_/B vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__or2_1
XFILLER_64_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2700__B_N _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4852_ _5618_/Q _4856_/A vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__or2_1
XFILLER_220_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3803_ _3532_/X _3780_/A _3791_/X _3802_/X vssd1 vssd1 vccd1 vccd1 _5468_/D sky130_fd_sc_hd__o22a_1
X_4783_ _5588_/Q _4784_/B _4782_/Y _4769_/X vssd1 vssd1 vccd1 vccd1 _5588_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2748__A1 _5617_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3734_ _5670_/Q _3600_/X _3602_/X _5654_/Q vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3665_ _5661_/Q _3600_/X _3602_/X _5645_/Q vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__a22o_1
X_5404_ _5404_/CLK _5404_/D vssd1 vssd1 vccd1 vccd1 _5404_/Q sky130_fd_sc_hd__dfxtp_1
X_3596_ _3596_/A vssd1 vssd1 vccd1 vccd1 _3596_/X sky130_fd_sc_hd__buf_6
XANTENNA__2769__B _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3173__A1 _5665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3173__B2 _5585_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5335_ _5686_/CLK _5335_/D vssd1 vssd1 vccd1 vccd1 _5335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5266_ _5266_/A vssd1 vssd1 vccd1 vccd1 _5731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_272_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4217_ _4483_/A _4213_/X _4215_/X _4216_/X vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__a211o_1
XFILLER_272_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2785__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3380__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5197_ _5193_/X _5196_/Y _5219_/S vssd1 vssd1 vccd1 vccd1 _5198_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__5161__A _5521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4148_ _4132_/A _4232_/B _3613_/X _4128_/B _4128_/A vssd1 vssd1 vccd1 vccd1 _4148_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_28_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_228_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4079_ _4274_/A _4079_/B _4079_/C vssd1 vssd1 vccd1 vccd1 _4280_/B sky130_fd_sc_hd__or3_1
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2951__C _3318_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4728__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4224__B _4307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3164__A1 _5599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3164__B2 _5615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4900__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5481__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A i_req_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5310__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5071__A _5761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2845__D _2967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4416__A1 _4050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3219__A2 _3133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4415__A _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4134__B _4301_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3465__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3450_ _3450_/A vssd1 vssd1 vccd1 vccd1 _5404_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3155__A1 _5645_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3155__B2 _5565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3381_ _3381_/A vssd1 vssd1 vccd1 vccd1 _5371_/D sky130_fd_sc_hd__clkbuf_1
X_5120_ _5131_/A _5131_/B _5156_/B vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_257_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2728__A_N _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5051_ _5528_/Q _5051_/B vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__and2_1
XFILLER_257_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4655__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4002_ _4379_/B _4379_/C vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__nand2_1
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2666__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4958__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5080__A1 _5705_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4904_ _5640_/Q _4897_/B _4903_/Y _4886_/X vssd1 vssd1 vccd1 vccd1 _5640_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_240_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3630__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4216__A2_N _4454_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4835_ _5611_/Q _4822_/B _4834_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5611_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5354__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4766_ _5581_/Q _4797_/B vssd1 vssd1 vccd1 vccd1 _4766_/X sky130_fd_sc_hd__or2_1
XFILLER_267_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3717_ _3732_/A _4418_/A vssd1 vssd1 vccd1 vccd1 _3717_/Y sky130_fd_sc_hd__nand2_2
XFILLER_193_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4697_ _4697_/A _4972_/A vssd1 vssd1 vccd1 vccd1 _4697_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5156__A _5156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3648_ _4229_/A vssd1 vssd1 vccd1 vccd1 _4454_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_146_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3579_ _5555_/Q _2720_/B _2726_/X _2729_/X _3588_/S vssd1 vssd1 vccd1 vccd1 _3579_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3697__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5318_ _5751_/Q _5295_/X _5317_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5751_/D sky130_fd_sc_hd__o211a_1
XFILLER_283_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2746__B_N _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5249_ _5249_/A vssd1 vssd1 vccd1 vccd1 _5726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__S1 _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4401__C _4600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4334__B1 _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5005__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4637__A1 _5527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5377__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2950_ _2949_/Y _2957_/B _3330_/C vssd1 vssd1 vccd1 vccd1 _3308_/D sky130_fd_sc_hd__o21a_1
XFILLER_15_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _5361_/Q _5360_/Q _3304_/A vssd1 vssd1 vccd1 vccd1 _2938_/B sky130_fd_sc_hd__or3_2
XANTENNA__2820__B1 _5331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4620_ _5229_/S _4618_/X _4619_/Y vssd1 vssd1 vccd1 vccd1 _4620_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__4799__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4551_ _5517_/Q _4550_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _4551_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3502_ _3502_/A vssd1 vssd1 vccd1 vccd1 _5430_/D sky130_fd_sc_hd__clkbuf_1
X_4482_ _4484_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _4485_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3433_ _5396_/Q _3048_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3434_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3001_/B _5365_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3365_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5103_ _5707_/Q _5235_/S _5101_/X _5102_/Y vssd1 vssd1 vccd1 vccd1 _5707_/D sky130_fd_sc_hd__a22o_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _5365_/Q vssd1 vssd1 vccd1 vccd1 _3295_/Y sky130_fd_sc_hd__inv_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5034_ _5034_/A vssd1 vssd1 vccd1 vccd1 _5697_/D sky130_fd_sc_hd__clkbuf_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4039__B _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2782__B _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3603__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4818_ _4684_/X _4799_/Y _4817_/X _4815_/X vssd1 vssd1 vccd1 vccd1 _5603_/D sky130_fd_sc_hd__o211a_1
XFILLER_278_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4564__B1 _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4749_ _4974_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4316__A0 _4127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4867__A1 _5624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput58 _3152_/X vssd1 vssd1 vccd1 vccd1 dbg_out[0] sky130_fd_sc_hd__buf_2
Xoutput69 _3157_/X vssd1 vssd1 vccd1 vccd1 dbg_out[1] sky130_fd_sc_hd__buf_2
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3134__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5044__A1 _4457_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3358__A1 _5362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4858__A1 _5620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3080_ _5403_/Q _3079_/B _3011_/A vssd1 vssd1 vccd1 vccd1 _3080_/X sky130_fd_sc_hd__o21ba_1
XFILLER_153_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4086__A2 _4239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3294__B1 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5035__A1 _4490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _5524_/Q _3923_/A _3981_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5524_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2933_ _5359_/Q _3330_/C _3775_/C vssd1 vssd1 vccd1 vccd1 _2934_/B sky130_fd_sc_hd__and3_1
X_5721_ _5721_/CLK _5721_/D vssd1 vssd1 vccd1 vccd1 _5721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5652_ _5654_/CLK _5652_/D vssd1 vssd1 vccd1 vccd1 _5652_/Q sky130_fd_sc_hd__dfxtp_2
X_2864_ _5457_/Q _5406_/Q vssd1 vssd1 vccd1 vccd1 _2865_/C sky130_fd_sc_hd__nor2_1
XANTENNA__4603__A _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4603_ _5771_/A vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__inv_2
XFILLER_248_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5583_ _5747_/CLK _5583_/D vssd1 vssd1 vccd1 vccd1 _5583_/Q sky130_fd_sc_hd__dfxtp_2
X_2795_ _5409_/Q vssd1 vssd1 vccd1 vccd1 _2849_/S sky130_fd_sc_hd__buf_4
XFILLER_190_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4534_ _4552_/C vssd1 vssd1 vccd1 vccd1 _4534_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4465_ _4463_/Y _4464_/X _4483_/A vssd1 vssd1 vccd1 vccd1 _4465_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4849__A1 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3416_ _3416_/A vssd1 vssd1 vccd1 vccd1 _5387_/D sky130_fd_sc_hd__clkbuf_1
X_4396_ _4396_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3347_ _5357_/Q _5356_/Q _3345_/Y _3346_/Y vssd1 vssd1 vccd1 vccd1 _5356_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5542__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3307_/A _3775_/B _3308_/A vssd1 vssd1 vccd1 vccd1 _3278_/Y sky130_fd_sc_hd__o21ai_1
X_5017_ _5017_/A vssd1 vssd1 vccd1 vccd1 _5689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__A1 _5132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3037__B1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3588__A1 _5319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3828__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4232__B _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3129__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3760__A1 _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5063__B _5462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_276_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input21_A i_mem_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4068__A2 _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3799__A _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4407__B _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3028__B1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__C1 _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3579__A1 _5555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3594__A4 _4466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5415__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3200__B1 _3149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5565__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3473__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5254__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4250_ _4300_/S _4250_/B vssd1 vssd1 vccd1 vccd1 _4250_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3201_ _5638_/Q _3143_/A _3145_/A _3200_/X vssd1 vssd1 vccd1 vccd1 _3201_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4700__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4181_ _4300_/S _4178_/X _4180_/Y _4468_/A vssd1 vssd1 vccd1 vccd1 _4181_/X sky130_fd_sc_hd__o211a_1
XFILLER_67_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2711__C1 _2710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3132_ input3/X input2/X input1/X vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__and3b_4
X_3063_ _4590_/B _3063_/B vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__or2_1
XFILLER_82_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_250_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3965_ _3965_/A _3965_/B vssd1 vssd1 vccd1 vccd1 _3965_/X sky130_fd_sc_hd__or2_1
XFILLER_250_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5704_ _5716_/CLK _5704_/D vssd1 vssd1 vccd1 vccd1 _5704_/Q sky130_fd_sc_hd__dfxtp_1
X_2916_ _3281_/A _3277_/A vssd1 vssd1 vccd1 vccd1 _3307_/A sky130_fd_sc_hd__and2_2
XANTENNA__4333__A _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3896_ _5503_/Q _3908_/B _3893_/A vssd1 vssd1 vccd1 vccd1 _3896_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4519__B1 _4529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5635_ _5653_/CLK _5635_/D vssd1 vssd1 vccd1 vccd1 _5635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2847_ input33/X _5428_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2850_/B sky130_fd_sc_hd__mux2_2
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4987__B _4987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5566_ _5674_/CLK _5566_/D vssd1 vssd1 vccd1 vccd1 _5566_/Q sky130_fd_sc_hd__dfxtp_4
X_2778_ _4523_/B vssd1 vssd1 vccd1 vccd1 _2778_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3742__B2 _5607_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4517_ _4533_/C _4527_/C vssd1 vssd1 vccd1 vccd1 _4517_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3383__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5497_ _5741_/CLK _5497_/D vssd1 vssd1 vccd1 vccd1 _5497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4448_ _4466_/A _4415_/A _4373_/A vssd1 vssd1 vccd1 vccd1 _4448_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4379_ _5445_/Q _4379_/B _4379_/C vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__and3_1
XFILLER_258_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5247__A1 _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_273_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4470__A2 _4449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4708__A1_N input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5438__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5588__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4897__B _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2698__A _5670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4143__D1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4694__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4418__A _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5013__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4997__A0 _5681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4153__A _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3750_ _4182_/B _3749_/X _4276_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ _2771_/A _2771_/B _5654_/Q _2806_/A vssd1 vssd1 vccd1 vccd1 _2701_/X sky130_fd_sc_hd__and4b_1
XFILLER_229_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3972__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3681_ _5529_/Q _5466_/Q vssd1 vssd1 vccd1 vccd1 _4076_/B sky130_fd_sc_hd__and2_1
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5420_ _5441_/CLK _5420_/D vssd1 vssd1 vccd1 vccd1 _5420_/Q sky130_fd_sc_hd__dfxtp_1
X_2632_ _5345_/Q vssd1 vssd1 vccd1 vccd1 _2761_/B sky130_fd_sc_hd__buf_2
XFILLER_64_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3724__A1 _5637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput204 _2785_/Y vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[1] sky130_fd_sc_hd__buf_2
X_5351_ _5716_/CLK _5351_/D vssd1 vssd1 vccd1 vccd1 _5351_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4600__B _4600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4302_ _4059_/B _4379_/C _4302_/S vssd1 vssd1 vccd1 vccd1 _4303_/B sky130_fd_sc_hd__mux2_1
X_5282_ _5737_/Q _5772_/A _5285_/S vssd1 vssd1 vccd1 vccd1 _5283_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4233_ _4231_/S _4071_/B _4232_/X vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__o21ai_1
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _2954_/X _4059_/C _4163_/X vssd1 vssd1 vccd1 vccd1 _4164_/Y sky130_fd_sc_hd__a21oi_1
X_3115_ _5705_/Q _5713_/Q _4651_/S vssd1 vssd1 vccd1 vccd1 _3116_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4095_ _4034_/A _4092_/Y _4101_/B vssd1 vssd1 vccd1 vccd1 _4213_/B sky130_fd_sc_hd__a21o_1
XANTENNA__2774__C _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3232__A _5461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3046_ _3085_/A _3053_/C _3046_/C vssd1 vssd1 vccd1 vccd1 _3046_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4047__B _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _5681_/Q _5335_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5730__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4063__A _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3948_ _3948_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _3948_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2766__A2 _2652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3879_ _3893_/A _3879_/B vssd1 vssd1 vccd1 vccd1 _3880_/A sky130_fd_sc_hd__and2_1
XFILLER_136_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5618_ _5650_/CLK _5618_/D vssd1 vssd1 vccd1 vccd1 _5618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3715__A1 _5642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5549_ _5674_/CLK _5549_/D vssd1 vssd1 vccd1 vccd1 _5549_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_151_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3191__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2668__D _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4676__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4140__A1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2687__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2684__C _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3651__B1 _3602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3403__A0 _2852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3954__A1 _5517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3706__A1 _5576_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3706__B2 _5592_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3317__A _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3182__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_338 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5603__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2875__B _5361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4920_ _4658_/X _4912_/Y _4919_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5646_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3642__B1 _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2996__A2 _2850_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4851_ _4674_/X _4836_/Y _4850_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5617_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_220_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3802_ _3802_/A _3802_/B _3802_/C _3802_/D vssd1 vssd1 vccd1 vccd1 _3802_/X sky130_fd_sc_hd__or4_2
X_4782_ _4970_/A _4784_/B vssd1 vssd1 vccd1 vccd1 _4782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2748__A2 _2652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3733_ _3726_/Y _3732_/Y _4231_/S vssd1 vssd1 vccd1 vccd1 _3733_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3926__S _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3664_ _4231_/S vssd1 vssd1 vccd1 vccd1 _4449_/S sky130_fd_sc_hd__buf_4
XFILLER_256_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5403_ _5404_/CLK _5403_/D vssd1 vssd1 vccd1 vccd1 _5403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3595_ _4128_/B vssd1 vssd1 vccd1 vccd1 _4469_/C sky130_fd_sc_hd__buf_2
XFILLER_133_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2769__C _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3173__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5334_ _5686_/CLK _5334_/D vssd1 vssd1 vccd1 vccd1 _5334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5265_ _5292_/A _5265_/B vssd1 vssd1 vccd1 vccd1 _5266_/A sky130_fd_sc_hd__and2_1
X_4216_ _3750_/X _4454_/D _4092_/B _2954_/X vssd1 vssd1 vccd1 vccd1 _4216_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_275_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5196_ _5196_/A _5196_/B vssd1 vssd1 vccd1 vccd1 _5196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_275_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4147_ _4146_/A _4142_/X _4146_/Y _4300_/S vssd1 vssd1 vccd1 vccd1 _4147_/X sky130_fd_sc_hd__a211o_1
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4078_ _3572_/X _4077_/Y _3673_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _4079_/C sky130_fd_sc_hd__o211a_1
X_3029_ _5081_/A _3010_/X _3026_/Y _3028_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3029_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2987__A2 _2852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3836__S _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3137__A _3137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3164__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5626__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4667__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2695__B _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_94 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3624__B1 _3608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3600__A _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4821__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3927__A1 _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3155__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3380_ _3379_/X _5371_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3381_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4104__A1 _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5050_ _5760_/A _5125_/A _5459_/Q vssd1 vssd1 vccd1 vccd1 _5050_/X sky130_fd_sc_hd__a21o_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4001_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__nand2_2
XANTENNA__4655__A2 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2666__A1 _5641_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2666__B2 _5673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2825__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4606__A _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5080__A2 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4903_ _4978_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4903_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3091__A1 _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4834_ _4985_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4834_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4765_ _4646_/X _4761_/Y _4764_/X _4745_/X vssd1 vssd1 vccd1 vccd1 _5580_/D sky130_fd_sc_hd__o211a_1
XFILLER_193_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3716_ _5562_/Q _3596_/X _3713_/X _3715_/X vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__o22a_4
XANTENNA__5649__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4696_ input22/X _4689_/X _4690_/X _4695_/Y vssd1 vssd1 vccd1 vccd1 _4972_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_146_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5156__B _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _4303_/A _3647_/B vssd1 vssd1 vccd1 vccd1 _3647_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_15_i_clk clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5747_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4343__A1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4343__B2 _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3578_ _5480_/Q _3532_/X _3577_/X vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__a21o_4
XANTENNA__2796__A _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5317_ _5317_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__or2_1
XFILLER_248_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_275_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5248_ _5261_/A _5248_/B vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__and2_1
XFILLER_275_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5179_ _5178_/X _5317_/A _5179_/S vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4803__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3082__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4582__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4401__D _4490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4334__B2 _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input51_A i_req_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4098__B1 _4192_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4637__A2 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2648__A1 _5579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3330__A _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__A1_N _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3073__A1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2880_ _5359_/Q _5358_/Q vssd1 vssd1 vccd1 vccd1 _3304_/A sky130_fd_sc_hd__nand2_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4573__A1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4550_ _5307_/A _4499_/B _4550_/S vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3501_ _5430_/Q input36/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3502_/A sky130_fd_sc_hd__mux2_1
XFILLER_183_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4481_ _5530_/Q _4458_/A _4480_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5530_/D sky130_fd_sc_hd__o211a_1
X_3432_ _3432_/A vssd1 vssd1 vccd1 vccd1 _5395_/D sky130_fd_sc_hd__clkbuf_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3363_/A vssd1 vssd1 vccd1 vccd1 _5364_/D sky130_fd_sc_hd__clkbuf_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _3790_/X _3943_/A _5235_/S vssd1 vssd1 vccd1 vccd1 _5102_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_257_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _5365_/Q _3292_/X _3293_/X _5334_/Q vssd1 vssd1 vccd1 vccd1 _5334_/D sky130_fd_sc_hd__a2bb2o_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5697_/Q _4362_/A _5135_/S vssd1 vssd1 vccd1 vccd1 _5034_/A sky130_fd_sc_hd__mux2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3836__A0 _5485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_382 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3240__A _5475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2782__C _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3064__A1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5471__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4817_ _5603_/Q _4819_/A vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__or2_1
XFILLER_178_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3386__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4071__A _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4748_ _5573_/Q _4747_/B _4747_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5573_/D sky130_fd_sc_hd__o211a_1
X_4679_ _4679_/A vssd1 vssd1 vccd1 vccd1 _4679_/X sky130_fd_sc_hd__buf_4
XANTENNA__4316__A1 _4148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4867__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput59 _3202_/X vssd1 vssd1 vccd1 vccd1 dbg_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3134__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4252__A0 _3717_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_304 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2718__A_N _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4004__B1 _3584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4858__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5016__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5344__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3818__A0 _5476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4156__A _4306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5494__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _3990_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _3981_/X sky130_fd_sc_hd__or2_1
X_5720_ _5721_/CLK _5720_/D vssd1 vssd1 vccd1 vccd1 _5720_/Q sky130_fd_sc_hd__dfxtp_1
X_2932_ _3791_/A vssd1 vssd1 vccd1 vccd1 _3293_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4794__A1 _5593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5651_ _5653_/CLK _5651_/D vssd1 vssd1 vccd1 vccd1 _5651_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2736__B_N _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2863_ _5331_/B vssd1 vssd1 vccd1 vccd1 _2863_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4602_ _4599_/Y _4601_/X _4532_/X vssd1 vssd1 vccd1 vccd1 _4602_/Y sky130_fd_sc_hd__a21oi_1
X_5582_ _5667_/CLK _5582_/D vssd1 vssd1 vccd1 vccd1 _5582_/Q sky130_fd_sc_hd__dfxtp_4
X_2794_ _5355_/Q vssd1 vssd1 vccd1 vccd1 _2794_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4533_ _5763_/A _5081_/A _4533_/C _5760_/A vssd1 vssd1 vccd1 vccd1 _4552_/C sky130_fd_sc_hd__and4_1
XANTENNA__3934__S _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4464_ _4419_/A _4419_/B _4483_/B _4438_/A _4408_/A vssd1 vssd1 vccd1 vccd1 _4464_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_171_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4849__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3415_ _2845_/A _5387_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3416_/A sky130_fd_sc_hd__mux2_1
XFILLER_264_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4395_ _4394_/Y _4177_/Y _4373_/Y _4141_/Y _4469_/D _4449_/S vssd1 vssd1 vccd1 vccd1
+ _4395_/X sky130_fd_sc_hd__mux4_1
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ _4987_/A _3346_/B vssd1 vssd1 vccd1 vccd1 _3346_/Y sky130_fd_sc_hd__nor2_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__A0 _5472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3277_ _3277_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3308_/C sky130_fd_sc_hd__nor2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5016_ _5689_/Q _5015_/Y _5030_/S vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3285__A1 _5361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3037__A1 _2840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3129__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5367__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3145__A _3145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_264_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3799__B _3799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3276__A1 _3308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3276__B2 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input14_A i_mem_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3028__A1 _2850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3579__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4776__A1 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3200__B2 _5574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2878__B _5362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output82_A _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3200_ _5654_/Q _3147_/A _3149_/A _5574_/Q vssd1 vssd1 vccd1 vccd1 _3200_/X sky130_fd_sc_hd__a22o_1
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4180_ _4300_/S _4180_/B vssd1 vssd1 vccd1 vccd1 _4180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3131_ _3131_/A vssd1 vssd1 vccd1 vccd1 _3131_/X sky130_fd_sc_hd__buf_4
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_282_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3062_ _3061_/Y _2850_/A _3089_/A vssd1 vssd1 vccd1 vccd1 _3062_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4216__B1 _4092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2833__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__A1 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3964_ _3963_/X _5313_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3965_/B sky130_fd_sc_hd__mux2_1
X_5703_ _5724_/CLK _5703_/D vssd1 vssd1 vccd1 vccd1 _5703_/Q sky130_fd_sc_hd__dfxtp_1
X_2915_ _5451_/Q _5486_/D _2914_/X vssd1 vssd1 vccd1 vccd1 _5451_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3895_ _5319_/A vssd1 vssd1 vccd1 vccd1 _3895_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4519__A1 _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5634_ _5653_/CLK _5634_/D vssd1 vssd1 vccd1 vccd1 _5634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2846_ input41/X _5435_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2850_/A sky130_fd_sc_hd__mux2_2
XFILLER_136_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5565_ _5674_/CLK _5565_/D vssd1 vssd1 vccd1 vccd1 _5565_/Q sky130_fd_sc_hd__dfxtp_4
X_2777_ _5550_/Q _2720_/B _2770_/X _2776_/X vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__o22ai_4
XFILLER_275_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3742__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4516_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4634_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_2_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5496_ _5741_/CLK _5496_/D vssd1 vssd1 vccd1 vccd1 _5496_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2950__B1 _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4447_ _4176_/Y _4140_/Y _4447_/S vssd1 vssd1 vccd1 vccd1 _4447_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ _3617_/A _4305_/B _4224_/X vssd1 vssd1 vccd1 vccd1 _4378_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_258_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input6_A i_mem_ack vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3329_ _5347_/Q _3780_/A _2934_/X vssd1 vssd1 vccd1 vccd1 _5347_/D sky130_fd_sc_hd__o21a_1
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_9 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_258_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_233_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4207__B1 _4271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4758__A1 _5578_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__A _5514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5183__A1 _5523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3574__S _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3194__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4930__A1 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2698__B _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output120_A _5552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3749__S _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5532__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2700_ _2806_/A _2771_/A _2771_/B _5590_/Q vssd1 vssd1 vccd1 vccd1 _2700_/X sky130_fd_sc_hd__and4bb_1
X_3680_ _3673_/A _3673_/B _4076_/A vssd1 vssd1 vccd1 vccd1 _3683_/B sky130_fd_sc_hd__a21o_1
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ _5346_/Q vssd1 vssd1 vccd1 vccd1 _2682_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3484__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5265__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3185__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3724__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5350_ _5716_/CLK _5350_/D vssd1 vssd1 vccd1 vccd1 _5350_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput205 _2778_/Y vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_57_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5682__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4301_ _4118_/B _3717_/Y _4301_/S vssd1 vssd1 vccd1 vccd1 _4301_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5281_ _5281_/A vssd1 vssd1 vccd1 vccd1 _5736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_245_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4232_ _4301_/S _4232_/B vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__or2_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2828__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4163_ _2904_/X _4052_/A _4403_/B _2936_/X _4162_/X vssd1 vssd1 vccd1 vccd1 _4163_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3114_ _3114_/A vssd1 vssd1 vccd1 vccd1 _3114_/X sky130_fd_sc_hd__clkbuf_1
X_4094_ _4034_/A _4093_/Y _4040_/X vssd1 vssd1 vccd1 vccd1 _4101_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__2774__D _5630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3232__B _4988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3045_ _5396_/Q _3045_/B vssd1 vssd1 vccd1 vccd1 _3046_/C sky130_fd_sc_hd__nor2_1
XFILLER_208_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3660__A1 _5551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4996_ _4996_/A vssd1 vssd1 vccd1 vccd1 _5680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_211_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3947_ _4552_/B _5729_/Q _5329_/A vssd1 vssd1 vccd1 vccd1 _3947_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3878_ _5497_/Q _5307_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3879_/B sky130_fd_sc_hd__mux2_1
X_5617_ _5650_/CLK _5617_/D vssd1 vssd1 vccd1 vccd1 _5617_/Q sky130_fd_sc_hd__dfxtp_4
X_2829_ _2829_/A _2829_/B vssd1 vssd1 vccd1 vccd1 _3003_/C sky130_fd_sc_hd__nand2_1
XANTENNA__2799__A _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3394__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3176__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3715__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5548_ _5747_/CLK _5548_/D vssd1 vssd1 vccd1 vccd1 _5548_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_151_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5479_ _5741_/CLK _5479_/D vssd1 vssd1 vccd1 vccd1 _5479_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4140__A2 _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5405__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3142__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A1 _5662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__B2 _5646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5555__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_224 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4701__B _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3706__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2914__B1 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output168_A _3082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4667__A0 _5708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5024__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5092__B1 _5706_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__A1 _5650_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3642__B2 _5602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4850_ _5617_/Q _4856_/A vssd1 vssd1 vccd1 vccd1 _4850_/X sky130_fd_sc_hd__or2_1
XFILLER_60_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3801_ _3775_/A _2937_/Y _2951_/B _2934_/B vssd1 vssd1 vccd1 vccd1 _3802_/D sky130_fd_sc_hd__a211o_1
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4781_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4784_/B sky130_fd_sc_hd__buf_4
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3732_ _3732_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _3732_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3663_ _4302_/S vssd1 vssd1 vccd1 vccd1 _4231_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__3158__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5402_ _5492_/CLK _5402_/D vssd1 vssd1 vccd1 vccd1 _5402_/Q sky130_fd_sc_hd__dfxtp_1
X_3594_ _3747_/A _4067_/A _4379_/B _4466_/B _5454_/Q vssd1 vssd1 vccd1 vccd1 _4128_/B
+ sky130_fd_sc_hd__o41ai_4
XFILLER_256_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2769__D _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5333_ _5686_/CLK _5333_/D vssd1 vssd1 vccd1 vccd1 _5333_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3942__S _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5428__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5264_ _5731_/Q _5766_/A _5285_/S vssd1 vssd1 vccd1 vccd1 _5265_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4215_ _2904_/X _4091_/B _4214_/X _4096_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4215_/X
+ sky130_fd_sc_hd__a221o_1
X_5195_ _5753_/Q _3840_/X _5194_/X vssd1 vssd1 vccd1 vccd1 _5196_/B sky130_fd_sc_hd__a21oi_1
XFILLER_228_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3243__A _4988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ _4146_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5578__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4077_ _5529_/Q _5466_/Q vssd1 vssd1 vccd1 vccd1 _4077_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3618__D1 _3549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5083__B1 _5051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3028_ _2850_/B _3027_/X _3343_/C vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4979_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4979_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3397__A0 _2840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4802__A _5596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5310__A1 _2743_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2695__C _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_219_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4683__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5074__B1 _5125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3624__A1 _5569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3624__B2 _5585_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3388__A0 _2840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2886__B _5360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4104__A2 _4105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3063__A _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ _4059_/A _4000_/B vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__nor2_2
XFILLER_284_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2666__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5065__B1 _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ _5639_/Q _4897_/B _4901_/Y _4886_/X vssd1 vssd1 vccd1 vccd1 _5639_/D sky130_fd_sc_hd__o211a_1
X_4833_ _5610_/Q _4822_/B _4832_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5610_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2774__A_N _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2841__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4764_ _5580_/Q _4797_/B vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__or2_1
XFILLER_193_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3715_ _5642_/Q _3605_/X _3606_/X _3714_/X vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__a211o_1
XFILLER_186_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4695_ _5713_/Q vssd1 vssd1 vccd1 vccd1 _4695_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3238__A _5479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3646_ _4161_/B _4071_/B _4302_/S vssd1 vssd1 vccd1 vccd1 _3647_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4343__A2 _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3577_ _5558_/Q _2720_/B _2699_/X _2702_/X _3588_/S vssd1 vssd1 vccd1 vccd1 _3577_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5316_ _5750_/Q _5295_/X _5315_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5750_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4069__A _4467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5247_ _5726_/Q _4533_/C _5253_/S vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3303__B1 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _4490_/B _5177_/Y _5200_/B vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__mux2_1
XFILLER_263_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4129_ _4129_/A vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4532__A _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3148__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4678__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5743__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input44_A i_req_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2647__A_N _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2648__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3058__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output200_A _5321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4270__A1 _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3073__A2 _3063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4161__B _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3500_ _3500_/A vssd1 vssd1 vccd1 vccd1 _5429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4480_ _4482_/B _4485_/A _4458_/Y _4479_/Y vssd1 vssd1 vccd1 vccd1 _4480_/X sky130_fd_sc_hd__a211o_1
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3431_ _5395_/Q _3043_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3432_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3492__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _3003_/A _5364_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3363_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4730__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5101_ _4537_/B _5156_/B _5109_/A _5100_/Y _3790_/X vssd1 vssd1 vccd1 vccd1 _5101_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3293_/A vssd1 vssd1 vccd1 vccd1 _3293_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_253_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5032_ _5032_/A vssd1 vssd1 vccd1 vccd1 _5135_/S sky130_fd_sc_hd__buf_4
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2836__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_394 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_253_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_213_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3240__B _5474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2782__D _5597_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5616__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4816_ _4679_/X _4799_/Y _4814_/X _4815_/X vssd1 vssd1 vccd1 vccd1 _5602_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4549__C1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5210__A0 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4071__B _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4747_ _4972_/A _4747_/B vssd1 vssd1 vccd1 vccd1 _4747_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4678_ _5710_/Q _4677_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4316__A2 _4149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3629_ _5568_/Q _3607_/A _3608_/A _5584_/Q vssd1 vssd1 vccd1 vccd1 _3629_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_276_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4527__A _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5122__S _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4252__A1 _4307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__A1 _5479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4960__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3606__A _3606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5093__A _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4437__A _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3341__A _5300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5639__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_i_clk clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5665_/CLK sky130_fd_sc_hd__clkbuf_16
X_3980_ _3979_/X _5321_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__mux2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _3800_/C _3791_/B _3318_/A _5241_/B vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__or4_1
XFILLER_250_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4794__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5268__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4172__A _4396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5650_ _5650_/CLK _5650_/D vssd1 vssd1 vccd1 vccd1 _5650_/Q sky130_fd_sc_hd__dfxtp_2
X_2862_ _3451_/S vssd1 vssd1 vccd1 vccd1 _3435_/S sky130_fd_sc_hd__buf_4
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4601_ _4600_/A _3895_/Y _4600_/Y _5294_/A vssd1 vssd1 vccd1 vccd1 _4601_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_29_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5528_/CLK sky130_fd_sc_hd__clkbuf_16
X_5581_ _5747_/CLK _5581_/D vssd1 vssd1 vccd1 vccd1 _5581_/Q sky130_fd_sc_hd__dfxtp_4
X_2793_ _2793_/A vssd1 vssd1 vccd1 vccd1 _5067_/B sky130_fd_sc_hd__buf_6
X_4532_ _4634_/A vssd1 vssd1 vccd1 vccd1 _4532_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4463_ _4430_/Y _4420_/B _4422_/B _4422_/A vssd1 vssd1 vccd1 vccd1 _4463_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3414_ _3414_/A vssd1 vssd1 vccd1 vccd1 _5386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_264_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4394_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4394_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_258_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3345_ _3345_/A vssd1 vssd1 vccd1 vccd1 _3345_/Y sky130_fd_sc_hd__inv_2
XFILLER_285_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3276_ _3308_/A _2943_/C _2957_/B _3775_/A vssd1 vssd1 vccd1 vccd1 _3802_/B sky130_fd_sc_hd__a22o_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_358 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _5015_/Y sky130_fd_sc_hd__inv_2
XFILLER_280_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4347__A _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3285__A2 _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4785__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3397__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3129__C input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4810__A _5600_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4942__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_i_clk_A i_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_254_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3276__A2 _2943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4225__A1 _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4776__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2787__A1 _5628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2787__B2 _5644_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output198_A _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3736__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3200__A2 _3147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output75_A _5769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2711__A1 _5621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3130_ _3130_/A vssd1 vssd1 vccd1 vccd1 _3131_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5461__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2894__B _5363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_227_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4167__A _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3061_ _3069_/C _3061_/B vssd1 vssd1 vccd1 vccd1 _3061_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4464__A1 _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3071__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4464__B2 _4408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4216__B2 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3963_ _5768_/A _5733_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3975__A0 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2914_ _3775_/A _2943_/C _3775_/C _3795_/A vssd1 vssd1 vccd1 vccd1 _2914_/X sky130_fd_sc_hd__a31o_1
X_5702_ _5724_/CLK _5702_/D vssd1 vssd1 vccd1 vccd1 _5702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3894_ _3894_/A vssd1 vssd1 vccd1 vccd1 _5502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_259_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5633_ _5667_/CLK _5633_/D vssd1 vssd1 vccd1 vccd1 _5633_/Q sky130_fd_sc_hd__dfxtp_2
X_2845_ _2845_/A _2845_/B _2845_/C _2967_/A vssd1 vssd1 vccd1 vccd1 _2851_/B sky130_fd_sc_hd__or4_1
XFILLER_12_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3727__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4924__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5564_ _5747_/CLK _5564_/D vssd1 vssd1 vccd1 vccd1 _5564_/Q sky130_fd_sc_hd__dfxtp_4
X_2776_ _2771_/Y _2772_/X _2773_/X _2774_/X _2775_/X vssd1 vssd1 vccd1 vccd1 _2776_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4515_ _5294_/A _4513_/X _4514_/X vssd1 vssd1 vccd1 vccd1 _4515_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_275_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5495_ _5741_/CLK _5495_/D vssd1 vssd1 vccd1 vccd1 _5495_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2788__C _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3246__A _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4446_ _2904_/X _4405_/B _4440_/A _2954_/X _4445_/X vssd1 vssd1 vccd1 vccd1 _4455_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_208_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4152__A0 _4148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4377_ _4377_/A vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2702__A1 _5622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3328_ _2771_/A _3780_/A _3327_/X vssd1 vssd1 vccd1 vccd1 _5346_/D sky130_fd_sc_hd__o21a_2
XFILLER_258_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3259_ _5528_/Q _3265_/A _5530_/Q vssd1 vssd1 vccd1 vccd1 _3259_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4077__A _5529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4207__B2 _4454_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4758__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5334__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3194__A1 _5605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3194__B2 _5621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4930__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2698__C _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5484__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4143__B1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4694__A1 _5556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4446__A1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4446__B2 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output113_A _5560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_269 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4906__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2630_ _5344_/Q vssd1 vssd1 vccd1 vccd1 _2681_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3185__A1 _5651_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3185__B2 _5571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput206 _2768_/Y vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__3066__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4300_ _4299_/X _4220_/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4428_/B sky130_fd_sc_hd__mux2_1
XFILLER_160_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5280_ _5292_/A _5280_/B vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__and2_1
XFILLER_4_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4231_ _4063_/A _4024_/B _4231_/S vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4162_ _2919_/X _4050_/A _4415_/A _4333_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4162_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4609__B _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3113_ _5704_/Q _5712_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3114_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4093_ _4161_/B vssd1 vssd1 vccd1 vccd1 _4093_/Y sky130_fd_sc_hd__inv_2
XFILLER_261_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3044_ _5396_/Q _3045_/B vssd1 vssd1 vccd1 vccd1 _3053_/C sky130_fd_sc_hd__and2_1
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2844__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3660__A2 _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5357__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4995_ _5680_/Q _5334_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3946_ _5515_/Q _3923_/X _3944_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5515_/D sky130_fd_sc_hd__o211a_1
XFILLER_23_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3877_ _5496_/Q _3874_/B _3876_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _5496_/D sky130_fd_sc_hd__o211a_1
XFILLER_164_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2828_ input49/X _5413_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _2829_/B sky130_fd_sc_hd__mux2_2
X_5616_ _5667_/CLK _5616_/D vssd1 vssd1 vccd1 vccd1 _5616_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3176__A1 _5633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5547_ _5665_/CLK _5547_/D vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__dfxtp_4
X_2759_ _5552_/Q _2720_/B _2755_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__o22ai_4
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5478_ _5741_/CLK _5478_/D vssd1 vssd1 vccd1 vccd1 _5478_/Q sky130_fd_sc_hd__dfxtp_4
X_4429_ _4428_/A _4471_/S _4375_/B _4427_/Y _4428_/Y vssd1 vssd1 vccd1 vccd1 _4429_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__5322__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4676__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3142__C input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A2 _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3167__A1 _5551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2914__A1 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4721__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3875__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5092__B2 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5040__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__A2 _3602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3800_ _3800_/A _3800_/B _3800_/C _3800_/D vssd1 vssd1 vccd1 vccd1 _3802_/C sky130_fd_sc_hd__or4_1
X_4780_ _4684_/X _4761_/Y _4779_/X _4769_/X vssd1 vssd1 vccd1 vccd1 _5587_/D sky130_fd_sc_hd__o211a_1
XFILLER_220_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3731_ _5556_/Q _3596_/X _3727_/X _3730_/X vssd1 vssd1 vccd1 vccd1 _4132_/B sky130_fd_sc_hd__o22a_4
XFILLER_146_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4180__A _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3662_ _4083_/B _4024_/B _4272_/S vssd1 vssd1 vccd1 vccd1 _3662_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3158__A1 _5662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3158__B2 _5582_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5401_ _5492_/CLK _5401_/D vssd1 vssd1 vccd1 vccd1 _5401_/Q sky130_fd_sc_hd__dfxtp_1
X_3593_ _4306_/A _4229_/A _4301_/S _4326_/A _4030_/A vssd1 vssd1 vccd1 vccd1 _4466_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5332_ _5332_/A vssd1 vssd1 vccd1 vccd1 _5757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2839__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5304__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5263_ _5263_/A vssd1 vssd1 vccd1 vccd1 _5292_/A sky130_fd_sc_hd__buf_2
XFILLER_141_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4214_ _2936_/X _4132_/B _2919_/X vssd1 vssd1 vccd1 vccd1 _4214_/X sky130_fd_sc_hd__a21o_1
XFILLER_141_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5194_ _5524_/Q _3932_/B _3864_/C _5504_/Q _5053_/X vssd1 vssd1 vccd1 vccd1 _5194_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_272_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4145_ _4143_/X _4144_/X _4447_/S vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__mux2_1
XFILLER_228_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4076_ _4076_/A _4076_/B vssd1 vssd1 vccd1 vccd1 _4079_/B sky130_fd_sc_hd__nor2_2
XFILLER_283_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5083__B2 _5530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3027_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3027_/X sky130_fd_sc_hd__buf_2
XANTENNA__4355__A _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4978_ _4978_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_211_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4594__B1 _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4802__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3929_ _5512_/Q _3923_/X _3928_/X _3848_/X vssd1 vssd1 vccd1 vccd1 _5512_/D sky130_fd_sc_hd__o211a_1
XFILLER_137_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3321__A1 _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2695__D _5606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3321__B2 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5522__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5074__A1 _5513_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5074__B2 _5761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3624__A2 _3607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4821__A1 _5604_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5672__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4204__S _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output180_A _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_269_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5035__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3312__A1 _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3063__B _3063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5065__B2 _4500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4901_ _4976_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4901_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2823__B1 _3458_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4903__A _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4832_ _4983_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4832_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4576__A0 _5520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4763_ _4781_/A vssd1 vssd1 vccd1 vccd1 _4797_/B sky130_fd_sc_hd__buf_4
XFILLER_267_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3714_ _5578_/Q _3607_/X _3608_/X _5594_/Q vssd1 vssd1 vccd1 vccd1 _3714_/X sky130_fd_sc_hd__a22o_1
X_4694_ _5556_/Q _4697_/A _4693_/Y _4670_/X vssd1 vssd1 vccd1 vccd1 _5556_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3238__B _5481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3645_ _5554_/Q _3596_/A _3642_/X _3644_/X vssd1 vssd1 vccd1 vccd1 _4071_/B sky130_fd_sc_hd__o22a_4
XFILLER_20_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_283_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3576_ _4419_/A _4408_/A _4050_/A vssd1 vssd1 vccd1 vccd1 _3590_/A sky130_fd_sc_hd__or3_1
XFILLER_283_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5315_ _5315_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__or2_1
XANTENNA__5545__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5246_ _5246_/A vssd1 vssd1 vccd1 vccd1 _5725_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4069__B _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177_ _5182_/A _5177_/B vssd1 vssd1 vccd1 vccd1 _5177_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_256_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4128_ _4128_/A _4128_/B _4128_/C vssd1 vssd1 vccd1 vccd1 _4129_/A sky130_fd_sc_hd__and3_1
XANTENNA__5695__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4059_ _4059_/A _4059_/B _4059_/C vssd1 vssd1 vccd1 vccd1 _4060_/B sky130_fd_sc_hd__or3_1
XFILLER_216_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3067__B1 _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4803__A1 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2814__A0 _5684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3148__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4098__A2 _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input37_A i_req_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3330__C _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5418__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_230_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3339__A _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3230__B1 _3458_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3781__A1 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5568__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3430_ _3430_/A vssd1 vssd1 vccd1 vccd1 _5394_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2897__B _5363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3361_ _3361_/A vssd1 vssd1 vccd1 vccd1 _5363_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _4536_/Y _5087_/Y _5098_/Y _5156_/B vssd1 vssd1 vccd1 vccd1 _5100_/Y sky130_fd_sc_hd__a31oi_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3292_ _5367_/Q _5366_/Q _3791_/A _3292_/D vssd1 vssd1 vccd1 vccd1 _3292_/X sky130_fd_sc_hd__or4_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5031_ _5031_/A vssd1 vssd1 vccd1 vccd1 _5696_/D sky130_fd_sc_hd__clkbuf_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3240__C _5477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4633__A _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4815_/X sky130_fd_sc_hd__buf_6
XFILLER_278_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3249__A _5508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3221__B1 _3145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4746_ _5572_/Q _4747_/B _4744_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5572_/D sky130_fd_sc_hd__o211a_1
XFILLER_193_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4677_ input12/X input19/X _4682_/S vssd1 vssd1 vccd1 vccd1 _4677_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4316__A3 _4150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3628_ _5616_/Q _3597_/A _3598_/A _5600_/Q _3627_/X vssd1 vssd1 vccd1 vccd1 _3628_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4721__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3559_ _5343_/Q _3601_/B _5341_/Q vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__nor3b_4
XFILLER_88_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5229_ _5527_/Q _5228_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _5230_/B sky130_fd_sc_hd__mux2_2
XANTENNA__4808__A _5599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4527__B _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4543__A _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5201__A1 _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4004__A2 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5710__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4692__A1_N input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5093__B _5125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4712__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4718__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3768__S _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2930_ _3799_/A _3317_/B vssd1 vssd1 vccd1 vccd1 _5241_/B sky130_fd_sc_hd__nor2_1
XFILLER_203_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2861_ _5300_/A _3343_/B vssd1 vssd1 vccd1 vccd1 _3451_/S sky130_fd_sc_hd__nor2_4
XANTENNA__5390__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4600_ _4600_/A _4600_/B vssd1 vssd1 vccd1 vccd1 _4600_/Y sky130_fd_sc_hd__nor2_1
XFILLER_248_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3203__B1 _3139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5580_ _5747_/CLK _5580_/D vssd1 vssd1 vccd1 vccd1 _5580_/Q sky130_fd_sc_hd__dfxtp_4
X_2792_ _2786_/X _2787_/X _2790_/X _2791_/X vssd1 vssd1 vccd1 vccd1 _2793_/A sky130_fd_sc_hd__o31a_1
XANTENNA__3754__A1 _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4531_ _5081_/A _4511_/X _3919_/X _4530_/X vssd1 vssd1 vccd1 vccd1 _5534_/D sky130_fd_sc_hd__o211a_1
XFILLER_156_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4462_ _4410_/A _4405_/A _4406_/Y _4409_/A _4322_/A vssd1 vssd1 vccd1 vccd1 _4462_/X
+ sky130_fd_sc_hd__a311o_1
X_3413_ _2835_/B _5386_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3414_/A sky130_fd_sc_hd__mux2_1
X_4393_ _3678_/Y _4255_/C _4392_/X _4043_/B vssd1 vssd1 vccd1 vccd1 _4399_/B sky130_fd_sc_hd__a22o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3344_ _3344_/A vssd1 vssd1 vccd1 vccd1 _5355_/D sky130_fd_sc_hd__clkbuf_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2847__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3275_ _3277_/A _2946_/A _3330_/C _5241_/C vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__a31o_1
XFILLER_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4628__A _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _5014_/A vssd1 vssd1 vccd1 vccd1 _5688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_285_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_213_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5733__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4363__A _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3745__A1 _5559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4729_ _5565_/Q _4759_/B vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__or2_1
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4810__B _4819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4302__S _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5344__D _5344_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4063__B_N _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4225__A2 _4223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3588__S _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2787__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3984__A1 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3736__A1 _5574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3736__B2 _5590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3617__A _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output68_A _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2711__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2894__C _5362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3060_ _5399_/Q _3060_/B vssd1 vssd1 vccd1 vccd1 _3061_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4167__B _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5756__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3672__B1 _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3962_ _5519_/Q _3923_/X _3961_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5519_/D sky130_fd_sc_hd__o211a_1
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701_ _5724_/CLK _5701_/D vssd1 vssd1 vccd1 vccd1 _5701_/Q sky130_fd_sc_hd__dfxtp_1
X_2913_ _3791_/A vssd1 vssd1 vccd1 vccd1 _3795_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_259_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3893_ _3893_/A _3893_/B vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__and2_1
XFILLER_259_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5632_ _5667_/CLK _5632_/D vssd1 vssd1 vccd1 vccd1 _5632_/Q sky130_fd_sc_hd__dfxtp_2
X_2844_ input43/X _5437_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3727__A1 _5668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3727__B2 _5652_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5563_ _5675_/CLK _5563_/D vssd1 vssd1 vccd1 vccd1 _5563_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_275_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2775_ _2727_/C _2775_/B _5646_/Q _2775_/D vssd1 vssd1 vccd1 vccd1 _2775_/X sky130_fd_sc_hd__and4b_1
XANTENNA__3527__A _5468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4514_ _5513_/Q _5459_/Q vssd1 vssd1 vccd1 vccd1 _4514_/X sky130_fd_sc_hd__and2_1
XFILLER_144_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5494_ _5741_/CLK _5494_/D vssd1 vssd1 vccd1 vccd1 _5494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2788__D _5564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4445_ _4418_/A _4333_/A _4444_/X _4419_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4445_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4152__A1 _4149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4376_ _4396_/A _4299_/X _4375_/Y _4347_/A vssd1 vssd1 vccd1 vccd1 _4376_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2702__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3327_ _5368_/Q _3335_/B _3335_/C _5371_/Q _3293_/A vssd1 vssd1 vccd1 vccd1 _3327_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5101__B1 _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3258_ _3265_/A _3255_/X _3256_/X _3265_/B vssd1 vssd1 vccd1 vccd1 _3258_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4077__B _5466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3189_ _5604_/Q _3133_/X _3135_/X _5620_/Q _3188_/X vssd1 vssd1 vccd1 vccd1 _3189_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4860__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_241_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4093__A _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3966__A1 _5520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4391__A1 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3194__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5629__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2698__D _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5754_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4143__A1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5686_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_264_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3654__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3900__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4731__A _5566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_28_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4382__A1 _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3185__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4382__B2 _3678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput207 _2760_/Y vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_141_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4230_ _4304_/S _4226_/X _4229_/X vssd1 vssd1 vccd1 vccd1 _4230_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4161_ _5446_/Q _4161_/B vssd1 vssd1 vccd1 vccd1 _4161_/X sky130_fd_sc_hd__and2_4
XFILLER_4_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_228_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3112_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3112_/X sky130_fd_sc_hd__clkbuf_1
X_4092_ _4161_/B _4092_/B vssd1 vssd1 vccd1 vccd1 _4092_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3043_ _5765_/A _3010_/X _3041_/Y _3042_/X _3016_/A vssd1 vssd1 vccd1 vccd1 _3043_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4994_ _4994_/A vssd1 vssd1 vccd1 vccd1 _5679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3945_ _5331_/A vssd1 vssd1 vccd1 vccd1 _3945_/X sky130_fd_sc_hd__buf_2
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4641__A _4950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3876_ _3948_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3876_/Y sky130_fd_sc_hd__nand2_1
X_5615_ _5667_/CLK _5615_/D vssd1 vssd1 vccd1 vccd1 _5615_/Q sky130_fd_sc_hd__dfxtp_2
X_2827_ input46/X _5412_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _2829_/A sky130_fd_sc_hd__mux2_2
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3176__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5546_ _5665_/CLK _5546_/D vssd1 vssd1 vccd1 vccd1 _5774_/A sky130_fd_sc_hd__dfxtp_4
X_2758_ _5616_/Q _2652_/X _2756_/X _2757_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2758_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_144_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3581__C1 _3528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5477_ _5722_/CLK _5477_/D vssd1 vssd1 vccd1 vccd1 _5477_/Q sky130_fd_sc_hd__dfxtp_4
X_2689_ _2679_/X _2680_/X _2687_/X _2688_/X vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__o31a_1
X_4428_ _4428_/A _4428_/B vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4220__S1 _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4676__A2 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4088__A _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4359_ _4483_/A _4352_/Y _4355_/X _4358_/X vssd1 vssd1 vccd1 vccd1 _4359_/X sky130_fd_sc_hd__a211o_1
XFILLER_235_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3636__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4833__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3866__S _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5451__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3167__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2914__A2 _2943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3627__B1 _3602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _5620_/Q _3597_/X _3606_/X _3728_/X _3729_/X vssd1 vssd1 vccd1 vccd1 _3730_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4461__A _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3661_ _4301_/S vssd1 vssd1 vccd1 vccd1 _4272_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3158__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5400_ _5492_/CLK _5400_/D vssd1 vssd1 vccd1 vccd1 _5400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3592_ _4045_/A _4419_/A _4408_/A _4050_/A vssd1 vssd1 vccd1 vccd1 _3747_/A sky130_fd_sc_hd__or4_4
X_5331_ _5331_/A _5331_/B _5331_/C vssd1 vssd1 vccd1 vccd1 _5332_/A sky130_fd_sc_hd__and3_1
XANTENNA__5292__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4107__A1 _4108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5262_ _5262_/A vssd1 vssd1 vccd1 vccd1 _5730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3315__C1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4213_ _4213_/A _4213_/B vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__xor2_1
XFILLER_114_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2669__A1 _5625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3866__A0 _5492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5193_ _5772_/A _5193_/B vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__and2_1
XFILLER_205_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4144_ _4466_/A _4059_/B _4469_/B _4469_/C _3613_/X vssd1 vssd1 vccd1 vccd1 _4144_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2855__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4075_ _4066_/Y _4323_/B _4090_/D _4074_/X vssd1 vssd1 vccd1 vccd1 _4194_/A sky130_fd_sc_hd__o31a_1
XFILLER_228_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3026_ _3085_/A _3026_/B _3031_/B vssd1 vssd1 vccd1 vccd1 _3026_/Y sky130_fd_sc_hd__nor3_1
XFILLER_243_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5474__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4977_ _5671_/Q _4972_/B _4976_/Y _4957_/X vssd1 vssd1 vccd1 vccd1 _5671_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4371__A _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4594__A1 _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3928_ _3965_/A _3928_/B vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__or2_1
XFILLER_211_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3859_ _5329_/A _3893_/A _3919_/A _5491_/Q vssd1 vssd1 vccd1 vccd1 _5491_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4346__A1 _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5529_ _5707_/CLK _5529_/D vssd1 vssd1 vccd1 vccd1 _5529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_105_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3857__B1 _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3321__A2 _2928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3609__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4546__A _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4282__B1 _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4821__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4279__A_N _4014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4281__A _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_226_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_269_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5347__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3312__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5497__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4900_ _5638_/Q _4897_/B _4899_/Y _4886_/X vssd1 vssd1 vccd1 vccd1 _5638_/D sky130_fd_sc_hd__o211a_1
XFILLER_280_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2823__A1 _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4831_ _5609_/Q _4822_/B _4830_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5609_/D sky130_fd_sc_hd__o211a_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4903__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4762_ _5682_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__and2_1
XFILLER_193_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_267_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3713_ _5626_/Q _3597_/X _3598_/X _5610_/Q _3712_/X vssd1 vssd1 vccd1 vccd1 _3713_/X
+ sky130_fd_sc_hd__a221o_2
X_4693_ _4697_/A _4970_/A vssd1 vssd1 vccd1 vccd1 _4693_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4328__A1 _3555_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3644_ _5666_/Q _3600_/X _3606_/A _3643_/X vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3238__C _5480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3575_ _5483_/Q _5323_/A _3588_/S vssd1 vssd1 vccd1 vccd1 _4050_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3535__A _4083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5314_ _5749_/Q _5295_/X _5313_/X _4979_/X vssd1 vssd1 vccd1 vccd1 _5749_/D sky130_fd_sc_hd__o211a_1
XFILLER_216_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5245_ _5261_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__and2_1
XANTENNA__3303__A2 _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5176_ _4599_/B _5175_/X _4593_/Y vssd1 vssd1 vccd1 vccd1 _5177_/B sky130_fd_sc_hd__o21ai_2
XFILLER_256_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4127_ _4132_/A _4071_/B _3613_/X _4469_/C _4469_/B vssd1 vssd1 vccd1 vccd1 _4127_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_232_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_300 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_283_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4058_ _4059_/A _4059_/B _4059_/C vssd1 vssd1 vccd1 vccd1 _4441_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3067__A1 _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4803__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3009_ _5355_/Q _5678_/Q vssd1 vssd1 vccd1 vccd1 _3063_/B sky130_fd_sc_hd__nor2_2
XANTENNA__2814__A1 _5685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4319__A1 _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4178__S0 _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4276__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3058__A1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3330__D _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3766__C1 _3843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3230__A1 _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3781__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5046__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2897__C _5362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4730__A1 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3360_ _3003_/B _5363_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3361_/A sky130_fd_sc_hd__mux2_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2741__B1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _5365_/Q _5366_/Q _3290_/Y _3795_/A _5333_/Q vssd1 vssd1 vccd1 vccd1 _5333_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_151_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_257_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5030_ _5696_/Q _5156_/A _5030_/S vssd1 vssd1 vccd1 vccd1 _5031_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3802__B _3802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__D _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3240__D _5476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4914__A _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _5602_/Q _4819_/A vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__or2_1
XFILLER_178_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4549__A1 _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3249__B _5478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3221__A1 _5642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4745_ _5331_/A vssd1 vssd1 vccd1 vccd1 _4745_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5512__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3964__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4676_ _4642_/Y _4674_/X _4675_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _5553_/D sky130_fd_sc_hd__o211a_1
X_3627_ _5664_/Q _3600_/A _3602_/A _5648_/Q vssd1 vssd1 vccd1 vccd1 _3627_/X sky130_fd_sc_hd__a22o_1
XFILLER_227_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3558_ _4428_/A _4372_/B vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__nor2_8
XANTENNA__5662__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3489_ _3489_/A vssd1 vssd1 vccd1 vccd1 _5424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5228_ _5775_/A _5193_/B _5227_/X _5071_/B vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__a22o_1
XFILLER_248_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4808__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4096__A _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5159_ _5712_/Q _5158_/X _5233_/S vssd1 vssd1 vccd1 vccd1 _5160_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4527__C _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4237__B1 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4824__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4543__B _4543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3212__A1 _5560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4960__A1 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3920__C1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3903__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4476__B1 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_235_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3987__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__A1 _3091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5535__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2860_ _5357_/Q _2794_/Y _2823_/Y _2858_/X _3016_/A vssd1 vssd1 vccd1 vccd1 _3343_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3203__A1 _5671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3784__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2791_ _5548_/Q _2791_/B vssd1 vssd1 vccd1 vccd1 _2791_/X sky130_fd_sc_hd__or2_1
XFILLER_178_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4530_ _4585_/A _4525_/X _4528_/X _4529_/X vssd1 vssd1 vccd1 vccd1 _4530_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3754__A2 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4461_ _4600_/A _5051_/B vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__nand2_2
XANTENNA__2701__B _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3085__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3412_ _3412_/A vssd1 vssd1 vccd1 vccd1 _5385_/D sky130_fd_sc_hd__clkbuf_1
X_4392_ _5449_/Q _4043_/A _2904_/X vssd1 vssd1 vccd1 vccd1 _4392_/X sky130_fd_sc_hd__a21o_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _5331_/A _3343_/B _3343_/C vssd1 vssd1 vccd1 vccd1 _3344_/A sky130_fd_sc_hd__and3_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_132 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _5253_/S _3273_/X _3851_/B vssd1 vssd1 vccd1 vccd1 _5678_/D sky130_fd_sc_hd__a21o_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5688_/Q _3755_/Y _5030_/S vssd1 vssd1 vccd1 vccd1 _5014_/A sky130_fd_sc_hd__mux2_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3959__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4363__B _4363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2989_ _2974_/Y _2852_/B _2845_/C _2988_/Y vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3745__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4942__A1 _5656_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4728_ _4646_/X _4724_/Y _4727_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5564_/D sky130_fd_sc_hd__o211a_1
X_4659_ _5550_/Q _4722_/A vssd1 vssd1 vccd1 vccd1 _4659_/X sky130_fd_sc_hd__or2_1
XFILLER_238_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2705__B1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4819__A _4819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5408__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4473__A3 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5558__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3736__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2802__A _5678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4729__A _5565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3121__A0 _5708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3672__B2 _5548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _3965_/A _3961_/B vssd1 vssd1 vccd1 vccd1 _3961_/X sky130_fd_sc_hd__or2_1
X_5700_ _5724_/CLK _5700_/D vssd1 vssd1 vccd1 vccd1 _5700_/Q sky130_fd_sc_hd__dfxtp_1
X_2912_ _2912_/A vssd1 vssd1 vccd1 vccd1 _5452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3892_ _5502_/Q _5317_/A _3905_/S vssd1 vssd1 vccd1 vccd1 _3893_/B sky130_fd_sc_hd__mux2_1
X_5631_ _5667_/CLK _5631_/D vssd1 vssd1 vccd1 vccd1 _5631_/Q sky130_fd_sc_hd__dfxtp_2
X_2843_ input40/X _5434_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2845_/C sky130_fd_sc_hd__mux2_2
XANTENNA__3188__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3727__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4924__A1 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5562_ _5675_/CLK _5562_/D vssd1 vssd1 vccd1 vccd1 _5562_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__2712__A _5557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2774_ _2775_/B _2789_/B _2774_/C _5630_/Q vssd1 vssd1 vccd1 vccd1 _2774_/X sky130_fd_sc_hd__and4b_1
X_4513_ _3935_/A _5015_/A _4626_/S vssd1 vssd1 vccd1 vccd1 _4513_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5493_ _5741_/CLK _5493_/D vssd1 vssd1 vccd1 vccd1 _5493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_343 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4444_ _2936_/X _4418_/A _2919_/X vssd1 vssd1 vccd1 vccd1 _4444_/X sky130_fd_sc_hd__a21o_1
XFILLER_144_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4152__A2 _4150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4375_ _4396_/A _4375_/B vssd1 vssd1 vccd1 vccd1 _4375_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3543__A _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3326_ _2771_/B _5486_/D _3325_/X vssd1 vssd1 vccd1 vccd1 _5345_/D sky130_fd_sc_hd__o21a_2
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5101__A1 _4537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5700__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3257_ _5349_/Q vssd1 vssd1 vccd1 vccd1 _3265_/B sky130_fd_sc_hd__inv_2
XANTENNA__5101__B2 _5100_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5492_/CLK sky130_fd_sc_hd__clkbuf_16
X_3188_ _5668_/Q _3137_/X _3139_/X _5588_/Q vssd1 vssd1 vccd1 vccd1 _3188_/X sky130_fd_sc_hd__a22o_1
XFILLER_226_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_214_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4612__B1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2754__A_N _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3179__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4376__C1 _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4391__A2 _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4143__A2 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5380__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3654__A1 _5630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3273__C_N _3252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input12_A i_mem_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_217_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5159__A1 _5158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_82 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2772__B_N _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4731__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4223__S _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4906__A1 _5641_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2917__B1 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput208 _5307_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_153_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_387 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5723__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4160_ _4160_/A vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__buf_4
X_3111_ _5711_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3112_/A sky130_fd_sc_hd__and2_1
XFILLER_255_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4091_ _4192_/A _4091_/B vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__and2b_1
XFILLER_255_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5095__B1 _5051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3042_ _2840_/D _3027_/X _3343_/C vssd1 vssd1 vccd1 vccd1 _3042_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3645__A1 _5554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2707__A _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2853__C1 _2829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4993_ _4690_/X _3790_/X _5720_/D vssd1 vssd1 vccd1 vccd1 _4994_/A sky130_fd_sc_hd__mux2_1
XFILLER_210_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3944_ _3948_/B _3942_/X _3943_/Y _3965_/A vssd1 vssd1 vccd1 vccd1 _3944_/X sky130_fd_sc_hd__a211o_1
XFILLER_211_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3875_ _5495_/Q _3874_/B _3874_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _5495_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5229__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3538__A _5470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5614_ _5653_/CLK _5614_/D vssd1 vssd1 vccd1 vccd1 _5614_/Q sky130_fd_sc_hd__dfxtp_1
X_2826_ _2826_/A _2835_/A vssd1 vssd1 vccd1 vccd1 _2830_/A sky130_fd_sc_hd__or2b_1
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5545_ _5665_/CLK _5545_/D vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2757_ _2789_/B _2782_/C _5648_/Q _2757_/D vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__and4b_1
XANTENNA__3972__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3581__B1 _2738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5476_ _5722_/CLK _5476_/D vssd1 vssd1 vccd1 vccd1 _5476_/Q sky130_fd_sc_hd__dfxtp_4
X_2688_ _5559_/Q _2791_/B vssd1 vssd1 vccd1 vccd1 _2688_/X sky130_fd_sc_hd__or2_1
X_4427_ _4469_/D _4146_/B _4426_/X vssd1 vssd1 vccd1 vccd1 _4427_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_132_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4530__C1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4358_ _5445_/Q _4031_/X _4348_/A _5449_/Q _4357_/X vssd1 vssd1 vccd1 vccd1 _4358_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2687__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input4_A dbg_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3309_ _3309_/A _3322_/A _3309_/C vssd1 vssd1 vccd1 vccd1 _3310_/B sky130_fd_sc_hd__or3_2
XFILLER_98_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4289_ _4537_/B _4522_/B _4289_/C _4289_/D vssd1 vssd1 vccd1 vccd1 _4362_/C sky130_fd_sc_hd__or4_1
XFILLER_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3636__A1 _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3636__B2 _5651_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4597__C1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4832__A _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5746__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3572__B1 _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2914__A3 _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3324__B1 _3323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5077__A0 _5060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3627__A1 _5664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3627__B2 _5648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4461__B _5051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _5551_/Q _3596_/A _3657_/X _3659_/X vssd1 vssd1 vccd1 vccd1 _4024_/B sky130_fd_sc_hd__o22a_4
XANTENNA__5001__A0 _5683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3591_ _4128_/A vssd1 vssd1 vccd1 vccd1 _4469_/B sky130_fd_sc_hd__buf_2
XFILLER_186_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5329_/Y _4690_/X _5720_/Q vssd1 vssd1 vccd1 vccd1 _5331_/C sky130_fd_sc_hd__mux2_1
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4760__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5261_ _5261_/A _5261_/B vssd1 vssd1 vccd1 vccd1 _5262_/A sky130_fd_sc_hd__and2_1
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5304__A1 _2768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4212_ _3615_/X _4468_/B _4468_/A vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3315__B1 _3310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5192_ _5192_/A _5187_/B vssd1 vssd1 vccd1 vccd1 _5198_/B sky130_fd_sc_hd__or2b_1
XANTENNA__3866__A1 _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2669__A2 _2652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4143_ _4466_/A _4415_/A _4469_/B _4469_/C _3613_/X vssd1 vssd1 vccd1 vccd1 _4143_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__4917__A _5645_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4074_ _4072_/Y _4070_/A _4073_/A vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3618__A1 _5480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3540__B _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3025_ _5392_/Q _5391_/Q _5390_/Q vssd1 vssd1 vccd1 vccd1 _3031_/B sky130_fd_sc_hd__and3_1
XFILLER_221_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5619__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3967__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5756_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_251_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4976_ _4976_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_251_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4594__A2 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3927_ _3926_/X _5067_/B _3984_/S vssd1 vssd1 vccd1 vccd1 _3928_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3268__A _5471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3858_ _5723_/Q _3893_/A _3919_/A _5490_/Q vssd1 vssd1 vccd1 vccd1 _5490_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5598_/CLK sky130_fd_sc_hd__clkbuf_16
X_2809_ _5341_/Q vssd1 vssd1 vccd1 vccd1 _3601_/C sky130_fd_sc_hd__buf_4
X_3789_ _3789_/A vssd1 vssd1 vccd1 vccd1 _5463_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2900__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5528_ _5528_/CLK _5528_/D vssd1 vssd1 vccd1 vccd1 _5528_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_59_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5459_ _5743_/CLK _5459_/D vssd1 vssd1 vccd1 vccd1 _5459_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_132_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_219_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5059__B1 _5460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3609__A1 _5579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3609__B2 _5595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4282__A1 _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__A _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__A0 _4482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_360 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3906__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4742__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3117__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_257_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4737__A _5569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2823__A2 _3346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4830_ _4981_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4830_/Y sky130_fd_sc_hd__nand2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4761_ _5682_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4761_/Y sky130_fd_sc_hd__nand2_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3784__A0 _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3712_ _5674_/Q _3600_/X _3602_/X _5658_/Q vssd1 vssd1 vccd1 vccd1 _3712_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4692_ input21/X _4689_/X _4690_/X _4691_/Y vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_267_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3643_ _5634_/Q _3605_/A _3607_/A _5570_/Q vssd1 vssd1 vccd1 vccd1 _3643_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3238__D _5483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2720__A _5556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3574_ _5485_/Q _2650_/Y _3588_/S vssd1 vssd1 vccd1 vccd1 _4408_/A sky130_fd_sc_hd__mux2_2
XFILLER_161_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5313_ _5313_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__or2_1
XFILLER_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5244_ _5725_/Q _4527_/C _5253_/S vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4647__A _5680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5175_ _5770_/A _5193_/B _5174_/Y _5196_/A vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5242__S _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3551__A _5474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _5454_/Q _4161_/B _3613_/X _4128_/B _4128_/A vssd1 vssd1 vccd1 vccd1 _4394_/A
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5441__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4057_ _5453_/Q vssd1 vssd1 vccd1 vccd1 _4171_/A sky130_fd_sc_hd__clkinv_2
XFILLER_45_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3008_ _5760_/A vssd1 vssd1 vccd1 vccd1 _4527_/C sky130_fd_sc_hd__buf_4
XFILLER_271_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5065__A2_N _5062_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2814__A2 _5686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5591__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _5663_/Q _4985_/B vssd1 vssd1 vccd1 vccd1 _4959_/X sky130_fd_sc_hd__or2_1
XFILLER_177_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2750__A1 _2744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4178__S1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4991__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3270__A_N _5470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2805__A _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3230__A2 _3346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_224 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4231__S _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4191__B1 _4192_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4730__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2741__A1 _5586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5464__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3290_ _3300_/B vssd1 vssd1 vccd1 vccd1 _3290_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4467__A _4467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4246__A1 _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4813_ _4674_/X _4799_/Y _4812_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _5601_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4549__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3757__A0 _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _4970_/A _4747_/B vssd1 vssd1 vccd1 vccd1 _4744_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3221__A2 _3143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_i_clk_A clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4675_ _5553_/Q _4687_/A vssd1 vssd1 vccd1 vccd1 _4675_/X sky130_fd_sc_hd__or2_1
XANTENNA__3546__A _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3626_ _3622_/X _3623_/X _3625_/X _3596_/A _5553_/Q vssd1 vssd1 vccd1 vccd1 _4232_/B
+ sky130_fd_sc_hd__o32a_4
XANTENNA__4706__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3557_ _4474_/A _4124_/A _4067_/A _3556_/X vssd1 vssd1 vccd1 vccd1 _4372_/B sky130_fd_sc_hd__a211o_4
XANTENNA__3980__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5761__A _5761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3488_ _5424_/Q input29/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3489_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5227_ _5756_/Q _3840_/X _5226_/X vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3281__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _5157_/X _5313_/A _5179_/S vssd1 vssd1 vccd1 vccd1 _5158_/X sky130_fd_sc_hd__mux2_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _4370_/B _4109_/B vssd1 vssd1 vccd1 vccd1 _4386_/C sky130_fd_sc_hd__or2_1
XFILLER_256_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5089_ _5200_/B _5087_/Y _5088_/X _5179_/S vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__a31o_1
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4824__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2874__C_N _5362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5337__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5201__A3 _5225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4840__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3212__A2 _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4960__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4173__A0 _4149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_284_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input42_A i_req_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4476__A1 _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output129_A _5689_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2660__A_N _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4226__S _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4936__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2790_ _5612_/Q _2652_/X _2788_/X _2789_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2790_/X
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__4400__A1 _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3203__A2 _3137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_20_i_clk_A clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4460_ _5528_/Q _4458_/A _4459_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5528_/D sky130_fd_sc_hd__o211a_1
XFILLER_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3411_ _2967_/A _5385_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3412_/A sky130_fd_sc_hd__mux2_1
X_4391_ _2936_/X _4363_/A _4363_/B _4390_/X vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__a31o_1
XFILLER_264_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3342_ _5263_/A vssd1 vssd1 vccd1 vccd1 _5331_/A sky130_fd_sc_hd__buf_6
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3273_ _3273_/A _3273_/B _3252_/B vssd1 vssd1 vccd1 vccd1 _3273_/X sky130_fd_sc_hd__or3b_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A vssd1 vssd1 vccd1 vccd1 _5687_/D sky130_fd_sc_hd__clkbuf_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__C1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4925__A _5649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3975__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2988_ _5398_/Q vssd1 vssd1 vccd1 vccd1 _2988_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4727_ _5564_/Q _4759_/B vssd1 vssd1 vccd1 vccd1 _4727_/X sky130_fd_sc_hd__or2_1
XFILLER_147_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4942__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4658_ _4658_/A vssd1 vssd1 vccd1 vccd1 _4658_/X sky130_fd_sc_hd__buf_4
X_3609_ _5579_/Q _3607_/X _3608_/X _5595_/Q vssd1 vssd1 vccd1 vccd1 _3609_/X sky130_fd_sc_hd__a22o_1
X_4589_ _4590_/B _4581_/B _4585_/X _4588_/X _3919_/X vssd1 vssd1 vccd1 vccd1 _5541_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2705__A1 _5573_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3902__A0 _5505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2705__B2 _5605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4630__A1 _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4918__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4570__A _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3197__A1 _5557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2802__B _3851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2944__A1 _2938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4729__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4449__A1 _4424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3125__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4515__B1_N _4514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5502__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4745__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3960_ _3959_/X _5311_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3961_/B sky130_fd_sc_hd__mux2_1
X_2911_ _2904_/X _2910_/X _3337_/B vssd1 vssd1 vccd1 vccd1 _2912_/A sky130_fd_sc_hd__mux2_1
X_3891_ _3891_/A vssd1 vssd1 vccd1 vccd1 _5501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_250_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5630_ _5653_/CLK _5630_/D vssd1 vssd1 vccd1 vccd1 _5630_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4909__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2842_ input34/X _5429_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2845_/B sky130_fd_sc_hd__mux2_2
XANTENNA__3188__A1 _5668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3188__B2 _5588_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2773_ _2774_/C _2789_/B _2789_/C _5582_/Q vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__and4bb_1
XFILLER_191_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4924__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5561_ _5675_/CLK _5561_/D vssd1 vssd1 vccd1 vccd1 _5561_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__2712__B _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2935__A1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4512_ _4550_/S vssd1 vssd1 vccd1 vccd1 _4626_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_156_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5492_ _5492_/CLK _5492_/D vssd1 vssd1 vccd1 vccd1 _5492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4443_ _4422_/B _4443_/B _4483_/A vssd1 vssd1 vccd1 vccd1 _4443_/X sky130_fd_sc_hd__and3b_1
XFILLER_208_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4374_ _4140_/Y _4141_/Y _4177_/Y _4373_/Y _4272_/S _4146_/A vssd1 vssd1 vccd1 vccd1
+ _4375_/B sky130_fd_sc_hd__mux4_1
XFILLER_208_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4152__A3 _4151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3543__B _4307_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3360__A1 _5363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3325_ _5369_/Q _3335_/B _3335_/C _5372_/Q _3293_/A vssd1 vssd1 vccd1 vccd1 _3325_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_224_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3256_ _5529_/Q _5350_/Q _5351_/Q vssd1 vssd1 vccd1 vccd1 _3256_/X sky130_fd_sc_hd__or3b_1
XANTENNA__5101__A2 _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_273_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3187_ _5555_/Q _3131_/X _3184_/X _3186_/X vssd1 vssd1 vccd1 vccd1 _3187_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5250__S _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4860__A1 _5621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4299__S0 _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4612__A1 _5198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3179__A1 _5602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3179__B2 _5618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3718__B _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4391__A3 _4363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5525__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4851__A1 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3654__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5675__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2813__A _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4906__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output196_A _5479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2917__A1 _3307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput209 _2743_/Y vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_153_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5316__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output73_A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3110_ _3110_/A vssd1 vssd1 vccd1 vccd1 _3110_/X sky130_fd_sc_hd__clkbuf_1
X_4090_ _4090_/A _4090_/B _4323_/B _4090_/D vssd1 vssd1 vccd1 vccd1 _4194_/B sky130_fd_sc_hd__or4_1
XFILLER_255_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5095__B2 _5531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3041_ _3085_/A _3045_/B _3041_/C vssd1 vssd1 vccd1 vccd1 _3041_/Y sky130_fd_sc_hd__nor3_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3645__A2 _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2853__B1 _2829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4992_ _4992_/A vssd1 vssd1 vccd1 vccd1 _5677_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_223_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ _3943_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _3943_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4704__A1_N input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3874_ _3943_/A _3874_/B vssd1 vssd1 vccd1 vccd1 _3874_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4358__B1 _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5613_ _5653_/CLK _5613_/D vssd1 vssd1 vccd1 vccd1 _5613_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_176_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2825_ input35/X _5411_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2835_/A sky130_fd_sc_hd__mux2_2
XFILLER_176_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5544_ _5665_/CLK _5544_/D vssd1 vssd1 vccd1 vccd1 _5772_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2756_ _2757_/D _2782_/B _2782_/C _5584_/Q vssd1 vssd1 vccd1 vccd1 _2756_/X sky130_fd_sc_hd__and4bb_1
XFILLER_191_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3581__A1 _5554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5548__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2687_ _5623_/Q _2652_/X _2684_/X _2685_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2687_/X
+ sky130_fd_sc_hd__a2111o_2
X_5475_ _5722_/CLK _5475_/D vssd1 vssd1 vccd1 vccd1 _5475_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3554__A _4306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4426_ _4146_/A _4424_/Y _4425_/X _4471_/S _4372_/A vssd1 vssd1 vccd1 vccd1 _4426_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_132_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3333__B2 _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4357_ _5452_/Q _4029_/X _4356_/X vssd1 vssd1 vccd1 vccd1 _4357_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5698__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3308_ _3308_/A _3800_/B _3308_/C _3308_/D vssd1 vssd1 vccd1 vccd1 _3309_/C sky130_fd_sc_hd__or4_1
XFILLER_100_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4288_ _4500_/A _5015_/A vssd1 vssd1 vccd1 vccd1 _4289_/D sky130_fd_sc_hd__nand2_1
XFILLER_140_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3239_ _5478_/Q _3270_/C _3270_/D _5470_/Q vssd1 vssd1 vccd1 vccd1 _5094_/B sky130_fd_sc_hd__and4b_1
XFILLER_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3636__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4833__A1 _5610_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4832__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4349__B1 _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_299 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4364__A3 _4041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3572__B2 _5548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_145_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3324__A1 _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4521__B1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_277_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3627__A2 _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3403__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output111_A _5558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output209_A _2743_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4588__B1 _4529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5404_/CLK sky130_fd_sc_hd__clkbuf_16
X_3590_ _3590_/A _4363_/A _3619_/A _3590_/D vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__nor4_4
XFILLER_173_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5260_ _5730_/Q _5765_/A _5285_/S vssd1 vssd1 vccd1 vccd1 _5261_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4211_ _4173_/X _4180_/B _4471_/S vssd1 vssd1 vccd1 vccd1 _4468_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191_ _5191_/A vssd1 vssd1 vccd1 vccd1 _5715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_268_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4142_ _4140_/Y _4141_/Y _4447_/S vssd1 vssd1 vccd1 vccd1 _4142_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4917__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4073_ _4073_/A _4072_/Y vssd1 vssd1 vccd1 vccd1 _4090_/D sky130_fd_sc_hd__or2b_1
XFILLER_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3618__A2 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3024_ _5391_/Q _5390_/Q _5392_/Q vssd1 vssd1 vccd1 vccd1 _3026_/B sky130_fd_sc_hd__a21oi_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4933__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4975_ _5670_/Q _4972_/B _4974_/Y _4957_/X vssd1 vssd1 vccd1 vccd1 _5670_/D sky130_fd_sc_hd__o211a_1
XFILLER_211_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3926_ _4527_/C _5725_/Q _5329_/A vssd1 vssd1 vccd1 vccd1 _3926_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5370__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3857_ _3853_/Y _3856_/X _4987_/A vssd1 vssd1 vccd1 vccd1 _5489_/D sky130_fd_sc_hd__a21oi_1
XFILLER_50_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3983__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_214 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5764__A _5764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2808_ _2808_/A _2808_/B vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__or2_1
X_3788_ _5463_/Q _3791_/D _3813_/S vssd1 vssd1 vccd1 vccd1 _3789_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5527_ _5741_/CLK _5527_/D vssd1 vssd1 vccd1 vccd1 _5527_/Q sky130_fd_sc_hd__dfxtp_2
X_2739_ _5666_/Q _2774_/C _2789_/B _2789_/C vssd1 vssd1 vccd1 vccd1 _2739_/X sky130_fd_sc_hd__and4_1
XANTENNA__3284__A _3304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5458_ _5716_/CLK _5458_/D vssd1 vssd1 vccd1 vccd1 _5458_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_172_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4409_ _4409_/A vssd1 vssd1 vccd1 vccd1 _4410_/B sky130_fd_sc_hd__inv_2
XFILLER_182_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5389_ _5722_/CLK _5389_/D vssd1 vssd1 vccd1 vccd1 _5389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_262_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3609__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_227_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4282__A2 _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__B _5132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5713__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5298__A1 _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_280_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4753__A _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5222__A1 _5325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5393__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _5579_/Q _4747_/B _4759_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5579_/D sky130_fd_sc_hd__o211a_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3711_ _4118_/B _3710_/X _4231_/S vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3784__A1 _3319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4691_ _5712_/Q vssd1 vssd1 vccd1 vccd1 _4691_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3642_ _5650_/Q _3602_/A _3598_/A _5602_/Q _3641_/X vssd1 vssd1 vccd1 vccd1 _3642_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3573_ _5484_/Q _5325_/A _3588_/S vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__mux2_2
XANTENNA__2720__B _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5312_ _5748_/Q _5295_/X _5311_/X _4979_/X vssd1 vssd1 vccd1 vccd1 _5748_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5243_ _5243_/A vssd1 vssd1 vccd1 vccd1 _5724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5174_ _5751_/Q _3840_/X _5173_/X vssd1 vssd1 vccd1 vccd1 _5174_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4647__B _4950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3004__D_N _2835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _4276_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4300_/S sky130_fd_sc_hd__xnor2_4
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_15_i_clk_A clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4056_ _4056_/A _4322_/A _4055_/X vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__or3b_1
XFILLER_271_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_271_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3007_ _3007_/A vssd1 vssd1 vccd1 vccd1 _5408_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5736__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4663__A _4663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2814__A3 _5687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3224__B1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4958_ _4658_/X _4949_/Y _4956_/X _4957_/X vssd1 vssd1 vccd1 vccd1 _5662_/D sky130_fd_sc_hd__o211a_1
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3909_ _5507_/Q _3874_/B _3908_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _5507_/D sky130_fd_sc_hd__o211a_1
X_4889_ _4674_/X _4874_/Y _4888_/X _4886_/X vssd1 vssd1 vccd1 vccd1 _5633_/D sky130_fd_sc_hd__o211a_1
XFILLER_177_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3726__B _4130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4838__A _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4488__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_215_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4660__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_230_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3215__B1 _3149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3766__A1 _4529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5609__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2741__A2 _2635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5740_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5650_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4246__A2 _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4483__A _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3099__A _5705_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4812_ _5601_/Q _4819_/A vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__or2_1
XFILLER_278_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3206__B1 _3145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_158 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3757__A1 _3755_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4743_ _4743_/A vssd1 vssd1 vccd1 vccd1 _4747_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_159_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4674_ _4674_/A vssd1 vssd1 vccd1 vccd1 _4674_/X sky130_fd_sc_hd__buf_4
XFILLER_174_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3625_ _5633_/Q _3605_/A _3606_/A _3624_/X vssd1 vssd1 vccd1 vccd1 _3625_/X sky130_fd_sc_hd__a211o_1
X_3556_ _4030_/A _3556_/B vssd1 vssd1 vccd1 vccd1 _3556_/X sky130_fd_sc_hd__xor2_2
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4658__A _4658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3487_ _3487_/A vssd1 vssd1 vccd1 vccd1 _5423_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5253__S _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5226_ _5527_/Q _3932_/B _3864_/C _5507_/Q _5053_/X vssd1 vssd1 vccd1 vccd1 _5226_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_229_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5157_ _5200_/B _5153_/Y _5166_/A _5156_/X vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3693__B1 _3572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4108_ _4108_/A _4108_/B _4108_/C vssd1 vssd1 vccd1 vccd1 _4109_/B sky130_fd_sc_hd__and3_1
X_5088_ _5060_/B _5077_/S _5086_/Y _4524_/X vssd1 vssd1 vccd1 vccd1 _5088_/X sky130_fd_sc_hd__a211o_1
XFILLER_56_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_256_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2906__A _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _4096_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _4091_/B sky130_fd_sc_hd__or2_1
XFILLER_112_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3501__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_248 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2641__A _5675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4173__A1 _4150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5218__A1_N _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3306__B_N _2938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_279_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4568__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4476__A2 _4485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A i_req_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3411__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3647__A _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5431__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4149__D1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2701__D _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4164__A1 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3410_ _3410_/A vssd1 vssd1 vccd1 vccd1 _5384_/D sky130_fd_sc_hd__clkbuf_1
X_4390_ _2919_/X _4363_/A _4363_/B _4333_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4390_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3911__A1 _5508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3341_ _5300_/A vssd1 vssd1 vccd1 vccd1 _5263_/A sky130_fd_sc_hd__clkinv_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5581__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _5347_/Q _5465_/Q _3267_/B _3761_/A vssd1 vssd1 vccd1 vccd1 _3273_/B sky130_fd_sc_hd__a31o_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5687_/Q _5333_/Q _5030_/S vssd1 vssd1 vccd1 vccd1 _5012_/A sky130_fd_sc_hd__mux2_1
XFILLER_285_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4925__B _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4624__C1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3978__A1 _5523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4941__A _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5775_ _5775_/A vssd1 vssd1 vccd1 vccd1 _5775_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2987_ _2973_/Y _2852_/A _2852_/B _2974_/Y _2986_/X vssd1 vssd1 vccd1 vccd1 _2987_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5225__C_N _5214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4726_ _4743_/A vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_147_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4657_ _5706_/Q _4656_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4658_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5772__A _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3608_ _3608_/A vssd1 vssd1 vccd1 vccd1 _3608_/X sky130_fd_sc_hd__buf_6
X_4588_ _4532_/X _4586_/Y _4587_/X _4529_/A vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__a31o_1
XFILLER_162_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_250 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2705__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3902__A1 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3539_ _2786_/X _2787_/X _2790_/X _2791_/X _3528_/A vssd1 vssd1 vccd1 vccd1 _3673_/B
+ sky130_fd_sc_hd__o311ai_4
XFILLER_254_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5209_ _5225_/B _5214_/B vssd1 vssd1 vccd1 vccd1 _5209_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_190_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3666__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4863__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5454__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4570__B _5311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5158__S _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3197__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2944__A2 _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4997__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3753__A_N _3750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3657__B1 _3602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_60 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_235_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3409__A0 _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2910_ _2943_/C _3283_/B _2957_/B _3775_/A vssd1 vssd1 vccd1 vccd1 _2910_/X sky130_fd_sc_hd__a22o_1
XFILLER_250_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3890_ _3893_/A _3890_/B vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__and2_1
XFILLER_259_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2841_ input45/X _5439_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2845_/A sky130_fd_sc_hd__mux2_2
XFILLER_231_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3188__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5560_ _5675_/CLK _5560_/D vssd1 vssd1 vccd1 vccd1 _5560_/Q sky130_fd_sc_hd__dfxtp_4
X_2772_ _5614_/Q _2775_/D vssd1 vssd1 vccd1 vccd1 _2772_/X sky130_fd_sc_hd__or2b_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2935__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4511_ _4581_/B vssd1 vssd1 vccd1 vccd1 _4511_/X sky130_fd_sc_hd__clkbuf_4
X_5491_ _5722_/CLK _5491_/D vssd1 vssd1 vccd1 vccd1 _5491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4137__A1 _4127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4442_ _4114_/A _4171_/B _4441_/X _4060_/B _4416_/Y vssd1 vssd1 vccd1 vccd1 _4443_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_171_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4373_ _4373_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2699__A1 _5574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3896__B1 _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4001__A _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _2806_/A _5486_/D _3323_/X vssd1 vssd1 vccd1 vccd1 _5344_/D sky130_fd_sc_hd__o21a_2
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3255_ _5528_/Q _5530_/Q _5351_/Q vssd1 vssd1 vccd1 vccd1 _3255_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4845__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3186_ _5635_/Q _3143_/X _3145_/X _3185_/X vssd1 vssd1 vccd1 vccd1 _3186_/X sky130_fd_sc_hd__a211o_1
XFILLER_273_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4860__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5477__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4299__S1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5767__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4612__A2 _4611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3820__A0 _5477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3179__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4376__A1 _4396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3584__C1 _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4709_ _4722_/A _4978_/A vssd1 vssd1 vccd1 vccd1 _4709_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5689_ _5716_/CLK _5689_/D vssd1 vssd1 vccd1 vccd1 _5689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4846__A _5615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3639__B1 _3606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4300__A1 _4220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4851__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4581__A _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3811__A0 _5473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4367__A1 _4386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2917__A2 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output189_A _5472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3327__C1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3878__A0 _5497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output66_A _5761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4827__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3040_ _5394_/Q _3039_/C _5395_/Q vssd1 vssd1 vccd1 vccd1 _3041_/C sky130_fd_sc_hd__a21oi_1
XFILLER_208_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4991_ _5677_/Q _5724_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _4992_/A sky130_fd_sc_hd__mux2_1
X_3942_ _5763_/A _5728_/Q _5329_/A vssd1 vssd1 vccd1 vccd1 _3942_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2723__B _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3873_ _5494_/Q _3874_/B _3872_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _5494_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4358__A1 _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5612_ _5747_/CLK _5612_/D vssd1 vssd1 vccd1 vccd1 _5612_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4358__B2 _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2824_ input24/X _5410_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _2826_/A sky130_fd_sc_hd__mux2_4
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5543_ _5665_/CLK _5543_/D vssd1 vssd1 vccd1 vccd1 _5771_/A sky130_fd_sc_hd__dfxtp_4
X_2755_ _5568_/Q _2644_/X _2752_/X _2753_/X _2754_/X vssd1 vssd1 vccd1 vccd1 _2755_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3581__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5474_ _5722_/CLK _5474_/D vssd1 vssd1 vccd1 vccd1 _5474_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_219_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2686_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__buf_6
XANTENNA__3554__B _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4425_ _4449_/S _4484_/A _4469_/B _4469_/C vssd1 vssd1 vccd1 vccd1 _4425_/X sky130_fd_sc_hd__and4_1
XFILLER_144_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3333__A2 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4530__A1 _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4356_ _5450_/Q _4067_/A _4232_/B _5446_/Q _4160_/A vssd1 vssd1 vccd1 vccd1 _4356_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_48_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3307_ _3307_/A _3330_/C _3775_/C vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__and3_1
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4287_ _4347_/A _4199_/B _4286_/X vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__4818__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3570__A _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3238_ _5479_/Q _5481_/Q _5480_/Q _5483_/Q vssd1 vssd1 vccd1 vccd1 _3270_/D sky130_fd_sc_hd__nor4_1
XANTENNA__4833__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3169_ _5600_/Q _3133_/X _3135_/X _5616_/Q _3168_/X vssd1 vssd1 vccd1 vccd1 _3169_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4597__A1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2780__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4279__C _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4521__A1 _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3324__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5642__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4809__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4588__A1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5200__A _5200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3260__A1 _5530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3548__C1 _3528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4760__A1 _5579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4189__C _5200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4210_ _4040_/X _4025_/Y _4036_/Y _4322_/A vssd1 vssd1 vccd1 vccd1 _4210_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3315__A2 _3318_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ _5715_/Q _5189_/X _5233_/S vssd1 vssd1 vccd1 vccd1 _5191_/A sky130_fd_sc_hd__mux2_1
X_4141_ _4466_/A _4363_/B _4373_/A vssd1 vssd1 vccd1 vccd1 _4141_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4072_ _4071_/A _4071_/B _4071_/C vssd1 vssd1 vccd1 vccd1 _4072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2718__B _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3023_ _3343_/C _3020_/X _3022_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3023_/X sky130_fd_sc_hd__o211a_1
XFILLER_283_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2734__A _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4974_ _4974_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4974_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5110__A _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3549__B _3549_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3925_ _3990_/A vssd1 vssd1 vccd1 vccd1 _3965_/A sky130_fd_sc_hd__buf_2
XANTENNA__5515__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3856_ _5329_/A _5723_/Q _3856_/C _5489_/Q vssd1 vssd1 vccd1 vccd1 _3856_/X sky130_fd_sc_hd__or4b_1
XANTENNA__3539__C1 _3528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2807_ _5684_/Q _5685_/Q _5686_/Q _5687_/Q _2771_/A _2771_/B vssd1 vssd1 vccd1 vccd1
+ _2808_/B sky130_fd_sc_hd__mux4_1
XFILLER_164_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_11_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3787_ _5462_/Q _3780_/A _3786_/X vssd1 vssd1 vccd1 vccd1 _5462_/D sky130_fd_sc_hd__o21a_1
X_5526_ _5756_/CLK _5526_/D vssd1 vssd1 vccd1 vccd1 _5526_/Q sky130_fd_sc_hd__dfxtp_2
X_2738_ _5618_/Q _2652_/X _2735_/X _2736_/X _2737_/X vssd1 vssd1 vccd1 vccd1 _2738_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_117_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5665__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3284__B _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_270 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5457_ _5743_/CLK _5457_/D vssd1 vssd1 vccd1 vccd1 _5457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2669_ _5625_/Q _2652_/A _2667_/X _2668_/X _2686_/A vssd1 vssd1 vccd1 vccd1 _2669_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_246_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4408_ _4408_/A _4484_/A vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__nor2_1
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5388_ _5722_/CLK _5388_/D vssd1 vssd1 vccd1 vccd1 _5388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4339_ _4087_/A _4089_/A _4339_/S vssd1 vssd1 vccd1 vccd1 _4339_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4396__A _4396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2817__A1 _5352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4742__A1 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_269_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5298__A2 _3843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_336 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4753__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5538__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3747_/A _3747_/B _4000_/B vssd1 vssd1 vccd1 vccd1 _3710_/X sky130_fd_sc_hd__or3_1
X_4690_ _4690_/A vssd1 vssd1 vccd1 vccd1 _4690_/X sky130_fd_sc_hd__buf_4
XANTENNA__5688__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3641_ _5618_/Q _3597_/A _3608_/A _5586_/Q vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__a22o_1
X_3572_ _3561_/X _3564_/X _3569_/X _3596_/A _5548_/Q vssd1 vssd1 vccd1 vccd1 _3572_/X
+ sky130_fd_sc_hd__o32a_2
XANTENNA__2744__B1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5311_ _5311_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__or2_1
XANTENNA__3941__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242_ _5724_/Q _5241_/X _5242_/S vssd1 vssd1 vccd1 vccd1 _5243_/A sky130_fd_sc_hd__mux2_1
X_5173_ _5522_/Q _3932_/B _3864_/C _5502_/Q vssd1 vssd1 vccd1 vccd1 _5173_/X sky130_fd_sc_hd__a22o_1
X_4124_ _4124_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__nor2_4
XFILLER_110_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 dbg_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_283_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4055_ _4403_/A _4055_/B _4059_/C vssd1 vssd1 vccd1 vccd1 _4055_/X sky130_fd_sc_hd__or3_1
XFILLER_256_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_283_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3006_ _5408_/Q _3011_/A _3346_/B vssd1 vssd1 vccd1 vccd1 _3007_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4155__S _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4016__A3 _4014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3224__A1 _5611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4957_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4957_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3224__B2 _5627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5775__A _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3908_ _4635_/B _3908_/B vssd1 vssd1 vccd1 vccd1 _3908_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4888_ _5633_/Q _4894_/A vssd1 vssd1 vccd1 vccd1 _4888_/X sky130_fd_sc_hd__or2_1
XFILLER_137_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2983__B1 _2845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3839_ _3839_/A vssd1 vssd1 vccd1 vccd1 _3840_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3295__A _5365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5509_ _5741_/CLK _5509_/D vssd1 vssd1 vccd1 vccd1 _5509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5015__A _5015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3160__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4854__A _5619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5722_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_262_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3215__A1 _5657_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4412__B1 _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3215__B2 _5577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2821__B _4988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3409__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater217_A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3151__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5360__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4764__A _5580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__A3 _4220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_196 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4651__A0 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_358 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3099__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4811_ _4668_/X _4799_/Y _4810_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _5600_/D sky130_fd_sc_hd__o211a_1
XFILLER_261_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3206__A1 _5639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4742_ _4684_/X _4724_/Y _4741_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5571_/D sky130_fd_sc_hd__o211a_1
XFILLER_159_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4673_ _5709_/Q _4672_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__mux2_1
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3624_ _5569_/Q _3607_/A _3608_/A _5585_/Q vssd1 vssd1 vccd1 vccd1 _3624_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4706__A1 _5559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3555_ _5454_/Q _4124_/B _3555_/C vssd1 vssd1 vccd1 vccd1 _3556_/B sky130_fd_sc_hd__and3_1
XFILLER_127_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4939__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2812__S0 _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3390__A0 _2840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3486_ _5423_/Q input28/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3487_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3562__B _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5225_ _5225_/A _5225_/B _5214_/B vssd1 vssd1 vccd1 vccd1 _5230_/A sky130_fd_sc_hd__or3b_1
XANTENNA__5703__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5156_ _5156_/A _5156_/B vssd1 vssd1 vccd1 vccd1 _5156_/X sky130_fd_sc_hd__and2_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3693__A1 _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_256_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4107_ _4108_/A _4108_/B _4108_/C vssd1 vssd1 vccd1 vccd1 _4370_/B sky130_fd_sc_hd__a21oi_2
XFILLER_256_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ _4524_/X _5086_/Y _5077_/S _5060_/B vssd1 vssd1 vccd1 vccd1 _5087_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_229_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4038_ _4192_/C vssd1 vssd1 vccd1 vccd1 _4038_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_271_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2757__A_N _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3804__A1_N _3775_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2641__B _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4173__A2 _4151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5383__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5122__A1 _5307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput190 _5473_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_239_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3899__S _3905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input28_A i_req_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5189__A1 _5319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4397__C1 _4372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4759__A _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5726__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3663__A _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3340_ _3340_/A vssd1 vssd1 vccd1 vccd1 _5354_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A1 _5708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _5055_/A _5461_/Q _3838_/C _3996_/B _4619_/B vssd1 vssd1 vccd1 vccd1 _3761_/A
+ sky130_fd_sc_hd__a41o_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5233_/S vssd1 vssd1 vccd1 vccd1 _5030_/S sky130_fd_sc_hd__buf_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3675__A1 _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4941__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5774_ _5774_/A vssd1 vssd1 vccd1 vccd1 _5774_/X sky130_fd_sc_hd__clkbuf_1
X_2986_ _2973_/Y _2852_/A _2840_/D _2975_/Y _2985_/X vssd1 vssd1 vccd1 vccd1 _2986_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_166_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4725_ _5681_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4743_/A sky130_fd_sc_hd__and2_2
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4656_ input8/X input15/X _4682_/S vssd1 vssd1 vccd1 vccd1 _4656_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3607_ _3607_/A vssd1 vssd1 vccd1 vccd1 _3607_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_162_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4587_ _4590_/B _4590_/C vssd1 vssd1 vccd1 vccd1 _4587_/X sky130_fd_sc_hd__or2_1
XANTENNA__4669__A _5552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5264__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3538_ _5470_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _3673_/A sky130_fd_sc_hd__nand2_2
XFILLER_115_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_254_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3292__B _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5104__A1 _5516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3469_ _5415_/Q input51/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3470_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3115__A0 _5705_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _4619_/B _5207_/X _4619_/Y vssd1 vssd1 vccd1 vccd1 _5214_/B sky130_fd_sc_hd__o21ai_4
XFILLER_130_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3666__A1 _5613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3666__B2 _5597_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5139_ _5539_/Q _5193_/B _5138_/X _5071_/B vssd1 vssd1 vccd1 vccd1 _5140_/B sky130_fd_sc_hd__a22o_1
XFILLER_229_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4615__B1 _4581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4918__A1 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5741_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2652__A _2652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_343 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5749__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5653_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4579__A _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3354__A0 _2829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3657__A1 _5663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3657__B2 _5647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4082__A1 _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4761__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4909__A1 _5642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2840_ _2840_/A _2840_/B _2840_/C _2840_/D vssd1 vssd1 vccd1 vccd1 _2851_/A sky130_fd_sc_hd__or4_1
XFILLER_148_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2771_ _2771_/A _2771_/B vssd1 vssd1 vccd1 vccd1 _2771_/Y sky130_fd_sc_hd__nor2_2
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4510_ _5347_/Q _5469_/Q _3761_/A _5253_/S vssd1 vssd1 vccd1 vccd1 _4581_/B sky130_fd_sc_hd__o31a_2
XANTENNA__3593__B1 _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5490_ _5722_/CLK _5490_/D vssd1 vssd1 vccd1 vccd1 _5490_/Q sky130_fd_sc_hd__dfxtp_1
X_4441_ _4441_/A _4441_/B vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__or2_1
XFILLER_171_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4372_ _4372_/A _4372_/B vssd1 vssd1 vccd1 vccd1 _4372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2699__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3323_ _5370_/Q _3335_/B _3335_/C _5373_/Q _3293_/A vssd1 vssd1 vccd1 vccd1 _3323_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4001__B _4363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3254_ _5350_/Q vssd1 vssd1 vccd1 vccd1 _3265_/A sky130_fd_sc_hd__inv_2
XFILLER_224_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3185_ _5651_/Q _3147_/X _3149_/X _5571_/Q vssd1 vssd1 vccd1 vccd1 _3185_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_214_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4952__A _5660_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3287__B _3802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5757_ _5757_/CLK _5757_/D vssd1 vssd1 vccd1 vccd1 _5757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2969_ _5401_/Q _2969_/B vssd1 vssd1 vccd1 vccd1 _2969_/X sky130_fd_sc_hd__and2_1
XFILLER_185_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_249_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4708_ input10/X _4689_/X _4690_/X _4707_/Y vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__o2bb2a_4
X_5688_ _5716_/CLK _5688_/D vssd1 vssd1 vccd1 vccd1 _5688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4639_ _5775_/A _4511_/X _3919_/A _4638_/X vssd1 vssd1 vccd1 vccd1 _5547_/D sky130_fd_sc_hd__o211a_1
XFILLER_135_357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3507__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5089__B1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3639__A1 _5635_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4846__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5421__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4862__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4581__B _4581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5571__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4367__A2 _4386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3575__A0 _5483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4772__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2917__A3 _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2783__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3417__S _3419_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3327__B1 _3335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3878__A1 _5307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output59_A _3202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2853__A2 _2852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _5032_/A vssd1 vssd1 vccd1 vccd1 _5720_/D sky130_fd_sc_hd__buf_4
XFILLER_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3941_ _5514_/Q _3923_/X _3940_/X _3848_/X vssd1 vssd1 vccd1 vccd1 _5514_/D sky130_fd_sc_hd__o211a_1
XFILLER_204_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3872_ _4523_/B _3874_/B vssd1 vssd1 vccd1 vccd1 _3872_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2723__C _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2823_ _3768_/S _3346_/B _3458_/C vssd1 vssd1 vccd1 vccd1 _2823_/Y sky130_fd_sc_hd__o21ai_1
X_5611_ _5675_/CLK _5611_/D vssd1 vssd1 vccd1 vccd1 _5611_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_176_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2754_ _2789_/C _2782_/B _2774_/C _5632_/Q vssd1 vssd1 vccd1 vccd1 _2754_/X sky130_fd_sc_hd__and4b_1
X_5542_ _5665_/CLK _5542_/D vssd1 vssd1 vccd1 vccd1 _5770_/A sky130_fd_sc_hd__dfxtp_4
X_5473_ _5743_/CLK _5473_/D vssd1 vssd1 vccd1 vccd1 _5473_/Q sky130_fd_sc_hd__dfxtp_4
X_2685_ _2782_/B _2782_/C _5655_/Q _2757_/D vssd1 vssd1 vccd1 vccd1 _2685_/X sky130_fd_sc_hd__and4b_1
XANTENNA__5108__A _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4424_ _4449_/S _4424_/B vssd1 vssd1 vccd1 vccd1 _4424_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4012__A _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4355_ _4355_/A _4355_/B _4355_/C vssd1 vssd1 vccd1 vccd1 _4355_/X sky130_fd_sc_hd__and3_1
XFILLER_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4947__A _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3851__A _5300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3306_ _3306_/A _2938_/X vssd1 vssd1 vccd1 vccd1 _3322_/A sky130_fd_sc_hd__or2b_1
XANTENNA__5444__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4286_ _4355_/A _4271_/Y _4277_/X _4285_/X vssd1 vssd1 vccd1 vccd1 _4286_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3570__B _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3237_ _5482_/Q _5485_/Q _5484_/Q vssd1 vssd1 vccd1 vccd1 _3270_/C sky130_fd_sc_hd__nor3_1
XANTENNA__3062__S _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3168_ _5664_/Q _3137_/X _3139_/X _5584_/Q vssd1 vssd1 vccd1 vccd1 _3168_/X sky130_fd_sc_hd__a22o_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5594__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3099_ _5705_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3100_/A sky130_fd_sc_hd__and2_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3557__B1 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2930__A _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4754__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2780__A1 _5581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2780__B2 _5661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4857__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4521__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3761__A _3761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4285__A1 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input10_A i_mem_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5200__B _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3761__B_N _3267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2840__A _2840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4760__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5467__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3671__A _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _4466_/A _4379_/C _4373_/A vssd1 vssd1 vccd1 vccd1 _4140_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_205_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2709__B_N _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4071_ _4071_/A _4071_/B _4071_/C vssd1 vssd1 vccd1 vccd1 _4073_/A sky130_fd_sc_hd__nor3_1
XANTENNA__2718__C _5652_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3022_ _4533_/C _3063_/B vssd1 vssd1 vccd1 vccd1 _3022_/X sky130_fd_sc_hd__or2_1
XFILLER_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4973_ _5669_/Q _4972_/B _4972_/Y _4957_/X vssd1 vssd1 vccd1 vccd1 _5669_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4007__A _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4984__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3924_ _5291_/S _3989_/S _3851_/B vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__a21oi_2
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3855_ _3988_/S vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__buf_4
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2806_ _2806_/A vssd1 vssd1 vccd1 vccd1 _2808_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__4736__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3786_ _3775_/A _2946_/A _2943_/C _3293_/A vssd1 vssd1 vccd1 vccd1 _3786_/X sky130_fd_sc_hd__a31o_1
XFILLER_164_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3565__B _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5525_ _5740_/CLK _5525_/D vssd1 vssd1 vccd1 vccd1 _5525_/Q sky130_fd_sc_hd__dfxtp_1
X_2737_ _2775_/D _2789_/B _2789_/C _5602_/Q vssd1 vssd1 vccd1 vccd1 _2737_/X sky130_fd_sc_hd__and4b_1
XANTENNA__2762__A1 _5631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3146__A_N input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2762__B2 _5647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5456_ _5743_/CLK _5456_/D vssd1 vssd1 vccd1 vccd1 _5456_/Q sky130_fd_sc_hd__dfxtp_1
X_2668_ _2733_/A _2747_/B _5657_/Q _2747_/D vssd1 vssd1 vccd1 vccd1 _2668_/X sky130_fd_sc_hd__and4b_1
XFILLER_172_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4407_ _4408_/A _4484_/A vssd1 vssd1 vccd1 vccd1 _4410_/A sky130_fd_sc_hd__nand2_1
XFILLER_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5387_ _5404_/CLK _5387_/D vssd1 vssd1 vccd1 vccd1 _5387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _4240_/S _4239_/B _4239_/A vssd1 vssd1 vccd1 vccd1 _4339_/S sky130_fd_sc_hd__a21o_1
XANTENNA__5192__B_N _5187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input2_A dbg_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4269_ _4269_/A _4269_/B vssd1 vssd1 vccd1 vccd1 _4269_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4267__A1 _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2925__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_264_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4019__A1 _5477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4975__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3756__A _5461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_215 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4742__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4587__A _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_265_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2835__A _2835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4966__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3640_ _3636_/X _3637_/X _3639_/X _3596_/A _5555_/Q vssd1 vssd1 vccd1 vccd1 _4161_/B
+ sky130_fd_sc_hd__o32a_4
XFILLER_146_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3571_ _3571_/A vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__buf_6
XANTENNA__2744__A1 _5569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2744__B2 _5601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5310_ _2743_/Y _5319_/B _5309_/X _4979_/X vssd1 vssd1 vccd1 vccd1 _5747_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4497__A _4537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5241_ _5241_/A _5241_/B _5241_/C _5241_/D vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__or4_1
XFILLER_114_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5172_ _5154_/A _5154_/B _5155_/A _5166_/B _5155_/B vssd1 vssd1 vccd1 vccd1 _5182_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4123_ _4372_/A vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__buf_2
XFILLER_268_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4249__A1 _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4054_ _4350_/A vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__clkinv_4
Xinput2 dbg_in[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
XFILLER_256_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_283_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3005_ _2996_/X _3002_/X _3004_/X vssd1 vssd1 vccd1 vccd1 _3011_/A sky130_fd_sc_hd__a21oi_2
XFILLER_283_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2680__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _5662_/Q _4985_/B vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__or2_1
XANTENNA__3224__A2 _3133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5632__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _5506_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4887_ _4668_/X _4874_/Y _4885_/X _4886_/X vssd1 vssd1 vccd1 vccd1 _5632_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5267__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3576__A _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3838_ _5055_/A _5094_/B _3838_/C vssd1 vssd1 vccd1 vccd1 _3839_/A sky130_fd_sc_hd__and3_1
X_3769_ _5456_/Q _3768_/X _5406_/D vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__mux2_1
XFILLER_192_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5508_ _5741_/CLK _5508_/D vssd1 vssd1 vccd1 vccd1 _5508_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5439_ _5722_/CLK _5439_/D vssd1 vssd1 vccd1 vccd1 _5439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4488__A1 _5531_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3515__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3160__A1 _5646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3160__B2 _5566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4854__B _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_215_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4660__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4870__A _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4948__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3215__A2 _3147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4176__B1 _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2726__A1 _5619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3425__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3151__A1 _5628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5505__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4764__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4651__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5655__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2662__B1 _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4810_ _5600_/Q _4819_/A vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__or2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3206__A2 _3143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_221_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _5571_/Q _4743_/A vssd1 vssd1 vccd1 vccd1 _4741_/X sky130_fd_sc_hd__or2_1
XANTENNA__3396__A _3419_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4672_ input11/X input18/X _4682_/S vssd1 vssd1 vccd1 vccd1 _4672_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3623_ _5617_/Q _3597_/A _3598_/A _5601_/Q vssd1 vssd1 vccd1 vccd1 _3623_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3554_ _4306_/A _4326_/A vssd1 vssd1 vccd1 vccd1 _3555_/C sky130_fd_sc_hd__nor2_2
XANTENNA__4939__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2812__S1 _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3843__B _3843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3485_ _3485_/A vssd1 vssd1 vccd1 vccd1 _5422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4020__A _4034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5224_ _5224_/A vssd1 vssd1 vccd1 vccd1 _5718_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3562__C _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5155_ _5155_/A _5155_/B _5154_/Y vssd1 vssd1 vccd1 vccd1 _5166_/A sky130_fd_sc_hd__or3b_1
XANTENNA__3693__A2 _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4106_ _4130_/B vssd1 vssd1 vccd1 vccd1 _4108_/B sky130_fd_sc_hd__inv_2
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5086_ _5081_/Y _5085_/X _5459_/Q vssd1 vssd1 vccd1 vccd1 _5086_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _4037_/A _4008_/X vssd1 vssd1 vccd1 vccd1 _4192_/C sky130_fd_sc_hd__nor2b_2
XFILLER_244_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_271_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2653__B1 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4690__A _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4939_ _4976_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_212_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2956__A1 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2641__C _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3905__A0 _5506_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3753__B _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5528__CLK _5528_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput180 _3435_/S vssd1 vssd1 vccd1 vccd1 o_req_ppl_submit sky130_fd_sc_hd__buf_2
Xoutput191 _5474_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[4] sky130_fd_sc_hd__buf_2
XFILLER_153_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5678__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2_0_i_clk clkbuf_2_3_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_i_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_262_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_247_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2701__A_N _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4936__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4105__A _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4149__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4759__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output89_A _3177_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _5470_/Q _5478_/Q _3270_/C _3270_/D vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__and4bb_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A2 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4775__A _5585_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3675__A2 _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4624__A1 _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_392 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4388__B1 _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5773_ _5773_/A vssd1 vssd1 vccd1 vccd1 _5773_/X sky130_fd_sc_hd__clkbuf_1
X_2985_ _2976_/Y _2840_/B _2840_/D _2975_/Y _2984_/X vssd1 vssd1 vccd1 vccd1 _2985_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4015__A _4306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4724_ _5681_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4724_/Y sky130_fd_sc_hd__nand2_4
XFILLER_238_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4655_ _4642_/Y _4653_/X _4654_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5549_/D sky130_fd_sc_hd__o211a_1
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3854__A _3854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3606_ _3606_/A vssd1 vssd1 vccd1 vccd1 _3606_/X sky130_fd_sc_hd__buf_4
XFILLER_162_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5441_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_238_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4586_ _4590_/B _4590_/C vssd1 vssd1 vccd1 vccd1 _4586_/Y sky130_fd_sc_hd__nand2_1
X_3537_ _3532_/X _3935_/A _3536_/Y vssd1 vssd1 vccd1 vccd1 _4229_/A sky130_fd_sc_hd__o21ai_4
XFILLER_103_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3292__C _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3468_ _3468_/A vssd1 vssd1 vccd1 vccd1 _5414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5207_ _5773_/A _5193_/B _5206_/Y _5196_/A vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4685__A _5555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4863__A1 _5622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3666__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3399_ _2840_/D _5379_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3400_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5138_ _5748_/Q _3840_/X _5137_/X vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2724__A_N _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_270_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5069_ _5704_/Q _5068_/Y _5135_/S vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__mux2_1
XFILLER_244_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4918__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3587__D1 _4006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3051__B1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5328__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5350__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3354__A1 _5360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4551__A0 _5517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input40_A i_req_data[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3657__A2 _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output127_A _5508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_250_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3939__A _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_250 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4909__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3042__B1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2770_ _5566_/Q _2644_/X _2664_/X _5598_/Q _2769_/X vssd1 vssd1 vccd1 vccd1 _2770_/X
+ sky130_fd_sc_hd__a221o_2
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3593__A1 _4306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4440_/A _4440_/B vssd1 vssd1 vccd1 vccd1 _4440_/X sky130_fd_sc_hd__or2_1
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4371_ _4483_/A _4371_/B _4371_/C vssd1 vssd1 vccd1 vccd1 _4384_/B sky130_fd_sc_hd__and3_1
XFILLER_171_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3896__A2 _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3322_ _3322_/A _3322_/B _3321_/X vssd1 vssd1 vccd1 vccd1 _3335_/C sky130_fd_sc_hd__or3b_4
XFILLER_112_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2747__A_N _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3253_ _5291_/S vssd1 vssd1 vccd1 vccd1 _5253_/S sky130_fd_sc_hd__buf_4
XANTENNA__4845__A1 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3184_ _5603_/Q _3133_/X _3135_/X _5619_/Q _3183_/X vssd1 vssd1 vccd1 vccd1 _3184_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_224_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2737__B _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4952__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_356 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5270__A1 _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2753__A _5664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3568__B _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5486__D _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5022__A1 _4543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5373__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5756_ _5756_/CLK _5756_/D vssd1 vssd1 vccd1 vccd1 _5756_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3033__B1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2968_ _5400_/Q _2966_/Y _2969_/B _5401_/Q vssd1 vssd1 vccd1 vccd1 _2968_/X sky130_fd_sc_hd__o22a_1
X_4707_ _5716_/Q vssd1 vssd1 vccd1 vccd1 _4707_/Y sky130_fd_sc_hd__inv_2
X_5687_ _5707_/CLK _5687_/D vssd1 vssd1 vccd1 vccd1 _5687_/Q sky130_fd_sc_hd__dfxtp_2
X_2899_ _2899_/A vssd1 vssd1 vccd1 vccd1 _3795_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4638_ _4634_/Y _4637_/X _4529_/X vssd1 vssd1 vccd1 vccd1 _4638_/X sky130_fd_sc_hd__a21o_1
XFILLER_265_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3336__A1 _5352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4569_ _5519_/Q _4599_/B vssd1 vssd1 vccd1 vccd1 _5154_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5089__A1 _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2928__A _2928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3639__A2 _3605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3523__S _3523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2647__B _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_217_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5716__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3759__A _5512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3272__B1 _3761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5013__A1 _3755_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3575__A1 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4827__A1 _5607_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3433__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3940_ _3948_/B _3938_/X _3939_/Y _3965_/A vssd1 vssd1 vccd1 vccd1 _3940_/X sky130_fd_sc_hd__a211o_1
XFILLER_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4460__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3871_ _5493_/Q _3874_/B _3870_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _5493_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2723__D _5635_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5610_ _5674_/CLK _5610_/D vssd1 vssd1 vccd1 vccd1 _5610_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2638__B_N _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2822_ _5457_/Q _3228_/A vssd1 vssd1 vccd1 vccd1 _3458_/C sky130_fd_sc_hd__nor2_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5541_ _5665_/CLK _5541_/D vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__dfxtp_2
X_2753_ _5664_/Q _2757_/D _2782_/B _2782_/C vssd1 vssd1 vccd1 vccd1 _2753_/X sky130_fd_sc_hd__and4_1
X_5472_ _5743_/CLK _5472_/D vssd1 vssd1 vccd1 vccd1 _5472_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2684_ _2757_/D _2782_/B _2782_/C _5591_/Q vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__and4bb_1
X_4423_ _4466_/A _4418_/A _4373_/A vssd1 vssd1 vccd1 vccd1 _4424_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__5108__B _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2788__B_N _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4012__B _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4354_ _3617_/A _4203_/X _4276_/B _3555_/C vssd1 vssd1 vccd1 vccd1 _4355_/C sky130_fd_sc_hd__a22oi_1
XFILLER_98_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4947__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3851__B _3851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3305_ _3330_/C _2943_/C _3775_/C _3800_/D vssd1 vssd1 vccd1 vccd1 _3306_/A sky130_fd_sc_hd__a31o_1
XFILLER_235_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4285_ _2936_/X _4012_/X _4279_/X _4284_/X vssd1 vssd1 vccd1 vccd1 _4285_/X sky130_fd_sc_hd__a211o_1
XFILLER_98_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4818__A1 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3570__C _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3236_ _4599_/B vssd1 vssd1 vccd1 vccd1 _4619_/B sky130_fd_sc_hd__buf_4
XFILLER_239_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5739__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4963__A _5665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3167_ _5551_/Q _3131_/X _3164_/X _3166_/X vssd1 vssd1 vccd1 vccd1 _3167_/X sky130_fd_sc_hd__o22a_2
XFILLER_251_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5654_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3098_ _3098_/A vssd1 vssd1 vccd1 vccd1 _3098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_214_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5739_ _5740_/CLK _5739_/D vssd1 vssd1 vccd1 vccd1 _5739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_276_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4506__B1 _4289_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2780__A2 _2635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4857__B _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4809__A1 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3568__A_N _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3796__A1 _5466_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4993__A0 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__B2 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3548__A1 _2744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output194_A _5477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2840__B _2840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5209__A _5225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output71_A _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4070_ _4070_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _4323_/B sky130_fd_sc_hd__nand2_1
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2718__D _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3021_ _5761_/A vssd1 vssd1 vccd1 vccd1 _4533_/C sky130_fd_sc_hd__buf_4
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4681__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_236_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_251_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4972_ _4972_/A _4972_/B vssd1 vssd1 vccd1 vccd1 _4972_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3787__A1 _5462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3923_ _3923_/A vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__buf_2
XANTENNA__4007__B _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3854_ _3854_/A vssd1 vssd1 vccd1 vccd1 _3988_/S sky130_fd_sc_hd__buf_4
X_2805_ _2806_/A _2805_/B vssd1 vssd1 vccd1 vccd1 _2805_/X sky130_fd_sc_hd__or2_1
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _5461_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4023__A _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5524_ _5756_/CLK _5524_/D vssd1 vssd1 vccd1 vccd1 _5524_/Q sky130_fd_sc_hd__dfxtp_1
X_2736_ _2774_/C _2789_/C _2789_/B _5570_/Q vssd1 vssd1 vccd1 vccd1 _2736_/X sky130_fd_sc_hd__and4bb_1
XFILLER_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5411__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2762__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5455_ _5692_/CLK _5455_/D vssd1 vssd1 vccd1 vccd1 _5455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2667_ _2747_/D _2733_/A _2747_/B _5593_/Q vssd1 vssd1 vccd1 vccd1 _2667_/X sky130_fd_sc_hd__and4bb_1
XFILLER_117_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4406_ _4055_/B _4403_/X _4440_/A _4052_/A vssd1 vssd1 vccd1 vccd1 _4406_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5386_ _5404_/CLK _5386_/D vssd1 vssd1 vccd1 vccd1 _5386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _4348_/C _4337_/B vssd1 vssd1 vccd1 vccd1 _4337_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5561__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4268_ _4454_/A _4265_/X _4267_/X _4454_/D vssd1 vssd1 vccd1 vccd1 _4269_/B sky130_fd_sc_hd__a211o_1
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3219_ _5610_/Q _3133_/A _3135_/A _5626_/Q _3218_/X vssd1 vssd1 vccd1 vccd1 _3219_/X
+ sky130_fd_sc_hd__a221o_1
X_4199_ _4468_/A _4199_/B vssd1 vssd1 vccd1 vccd1 _4199_/Y sky130_fd_sc_hd__nor2_1
XFILLER_227_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2925__B _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4019__A2 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5216__A1 _5526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5216__B2 _5506_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3860__A_N _5473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2660__B _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3950__A1 _5516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4868__A _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3772__A _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3711__S _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2835__B _2835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5207__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4108__A _4108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3218__B1 _3139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output207_A _2760_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3012__A _5355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5434__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3570_ _3601_/C _3599_/B _3601_/B vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__or3_1
XANTENNA__2997__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2744__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3941__A1 _5514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5584__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3682__A _3683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5143__A0 _4496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5240_/A vssd1 vssd1 vccd1 vccd1 _5723_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4497__B _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5171_ _5171_/A vssd1 vssd1 vccd1 vccd1 _5713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_216_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4326_/A _4122_/B vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__xor2_4
XANTENNA__2826__B_N _2835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4053_ _4403_/A _4055_/B _4059_/C vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__o21a_1
Xinput3 dbg_in[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__3457__B1 _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3004_ _5354_/Q _3004_/B _3004_/C _2835_/A vssd1 vssd1 vccd1 vccd1 _3004_/X sky130_fd_sc_hd__or4b_2
XFILLER_209_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4018__A _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3209__B1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2680__A1 _5639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2680__B2 _5671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4955_ _4653_/X _4949_/Y _4954_/X _4933_/X vssd1 vssd1 vccd1 vccd1 _5661_/D sky130_fd_sc_hd__o211a_1
XFILLER_196_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3906_ _5261_/A _3906_/B vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__and2_1
X_4886_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__buf_4
XANTENNA__3576__B _4408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2983__A2 _2850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3837_ _3837_/A vssd1 vssd1 vccd1 vccd1 _5485_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4185__A1 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4185__B2 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3768_ _5408_/D _5407_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3768_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5507_ _5741_/CLK _5507_/D vssd1 vssd1 vccd1 vccd1 _5507_/Q sky130_fd_sc_hd__dfxtp_1
X_2719_ _5620_/Q _2652_/X _2717_/X _2718_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2719_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3592__A _4045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3699_ _5577_/Q _3607_/X _3608_/X _5593_/Q vssd1 vssd1 vccd1 vccd1 _3699_/X sky130_fd_sc_hd__a22o_1
XFILLER_279_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5438_ _5441_/CLK _5438_/D vssd1 vssd1 vccd1 vccd1 _5438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4488__A2 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5369_ _5757_/CLK _5369_/D vssd1 vssd1 vccd1 vccd1 _5369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4893__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3160__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4620__B1_N _4619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4627__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2936__A _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_274_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4660__A2 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5457__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4870__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__A _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4176__A1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2726__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4884__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3151__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3441__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4636__C1 _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2662__A1 _2653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2662__B2 _5562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3677__A _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4272__S _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4679_/X _4724_/Y _4739_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5570_/D sky130_fd_sc_hd__o211a_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5182__B_N _5177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4671_ _4642_/Y _4668_/X _4669_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _5552_/D sky130_fd_sc_hd__o211a_1
XFILLER_186_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3622_ _5665_/Q _3600_/A _3602_/X _5649_/Q vssd1 vssd1 vccd1 vccd1 _3622_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3553_ _3532_/X _4523_/B _3533_/Y vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__o21ai_4
XFILLER_227_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3484_ _5422_/Q input27/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3485_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5223_ _5718_/Q _5222_/X _5233_/S vssd1 vssd1 vccd1 vccd1 _5224_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4020__B _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5154_ _5154_/A _5154_/B vssd1 vssd1 vccd1 vccd1 _5154_/Y sky130_fd_sc_hd__nand2_1
XFILLER_243_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ _4363_/A _4105_/B _4377_/A vssd1 vssd1 vccd1 vccd1 _4368_/B sky130_fd_sc_hd__and3_1
XANTENNA__4447__S _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5085_ _5082_/Y _5083_/Y _5084_/Y _5460_/Q vssd1 vssd1 vccd1 vccd1 _5085_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5132__A _5132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4036_ _4036_/A _4036_/B vssd1 vssd1 vccd1 vccd1 _4036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_271_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2653__A1 _5594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2653__B2 _5626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4938_ _5654_/Q _4935_/B _4937_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5654_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2956__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4869_ _5625_/Q _4859_/B _4868_/Y _4862_/X vssd1 vssd1 vccd1 vccd1 _5625_/D sky130_fd_sc_hd__o211a_1
XFILLER_177_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2641__D _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3905__A1 _5325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5307__A _5307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3753__C _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput170 _3091_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[15] sky130_fd_sc_hd__buf_2
Xoutput181 _5470_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[0] sky130_fd_sc_hd__buf_2
Xoutput192 _5475_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[5] sky130_fd_sc_hd__buf_2
XANTENNA__4330__A1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4330__B2 _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_247_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4881__A _5630_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3841__B1 _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_270_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4105__B _4105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4149__A1 _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4121__A _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4321__A1 _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4791__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3832__A0 _5483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5772_ _5772_/A vssd1 vssd1 vccd1 vccd1 _5772_/X sky130_fd_sc_hd__clkbuf_1
X_2984_ _2977_/Y _2845_/B _2840_/B _2976_/Y _2983_/X vssd1 vssd1 vccd1 vccd1 _2984_/X
+ sky130_fd_sc_hd__o221a_1
X_4723_ _5563_/Q _4697_/A _4722_/Y _4718_/X vssd1 vssd1 vccd1 vccd1 _5563_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4015__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4654_ _5549_/Q _4722_/A vssd1 vssd1 vccd1 vccd1 _4654_/X sky130_fd_sc_hd__or2_1
XFILLER_238_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3605_ _3605_/A vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__clkbuf_8
Xinput50 i_req_data[4] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
X_4585_ _4585_/A _4585_/B vssd1 vssd1 vccd1 vccd1 _4585_/X sky130_fd_sc_hd__and2_1
XANTENNA__3899__A0 _5504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4031__A _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3536_ _5471_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _3536_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3292__D _3292_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3467_ _5414_/Q input50/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3468_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3870__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4312__A1 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5206_ _5754_/Q _3840_/X _5205_/X vssd1 vssd1 vccd1 vccd1 _5206_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3398_ _3398_/A vssd1 vssd1 vccd1 vccd1 _5378_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4863__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5137_ _5519_/Q _3932_/B _3864_/C _5499_/Q vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__a22o_1
XFILLER_270_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5068_ _3790_/X _5065_/X _5067_/Y vssd1 vssd1 vccd1 vccd1 _5068_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_217_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_270_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2636__D _5643_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4019_ _5477_/Q _3532_/X _3579_/X vssd1 vssd1 vccd1 vccd1 _4034_/A sky130_fd_sc_hd__a21o_4
XFILLER_270_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2933__B _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3051__A1 _2852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5645__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4876__A _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3780__A _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input33_A i_req_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_234 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_231_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3042__A1 _2840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3593__A2 _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4370_ _4370_/A _4370_/B _4387_/A vssd1 vssd1 vccd1 vccd1 _4371_/C sky130_fd_sc_hd__or3_1
XFILLER_171_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3321_ _3799_/A _2928_/A _3795_/B _3281_/A _3278_/Y vssd1 vssd1 vccd1 vccd1 _3321_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4786__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3252_ _4987_/A _3252_/B vssd1 vssd1 vccd1 vccd1 _5741_/D sky130_fd_sc_hd__nor2_1
XFILLER_224_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4845__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3183_ _5667_/Q _3137_/X _3139_/X _5587_/Q vssd1 vssd1 vccd1 vccd1 _3183_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2737__C _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_226_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3805__A0 _5470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4716__A1_N input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2753__B _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5518__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4026__A _4034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3568__C _5644_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3569__C1 _3567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5755_ _5756_/CLK _5755_/D vssd1 vssd1 vccd1 vccd1 _5755_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3033__A1 _2845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2967_ _2967_/A vssd1 vssd1 vccd1 vccd1 _2969_/B sky130_fd_sc_hd__inv_2
XFILLER_194_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3865__A _3905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4706_ _5559_/Q _4697_/A _4705_/Y _4670_/X vssd1 vssd1 vccd1 vccd1 _5559_/D sky130_fd_sc_hd__o211a_1
X_5686_ _5686_/CLK _5686_/D vssd1 vssd1 vccd1 vccd1 _5686_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5668__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2898_ _2949_/B _3284_/B vssd1 vssd1 vccd1 vccd1 _2899_/A sky130_fd_sc_hd__or2_1
XFILLER_147_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4637_ _5527_/Q _5294_/A _4634_/A _4636_/X vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__a211o_1
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3336__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4568_ _5767_/A _4577_/C vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__or2_1
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3519_ _5439_/Q input45/X _3523_/S vssd1 vssd1 vccd1 vccd1 _3520_/A sky130_fd_sc_hd__mux2_1
X_4499_ _4543_/B _4499_/B vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__xor2_1
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5291__S _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4297__B1 _5453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2928__B _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3105__A _5708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2647__C _5659_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_217_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3272__A1 _5347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3775__A _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4772__A1 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4827__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5214__B _5214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_i_clk clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5743_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3870_ _3935_/A _3874_/B vssd1 vssd1 vccd1 vccd1 _3870_/Y sky130_fd_sc_hd__nand2_1
XFILLER_204_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ _2821_/A _4988_/B vssd1 vssd1 vccd1 vccd1 _3228_/A sky130_fd_sc_hd__nor2_2
XANTENNA__4212__A0 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5540_ _5756_/CLK _5540_/D vssd1 vssd1 vccd1 vccd1 _5768_/A sky130_fd_sc_hd__dfxtp_4
X_2752_ _2757_/D _2782_/B _2782_/C _5600_/Q vssd1 vssd1 vccd1 vccd1 _2752_/X sky130_fd_sc_hd__and4b_1
XFILLER_76_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5471_ _5743_/CLK _5471_/D vssd1 vssd1 vccd1 vccd1 _5471_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2683_ _2761_/B vssd1 vssd1 vccd1 vccd1 _2782_/C sky130_fd_sc_hd__buf_4
XFILLER_219_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4422_ _4422_/A _4422_/B _4422_/C vssd1 vssd1 vccd1 vccd1 _4422_/X sky130_fd_sc_hd__or3_1
XFILLER_117_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4515__A1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4353_ _3617_/A _4121_/B _4271_/A vssd1 vssd1 vccd1 vccd1 _4355_/B sky130_fd_sc_hd__o21ai_1
X_3304_ _3304_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3800_/D sky130_fd_sc_hd__nor2_1
X_4284_ _5449_/Q _4278_/C _4281_/X _5453_/Q _4283_/X vssd1 vssd1 vccd1 vccd1 _4284_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4818__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3235_ _5459_/Q vssd1 vssd1 vccd1 vccd1 _4599_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4374__S0 _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ _5631_/Q _3143_/X _3145_/X _3165_/X vssd1 vssd1 vccd1 vccd1 _3166_/X sky130_fd_sc_hd__a211o_1
XFILLER_239_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5340__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3097_ _5704_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3098_/A sky130_fd_sc_hd__and2_1
XFILLER_199_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5490__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3999_ _4045_/A vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__inv_2
XANTENNA__3595__A _4128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3557__A2 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4754__A1 _5576_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5738_ _5738_/CLK _5738_/D vssd1 vssd1 vccd1 vccd1 _5738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5675_/CLK _5669_/D vssd1 vssd1 vccd1 vccd1 _5669_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_276_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4506__A1 _4504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3190__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5315__A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4809__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_260_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3796__A2 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3001__C _3001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2737__A_N _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2840__C _2840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5209__B _5214_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output187_A _5485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5170__A1 _5169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3181__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__A _5225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output64_A _3227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5363__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3020_ _3019_/X _2840_/A _3089_/A vssd1 vssd1 vccd1 vccd1 _3020_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4971_ _5668_/Q _4972_/B _4970_/Y _4957_/X vssd1 vssd1 vccd1 vccd1 _5668_/D sky130_fd_sc_hd__o211a_1
XFILLER_221_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3787__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4984__A1 _5674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3922_ _5253_/S _3984_/S _3851_/B vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__a21o_2
XFILLER_189_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2995__B1 _2850_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3853_ _5722_/Q vssd1 vssd1 vccd1 vccd1 _3853_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2804_ _5680_/Q _5681_/Q _5682_/Q _5683_/Q _2771_/A _2771_/B vssd1 vssd1 vccd1 vccd1
+ _2805_/B sky130_fd_sc_hd__mux4_1
XANTENNA__4736__A1 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3784_ _4600_/A _3319_/A _3813_/S vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__mux2_1
X_2735_ _2789_/C _2789_/B _2774_/C _5634_/Q vssd1 vssd1 vccd1 vccd1 _2735_/X sky130_fd_sc_hd__and4b_1
X_5523_ _5740_/CLK _5523_/D vssd1 vssd1 vccd1 vccd1 _5523_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4023__B _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5454_ _5692_/CLK _5454_/D vssd1 vssd1 vccd1 vccd1 _5454_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_246_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2666_ _5641_/Q _2655_/X _2657_/X _5673_/Q vssd1 vssd1 vccd1 vccd1 _2666_/X sky130_fd_sc_hd__a22o_1
X_4405_ _4405_/A _4405_/B vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__and2_2
XANTENNA__5706__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5385_ _5404_/CLK _5385_/D vssd1 vssd1 vccd1 vccd1 _5385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3354__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4336_ _4335_/X _4087_/A _4350_/A vssd1 vssd1 vccd1 vccd1 _4337_/B sky130_fd_sc_hd__o21ai_1
XFILLER_259_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4267_ _4304_/S _3635_/Y _4266_/X vssd1 vssd1 vccd1 vccd1 _4267_/X sky130_fd_sc_hd__o21ba_1
XFILLER_113_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4974__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3218_ _5674_/Q _3137_/A _3139_/A _5594_/Q vssd1 vssd1 vccd1 vccd1 _3218_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4672__A0 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4198_ _4471_/S _4469_/D _4198_/C vssd1 vssd1 vccd1 vccd1 _4199_/B sky130_fd_sc_hd__and3_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4693__B _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _3149_/A vssd1 vssd1 vccd1 vccd1 _3149_/X sky130_fd_sc_hd__buf_4
XFILLER_199_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3227__A1 _5563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4975__A1 _5670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2986__B1 _2840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3529__S _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2660__C _5658_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4868__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5386__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3163__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_196 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2835__C _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3218__A1 _5674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3218__B2 _5594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3012__B _5678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4966__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3439__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4124__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2729__B1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5729__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5623_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3154__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5170_ _5713_/Q _5169_/Y _5233_/S vssd1 vssd1 vccd1 vccd1 _5171_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_268_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4121_ _4454_/A _4121_/B vssd1 vssd1 vccd1 vccd1 _4121_/X sky130_fd_sc_hd__or2_1
XFILLER_268_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3902__S _3905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _4052_/A _4052_/B vssd1 vssd1 vccd1 vccd1 _4059_/C sky130_fd_sc_hd__and2_1
XFILLER_232_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3457__A1 _3346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 dbg_in[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_83_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3003_ _3003_/A _3003_/B _3003_/C vssd1 vssd1 vccd1 vccd1 _3004_/C sky130_fd_sc_hd__or3_1
XFILLER_232_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_224_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3209__A1 _5608_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4018__B _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3209__B2 _5624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2680__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3614__D1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4954_ _5661_/Q _4985_/B vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__or2_1
XFILLER_196_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3905_ _5506_/Q _5325_/A _3905_/S vssd1 vssd1 vccd1 vccd1 _3906_/B sky130_fd_sc_hd__mux2_1
X_4885_ _5632_/Q _4894_/A vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__or2_1
XFILLER_189_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4034__A _4034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3576__C _4050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3836_ _5485_/Q _5389_/Q _5242_/S vssd1 vssd1 vccd1 vccd1 _3837_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3767_ _4987_/A _3767_/B vssd1 vssd1 vccd1 vccd1 _5443_/D sky130_fd_sc_hd__nor2_1
X_5506_ _5740_/CLK _5506_/D vssd1 vssd1 vccd1 vccd1 _5506_/Q sky130_fd_sc_hd__dfxtp_1
X_2718_ _2771_/A _2771_/B _5652_/Q _2806_/A vssd1 vssd1 vccd1 vccd1 _2718_/X sky130_fd_sc_hd__and4b_1
XANTENNA__4688__B _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3698_ _5625_/Q _3597_/X _3598_/X _5609_/Q _3697_/X vssd1 vssd1 vccd1 vccd1 _3698_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3592__B _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5134__A1 _2743_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5437_ _5441_/CLK _5437_/D vssd1 vssd1 vccd1 vccd1 _5437_/Q sky130_fd_sc_hd__dfxtp_1
X_2649_ _5563_/Q _2791_/B _2642_/X _2648_/X vssd1 vssd1 vccd1 vccd1 _4635_/B sky130_fd_sc_hd__o22ai_4
XFILLER_273_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5368_ _5757_/CLK _5368_/D vssd1 vssd1 vccd1 vccd1 _5368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4319_ _4300_/S _4396_/B _4318_/X vssd1 vssd1 vccd1 vccd1 _4320_/B sky130_fd_sc_hd__o21a_1
X_5299_ _5067_/B _5743_/Q _5325_/B vssd1 vssd1 vccd1 vccd1 _5300_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4209__A _4503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4643__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4948__A1 _5659_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__C1 _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4176__A2 _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4879__A _5629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3783__A _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4119__A _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_280_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_261_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2862__A _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3677__B _3751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3611__A1 _5563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5551__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4670_ _5331_/A vssd1 vssd1 vccd1 vccd1 _4670_/X sky130_fd_sc_hd__buf_2
XFILLER_186_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3621_ _3732_/A vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3552_ _3585_/B _3948_/A _3551_/Y vssd1 vssd1 vccd1 vccd1 _4030_/A sky130_fd_sc_hd__o21ai_4
X_3483_ _3483_/A vssd1 vssd1 vccd1 vccd1 _5421_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3127__A0 _5711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5222_ _5221_/X _5325_/A _5464_/Q vssd1 vssd1 vccd1 vccd1 _5222_/X sky130_fd_sc_hd__mux2_1
X_5153_ _5155_/B _5142_/B _5155_/A vssd1 vssd1 vccd1 vccd1 _5153_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_229_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4104_ _4363_/A _4105_/B _4377_/A vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__a21oi_2
XFILLER_243_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4627__A0 _5526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5084_ _5514_/Q _3931_/A _5055_/X _5490_/Q vssd1 vssd1 vccd1 vccd1 _5084_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_256_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5132__B _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4035_ _4028_/X _4032_/X _4033_/X _4034_/X vssd1 vssd1 vccd1 vccd1 _4036_/B sky130_fd_sc_hd__a211o_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4029__A _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2653__A2 _2635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2772__A _5614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _4974_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4937_/Y sky130_fd_sc_hd__nand2_1
XFILLER_268_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4868_ _4981_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4868_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3819_ _3819_/A vssd1 vssd1 vccd1 vccd1 _5476_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3807__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4799_ _5683_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4799_/Y sky130_fd_sc_hd__nand2_8
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4563__C1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput160 _5757_/Q vssd1 vssd1 vccd1 vccd1 o_mem_req sky130_fd_sc_hd__buf_2
XANTENNA__3669__A1 _5549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput171 _3023_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[1] sky130_fd_sc_hd__buf_2
Xoutput182 _5480_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[10] sky130_fd_sc_hd__buf_2
Xoutput193 _5476_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[6] sky130_fd_sc_hd__buf_2
XANTENNA__2947__A _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5323__A _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5424__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4618__A0 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4094__A1 _4034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4881__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5574__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4397__A2 _4396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4149__A2 _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4402__A _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4121__B _4121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3018__A _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater215_A _5539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2857__A _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2883__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3688__A _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5771_ _5771_/A vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__clkbuf_1
X_2983_ _2978_/Y _2850_/B _2845_/B _2977_/Y _2982_/X vssd1 vssd1 vccd1 vccd1 _2983_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4722_ _4722_/A _4985_/A vssd1 vssd1 vccd1 vccd1 _4722_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4653_ _4653_/A vssd1 vssd1 vccd1 vccd1 _4653_/X sky130_fd_sc_hd__buf_4
XFILLER_147_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3348__B1 _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput40 i_req_data[24] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3604_ _5627_/Q _3597_/X _3598_/X _5611_/Q _3603_/X vssd1 vssd1 vccd1 vccd1 _3604_/X
+ sky130_fd_sc_hd__a221o_1
Xinput51 i_req_data[5] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3899__A1 _5321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4584_ _5521_/Q _4583_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _4585_/B sky130_fd_sc_hd__mux2_1
X_3535_ _4083_/A vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__buf_4
XANTENNA__4031__B _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5447__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3466_ _3466_/A vssd1 vssd1 vccd1 vccd1 _5413_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3260__B1_N _5528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5205_ _5525_/Q _3932_/B _3864_/C _5505_/Q _5053_/X vssd1 vssd1 vccd1 vccd1 _5205_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3362__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3397_ _2840_/B _5378_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3398_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_229_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5136_ _5136_/A vssd1 vssd1 vccd1 vccd1 _5710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5067_ _5179_/S _5067_/B vssd1 vssd1 vccd1 vccd1 _5067_/Y sky130_fd_sc_hd__nand2_1
XFILLER_284_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_244_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_244_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _4030_/A _4063_/A vssd1 vssd1 vccd1 vccd1 _4087_/A sky130_fd_sc_hd__xor2_4
XFILLER_270_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3598__A _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2933__C _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3587__B1 _3584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5328__A1 _2650_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5053__A _5471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A i_req_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4892__A _5635_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5016__A0 _5689_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4116__B _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3593__A3 _4301_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3447__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4132__A _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3320_ _3281_/A _3283_/B _3308_/D _3282_/B vssd1 vssd1 vccd1 vccd1 _3322_/B sky130_fd_sc_hd__a211o_1
XANTENNA__4786__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3690__B _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3251_ _3245_/Y _3248_/X _3250_/X vssd1 vssd1 vccd1 vccd1 _3252_/B sky130_fd_sc_hd__o21ba_1
XFILLER_224_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3182_ _5554_/Q _3131_/X _3179_/X _3181_/X vssd1 vssd1 vccd1 vccd1 _3182_/X sky130_fd_sc_hd__o22a_1
XFILLER_224_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2737__D _5602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_240_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5007__A0 _5686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4307__A _4307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2753__C _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4026__B _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3568__D _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3569__B1 _3606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5754_ _5754_/CLK _5754_/D vssd1 vssd1 vccd1 vccd1 _5754_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4230__A1 _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ _2966_/A vssd1 vssd1 vccd1 vccd1 _2966_/Y sky130_fd_sc_hd__inv_2
X_4705_ _4722_/A _4976_/A vssd1 vssd1 vccd1 vccd1 _4705_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3584__A3 _2711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5685_ _5685_/CLK _5685_/D vssd1 vssd1 vccd1 vccd1 _5685_/Q sky130_fd_sc_hd__dfxtp_2
X_2897_ _5364_/Q _5363_/Q _5362_/Q vssd1 vssd1 vccd1 vccd1 _3284_/B sky130_fd_sc_hd__or3_4
XANTENNA__4042__A _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4636_ _4635_/A _4482_/B _4635_/Y _5229_/S vssd1 vssd1 vccd1 vccd1 _4636_/X sky130_fd_sc_hd__o211a_1
XFILLER_162_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4567_ _5767_/A _4577_/C vssd1 vssd1 vccd1 vccd1 _4567_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3881__A _3956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3741__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3518_ _3518_/A vssd1 vssd1 vccd1 vccd1 _5438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4498_ _4498_/A _4498_/B vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__xnor2_1
XFILLER_143_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3449_ _5404_/Q _3087_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3450_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3105__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2647__D _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5119_ _5131_/A _5131_/B vssd1 vssd1 vccd1 vccd1 _5119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_214_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3820__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4651__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5612__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4772__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5048__A _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2783__A1 _5613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4509__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3791__A _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3015__B _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5230__B _5230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4460__A1 _5528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2870__A _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2820_ _2803_/X _2817_/X _5331_/B _2821_/A input4/X vssd1 vssd1 vccd1 vccd1 _4988_/B
+ sky130_fd_sc_hd__a2111oi_4
XANTENNA__4748__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2751_ _2751_/A vssd1 vssd1 vccd1 vccd1 _5307_/A sky130_fd_sc_hd__buf_4
XANTENNA__3971__A0 _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5470_ _5743_/CLK _5470_/D vssd1 vssd1 vccd1 vccd1 _5470_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_184_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2682_ _2682_/A vssd1 vssd1 vccd1 vccd1 _2782_/B sky130_fd_sc_hd__buf_4
X_4421_ _4422_/A _4422_/B _4422_/C vssd1 vssd1 vccd1 vccd1 _4421_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4797__A _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3905__S _3905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3723__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4352_ _4352_/A _4352_/B vssd1 vssd1 vccd1 vccd1 _4352_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4920__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3303_ _3295_/Y _5366_/Q _3290_/Y _3795_/A _5340_/Q vssd1 vssd1 vccd1 vccd1 _5340_/D
+ sky130_fd_sc_hd__a32o_1
X_4283_ _5450_/Q _4229_/A _3692_/X _4281_/A _4282_/X vssd1 vssd1 vccd1 vccd1 _4283_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_140_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2684__B_N _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3234_ _5300_/A vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__buf_4
XFILLER_140_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4374__S1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3165_ _5647_/Q _3147_/X _3149_/X _5567_/Q vssd1 vssd1 vccd1 vccd1 _3165_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3096_ _3096_/A vssd1 vssd1 vccd1 vccd1 _3096_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4451__A1 _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5635__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3876__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4471__S _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3998_ _5467_/Q _4289_/C _5291_/S vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__o21a_2
XFILLER_210_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4754__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5737_ _5738_/CLK _5737_/D vssd1 vssd1 vccd1 vccd1 _5737_/Q sky130_fd_sc_hd__dfxtp_1
X_2949_ _2949_/A _2949_/B vssd1 vssd1 vccd1 vccd1 _2949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5668_ _5675_/CLK _5668_/D vssd1 vssd1 vccd1 vccd1 _5668_/Q sky130_fd_sc_hd__dfxtp_4
X_4619_ _5525_/Q _4619_/B vssd1 vssd1 vccd1 vccd1 _4619_/Y sky130_fd_sc_hd__nand2_2
X_5599_ _5738_/CLK _5599_/D vssd1 vssd1 vccd1 vccd1 _5599_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3714__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4500__A _4500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4911__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3190__A1 _5652_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3190__B2 _5572_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5331__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2840__D _2840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4700__A1_N input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3705__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4902__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3181__A1 _5634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5225__B _5225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5508__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3026__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_283_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2865__A _5678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5658__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4970_ _4970_/A _4972_/B vssd1 vssd1 vccd1 vccd1 _4970_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4433__A1 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3921_ _3989_/S vssd1 vssd1 vccd1 vccd1 _3984_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__4984__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3852_ _3893_/A _3856_/C _3919_/A _5488_/Q vssd1 vssd1 vccd1 vccd1 _5488_/D sky130_fd_sc_hd__a22o_1
XFILLER_149_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2803_ _5720_/Q _5442_/Q vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__or2b_1
XANTENNA__4736__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3783_ _4635_/A vssd1 vssd1 vccd1 vccd1 _4600_/A sky130_fd_sc_hd__buf_4
X_5522_ _5740_/CLK _5522_/D vssd1 vssd1 vccd1 vccd1 _5522_/Q sky130_fd_sc_hd__dfxtp_1
X_2734_ _2747_/D vssd1 vssd1 vccd1 vccd1 _2774_/C sky130_fd_sc_hd__buf_8
X_5453_ _5692_/CLK _5453_/D vssd1 vssd1 vccd1 vccd1 _5453_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2665_ _5577_/Q _2644_/X _2664_/X _5609_/Q vssd1 vssd1 vccd1 vccd1 _2665_/X sky130_fd_sc_hd__a22o_1
XFILLER_160_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4404_ _4419_/A _4418_/A vssd1 vssd1 vccd1 vccd1 _4405_/B sky130_fd_sc_hd__or2_1
XANTENNA__4320__A _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5384_ _5722_/CLK _5384_/D vssd1 vssd1 vccd1 vccd1 _5384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3172__A1 _5552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4335_ _4010_/X _4016_/X _4084_/B vssd1 vssd1 vccd1 vccd1 _4335_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4266_ _4304_/S _4303_/A _3662_/X _3617_/A vssd1 vssd1 vccd1 vccd1 _4266_/X sky130_fd_sc_hd__a31o_1
XFILLER_140_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4974__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3217_ _5561_/Q _3131_/A _3214_/X _3216_/X vssd1 vssd1 vccd1 vccd1 _3217_/X sky130_fd_sc_hd__o22a_2
XFILLER_274_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4672__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4197_ _4099_/X _4195_/X _4196_/Y vssd1 vssd1 vccd1 vccd1 _4208_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3148_ input3/X input2/X input1/X vssd1 vssd1 vccd1 vccd1 _3149_/A sky130_fd_sc_hd__nor3b_4
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _5403_/Q _3079_/B vssd1 vssd1 vccd1 vccd1 _3084_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3227__A2 _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4975__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2738__A1 _5618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2660__D _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5685_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3163__A1 _5663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4360__B1 _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3163__B2 _5583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2910__A1 _2943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2910__B2 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3871__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3218__A2 _3137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4966__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2729__A1 _5587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3926__A0 _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_60_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3455__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3154__A1 _5597_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4351__B1 _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3154__B2 _5613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2901__A1 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4120_ _4229_/A _4221_/A _4221_/B _4307_/A _4119_/Y vssd1 vssd1 vccd1 vccd1 _4121_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5480__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_315 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4051_ _4403_/B vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__clkinv_2
XFILLER_209_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 i_irq vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_3002_ _2962_/Y _2850_/C _2830_/Y _3001_/X vssd1 vssd1 vccd1 vccd1 _3002_/X sky130_fd_sc_hd__o211a_1
XFILLER_232_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2665__B1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3209__A2 _3133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4953_ _4646_/X _4949_/Y _4952_/X _4933_/X vssd1 vssd1 vccd1 vccd1 _5660_/D sky130_fd_sc_hd__o211a_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3904_ _3904_/A vssd1 vssd1 vccd1 vccd1 _5505_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4315__A _4496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3090__B1 _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4884_ _4663_/X _4874_/Y _4883_/X _4862_/X vssd1 vssd1 vccd1 vccd1 _5631_/D sky130_fd_sc_hd__o211a_1
XFILLER_189_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3835_ _3835_/A vssd1 vssd1 vccd1 vccd1 _5484_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4034__B _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3917__B1 _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3766_ _4529_/A _3764_/X _3765_/Y _3843_/B vssd1 vssd1 vccd1 vccd1 _3767_/B sky130_fd_sc_hd__o211a_1
XFILLER_257_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5505_ _5740_/CLK _5505_/D vssd1 vssd1 vccd1 vccd1 _5505_/Q sky130_fd_sc_hd__dfxtp_1
X_2717_ _2806_/A _2771_/A _2775_/B _5588_/Q vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__and4bb_1
XFILLER_133_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3697_ _5673_/Q _3600_/X _3602_/X _5657_/Q vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3592__C _4408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4050__A _4050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5436_ _5441_/CLK _5436_/D vssd1 vssd1 vccd1 vccd1 _5436_/Q sky130_fd_sc_hd__dfxtp_1
X_2648_ _5579_/Q _2644_/X _2645_/X _2686_/A _2647_/X vssd1 vssd1 vccd1 vccd1 _2648_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4342__B1 _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5367_ _5716_/CLK _5367_/D vssd1 vssd1 vccd1 vccd1 _5367_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4985__A _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4893__A1 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4318_ _4469_/D _4317_/X _4248_/X _4396_/A vssd1 vssd1 vccd1 vccd1 _4318_/X sky130_fd_sc_hd__a211o_1
XFILLER_259_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5298_ _4619_/B _3843_/B _5294_/B vssd1 vssd1 vccd1 vccd1 _5325_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4249_ _4469_/D _4247_/X _4248_/X vssd1 vssd1 vccd1 vccd1 _4250_/B sky130_fd_sc_hd__a21oi_1
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4948__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5353__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4879__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input56_A i_req_data_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4895__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4884__A1 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3304__A _3304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4636__A1 _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4119__B _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output212_A _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4135__A _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__B1 _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3611__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3620_ _3747_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3732_/A sky130_fd_sc_hd__nor2_2
XANTENNA__4572__B1 _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3551_ _5474_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _3551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3482_ _5421_/Q input26/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__mux2_1
X_5221_ _4457_/D _5220_/Y _5231_/S vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5152_ _5148_/Y _5151_/X _5219_/S vssd1 vssd1 vccd1 vccd1 _5155_/A sky130_fd_sc_hd__mux2_1
XFILLER_229_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4103_ _4103_/A _4103_/B vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__nand2_2
XFILLER_243_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5083_ _5487_/Q _3840_/A _5051_/B _5530_/Q vssd1 vssd1 vccd1 vccd1 _5083_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_110_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2756__C _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4034_ _4034_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4034_/X sky130_fd_sc_hd__and2_1
XFILLER_49_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4029__B _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5376__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5052__A1 _5508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5052__B2 _5492_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4936_ _5653_/Q _4935_/B _4935_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5653_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4045__A _4045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_130 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_268_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4867_ _5624_/Q _4859_/B _4866_/Y _4862_/X vssd1 vssd1 vccd1 vccd1 _5624_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3884__A _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3818_ _5476_/Q _5380_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3819_/A sky130_fd_sc_hd__mux2_1
X_4798_ _5595_/Q _4784_/B _4797_/Y _4791_/X vssd1 vssd1 vccd1 vccd1 _5595_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3366__A1 _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3749_ _3733_/X _3748_/X _4454_/B vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5419_ _5757_/CLK _5419_/D vssd1 vssd1 vccd1 vccd1 _5419_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput150 _3128_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[15] sky130_fd_sc_hd__buf_2
Xoutput161 _3113_/S vssd1 vssd1 vccd1 vccd1 o_mem_sel[0] sky130_fd_sc_hd__buf_2
XANTENNA__3669__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 _3029_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[2] sky130_fd_sc_hd__buf_2
Xoutput183 _5481_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[11] sky130_fd_sc_hd__buf_2
Xoutput194 _5477_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_101_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4618__A1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5291__A1 _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5719__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3841__A2 _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5658_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2902__S _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4402__B _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output162_A _3096_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3733__S _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5282__A1 _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2873__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3688__B _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _5770_/A vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4388__A3 _4041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2982_ _2978_/Y _2850_/B _2840_/A _2979_/Y _2981_/X vssd1 vssd1 vccd1 vccd1 _2982_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ input13/X _4689_/X _4690_/X _4720_/Y vssd1 vssd1 vccd1 vccd1 _4985_/A sky130_fd_sc_hd__o2bb2a_4
X_4652_ _5705_/Q _4651_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3348__A1 _5357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 i_req_data[15] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
X_3603_ _5675_/Q _3600_/X _3602_/X _5659_/Q vssd1 vssd1 vccd1 vccd1 _3603_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4545__B1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput41 i_req_data[25] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
X_4583_ _5315_/A _4362_/A _4626_/S vssd1 vssd1 vccd1 vccd1 _4583_/X sky130_fd_sc_hd__mux2_1
Xinput52 i_req_data[6] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3534_ _3532_/X _4523_/B _3533_/Y vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__o21a_2
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3465_ _5413_/Q input49/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5204_ _5204_/A vssd1 vssd1 vccd1 vccd1 _5716_/D sky130_fd_sc_hd__clkbuf_1
X_3396_ _3419_/S vssd1 vssd1 vccd1 vccd1 _3415_/S sky130_fd_sc_hd__buf_4
XFILLER_254_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5135_ _5710_/Q _5134_/X _5135_/S vssd1 vssd1 vccd1 vccd1 _5136_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5066_ _5464_/Q vssd1 vssd1 vccd1 vccd1 _5179_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__5273__A1 _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3879__A _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4017_ _4067_/A _4232_/B vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__xor2_4
XFILLER_84_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4481__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_225_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3587__A1 _5479_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4919_ _5646_/Q _4947_/B vssd1 vssd1 vccd1 vccd1 _4919_/X sky130_fd_sc_hd__or2_1
XANTENNA__3818__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4503__A _4503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5541__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4892__B _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5264__A1 _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input19_A i_mem_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2693__A _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5691__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3578__A1 _5480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3593__A4 _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4132__B _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output87_A _3167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2868__A _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3463__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3690__C _3690_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3250_ _3250_/A _3270_/C _3270_/D _3250_/D vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__and4_1
XFILLER_3_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3181_ _5634_/Q _3143_/X _3145_/X _3180_/X vssd1 vssd1 vccd1 vccd1 _3181_/X sky130_fd_sc_hd__a211o_1
XFILLER_78_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4058__A2 _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3266__B1 _5347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4307__B _4307_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2753__D _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4215__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3569__A1 _5564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5753_ _5754_/CLK _5753_/D vssd1 vssd1 vccd1 vccd1 _5753_/Q sky130_fd_sc_hd__dfxtp_1
X_2965_ _5402_/Q vssd1 vssd1 vccd1 vccd1 _2965_/Y sky130_fd_sc_hd__inv_2
X_4704_ input9/X _4689_/X _4690_/X _4703_/Y vssd1 vssd1 vccd1 vccd1 _4976_/A sky130_fd_sc_hd__o2bb2a_4
X_5684_ _5686_/CLK _5684_/D vssd1 vssd1 vccd1 vccd1 _5684_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5414__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2896_ _3281_/C vssd1 vssd1 vccd1 vccd1 _3775_/C sky130_fd_sc_hd__buf_2
X_4635_ _4635_/A _4635_/B vssd1 vssd1 vccd1 vccd1 _4635_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4042__B _4363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4566_ _5766_/A _4511_/X _3919_/A _4565_/X vssd1 vssd1 vccd1 vccd1 _5538_/D sky130_fd_sc_hd__o211a_1
XFILLER_265_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3741__A1 _5671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3881__B _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3517_ _5438_/Q input44/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3518_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5564__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2778__A _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4497_ _4537_/B _4522_/B vssd1 vssd1 vccd1 vccd1 _4498_/B sky130_fd_sc_hd__xor2_1
XANTENNA__3373__S _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3448_ _3448_/A vssd1 vssd1 vccd1 vccd1 _5403_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4151__D1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ input28/X _5423_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3379_/X sky130_fd_sc_hd__mux2_1
XFILLER_281_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5114_/Y _5117_/X _5219_/S vssd1 vssd1 vccd1 vccd1 _5131_/B sky130_fd_sc_hd__mux2_1
XFILLER_281_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5049_ _5055_/A _3838_/C _3996_/B _5460_/Q vssd1 vssd1 vccd1 vccd1 _5125_/A sky130_fd_sc_hd__a31o_2
XFILLER_27_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3272__A3 _3267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_213_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5329__A _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3775__C _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5048__B _5462_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4509__B1 _4507_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3980__A1 _5321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2783__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2688__A _5559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4408__A _4408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output125_A _5557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5003__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4460__A2 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5437__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_231_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2750_ _2744_/X _2745_/X _2748_/X _2749_/X vssd1 vssd1 vccd1 vccd1 _2751_/A sky130_fd_sc_hd__o31a_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5587__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2681_ _2681_/A vssd1 vssd1 vccd1 vccd1 _2757_/D sky130_fd_sc_hd__buf_4
XFILLER_129_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_5_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4420_ _4483_/B _4420_/B vssd1 vssd1 vccd1 vccd1 _4422_/C sky130_fd_sc_hd__xnor2_1
XFILLER_184_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4797__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3723__A1 _5573_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ _4087_/B _4339_/S _4087_/A vssd1 vssd1 vccd1 vccd1 _4352_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3302_ _3295_/Y _3300_/X _3293_/X _5339_/Q vssd1 vssd1 vccd1 vccd1 _5339_/D sky130_fd_sc_hd__a2bb2o_1
X_4282_ _4229_/A _4281_/A _5452_/Q vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__o21a_1
X_3233_ _3233_/A vssd1 vssd1 vccd1 vccd1 _3250_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3164_ _5599_/Q _3133_/X _3135_/X _5615_/Q _3163_/X vssd1 vssd1 vccd1 vccd1 _3164_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5228__A1 _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3095_ _5688_/Q _5677_/Q vssd1 vssd1 vccd1 vccd1 _3096_/A sky130_fd_sc_hd__or2b_1
XFILLER_254_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3876__B _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3368__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3997_ _5461_/Q _5051_/B vssd1 vssd1 vccd1 vccd1 _4289_/C sky130_fd_sc_hd__and2_2
XANTENNA__3411__A0 _2967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5736_ _5738_/CLK _5736_/D vssd1 vssd1 vccd1 vccd1 _5736_/Q sky130_fd_sc_hd__dfxtp_1
X_2948_ _3799_/B _3284_/B _5241_/D vssd1 vssd1 vccd1 vccd1 _3318_/C sky130_fd_sc_hd__o21bai_4
XFILLER_210_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_276_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3962__A1 _5519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4988__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5667_ _5667_/CLK _5667_/D vssd1 vssd1 vccd1 vccd1 _5667_/Q sky130_fd_sc_hd__dfxtp_4
X_2879_ _2879_/A vssd1 vssd1 vccd1 vccd1 _3799_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_276_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4618_ _5323_/A _4617_/Y _4626_/S vssd1 vssd1 vccd1 vccd1 _4618_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5598_ _5598_/CLK _5598_/D vssd1 vssd1 vccd1 vccd1 _5598_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_135_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3714__A1 _5578_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3714__B2 _5594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4549_ _4552_/B _4511_/X _4545_/Y _4548_/X _3919_/X vssd1 vssd1 vccd1 vccd1 _5536_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4500__B _5015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3190__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5331__B _5331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4228__A _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4662__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3705__A1 _5624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3705__B2 _5608_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3307__A _3307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3181__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2865__B _5300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__A2 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4138__A _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2881__A _5361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3920_ _5511_/Q _3918_/B _3918_/Y _3919_/X vssd1 vssd1 vccd1 vccd1 _5511_/D sky130_fd_sc_hd__o211a_1
XFILLER_189_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3641__B1 _3608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3851_ _5300_/A _3851_/B vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__nor2_4
X_2802_ _5678_/Q _3851_/B _2802_/C vssd1 vssd1 vccd1 vccd1 _2821_/A sky130_fd_sc_hd__or3_2
X_3782_ _5461_/Q vssd1 vssd1 vccd1 vccd1 _4635_/A sky130_fd_sc_hd__buf_4
XFILLER_157_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5521_ _5740_/CLK _5521_/D vssd1 vssd1 vccd1 vccd1 _5521_/Q sky130_fd_sc_hd__dfxtp_2
X_2733_ _2733_/A vssd1 vssd1 vccd1 vccd1 _2789_/B sky130_fd_sc_hd__buf_8
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5146__A0 _5711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5452_ _5528_/CLK _5452_/D vssd1 vssd1 vccd1 vccd1 _5452_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2664_ _2681_/A _2733_/A _2747_/B vssd1 vssd1 vccd1 vccd1 _2664_/X sky130_fd_sc_hd__and3b_4
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4403_ _4403_/A _4403_/B vssd1 vssd1 vccd1 vccd1 _4403_/X sky130_fd_sc_hd__or2_1
XFILLER_172_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5383_ _5404_/CLK _5383_/D vssd1 vssd1 vccd1 vccd1 _5383_/Q sky130_fd_sc_hd__dfxtp_1
X_4334_ _4320_/Y _4332_/X _4438_/B _4071_/B vssd1 vssd1 vccd1 vccd1 _5132_/A sky130_fd_sc_hd__o2bb2a_4
XANTENNA__3172__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4265_ _3733_/X _3647_/Y _4304_/S vssd1 vssd1 vccd1 vccd1 _4265_/X sky130_fd_sc_hd__mux2_1
X_3216_ _5641_/Q _3143_/A _3145_/A _3215_/X vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5602__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2775__B _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4196_ _4099_/X _4195_/X _4483_/A vssd1 vssd1 vccd1 vccd1 _4196_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_274_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3147_ _3147_/A vssd1 vssd1 vccd1 vccd1 _3147_/X sky130_fd_sc_hd__buf_4
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4064__A_N _4024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3078_ _5772_/A _3010_/X _3077_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3078_/X sky130_fd_sc_hd__o211a_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3887__A _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5752__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2791__A _5548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2986__A2 _2852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4188__A1 _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2738__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5719_ _5721_/CLK _5719_/D vssd1 vssd1 vccd1 vccd1 _5719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3826__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4511__A _4581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3699__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4896__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3163__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4360__B2 _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4657__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2966__A _2966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2685__B _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3623__B1 _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_362 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4179__A1 _4148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2729__A2 _2635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output192_A _5475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4887__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3154__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5625__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2901__A2 _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2876__A _3317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3471__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4050_/A _4415_/A vssd1 vssd1 vccd1 vccd1 _4403_/B sky130_fd_sc_hd__and2_1
XFILLER_256_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3001_ _3001_/A _3001_/B _3001_/C _3001_/D vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__or4_2
XANTENNA__3311__C1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput6 i_mem_ack vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2665__A1 _5577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2665__B2 _5609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4952_ _5660_/Q _4985_/B vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__or2_1
XANTENNA__3614__B1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4811__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3903_ _5261_/A _3903_/B vssd1 vssd1 vccd1 vccd1 _3904_/A sky130_fd_sc_hd__and2_1
X_4883_ _5631_/Q _4910_/B vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__or2_1
XFILLER_177_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3090__A1 _2850_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3834_ _5484_/Q _5388_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3835_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3917__A1 _3843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3765_ _4527_/C _4529_/A vssd1 vssd1 vccd1 vccd1 _3765_/Y sky130_fd_sc_hd__nand2_1
XFILLER_192_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3646__S _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2716_ _5636_/Q _2655_/X _2657_/X _5668_/Q vssd1 vssd1 vccd1 vccd1 _2716_/X sky130_fd_sc_hd__a22o_1
XFILLER_257_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5504_ _5740_/CLK _5504_/D vssd1 vssd1 vccd1 vccd1 _5504_/Q sky130_fd_sc_hd__dfxtp_1
X_3696_ _3650_/Y _3675_/X _3678_/Y _3695_/X vssd1 vssd1 vccd1 vccd1 _3696_/X sky130_fd_sc_hd__a31o_1
X_5435_ _5722_/CLK _5435_/D vssd1 vssd1 vccd1 vccd1 _5435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3592__D _4050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4050__B _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2647_ _2733_/A _2747_/B _5659_/Q _2747_/D vssd1 vssd1 vccd1 vccd1 _2647_/X sky130_fd_sc_hd__and4b_1
XFILLER_105_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4878__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4342__A1 _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5366_ _5757_/CLK _5366_/D vssd1 vssd1 vccd1 vccd1 _5366_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4985__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4893__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3696__A3 _3678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4317_ _4151_/X _4154_/X _4447_/S vssd1 vssd1 vccd1 vccd1 _4317_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5297_ _5294_/A _2785_/Y _5294_/B _5296_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5742_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_273_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4248_ _4454_/B _4449_/S _4248_/C vssd1 vssd1 vccd1 vccd1 _4248_/X sky130_fd_sc_hd__and3_1
XFILLER_259_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4179_ _4394_/A _4148_/X _4133_/X _4127_/X _4146_/A _4449_/S vssd1 vssd1 vccd1 vccd1
+ _4180_/B sky130_fd_sc_hd__mux4_1
XFILLER_82_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_255_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5648__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4869__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4895__B _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4884__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2696__A _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A i_req_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4636__A2 _4482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5011__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3072__A1 _2967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3550_ _3550_/A vssd1 vssd1 vccd1 vccd1 _4067_/A sky130_fd_sc_hd__buf_6
XFILLER_127_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3481_ _3481_/A vssd1 vssd1 vccd1 vccd1 _5420_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220_ _5220_/A _5225_/A vssd1 vssd1 vccd1 vccd1 _5220_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_142_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2908__C_N _5362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5151_ _5768_/A _5193_/B _5150_/Y _5196_/A vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__o2bb2a_1
X_4102_ _4102_/A _4102_/B vssd1 vssd1 vccd1 vccd1 _4386_/B sky130_fd_sc_hd__or2_2
X_5082_ _5494_/Q _5082_/B vssd1 vssd1 vccd1 vccd1 _5082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2756__D _5584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4033_ _4033_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4033_/X sky130_fd_sc_hd__and2_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4326__A _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5707_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_252_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4935_ _4972_/A _4935_/B vssd1 vssd1 vccd1 vccd1 _4935_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4045__B _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4260__B1 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4866_ _4978_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_268_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_165_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3817_ _3817_/A vssd1 vssd1 vccd1 vccd1 _5475_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3376__S _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4797_ _4985_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4797_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4563__A1 _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ _3740_/X _3747_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _3748_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3679_ _4302_/S _4076_/A vssd1 vssd1 vccd1 vccd1 _4278_/A sky130_fd_sc_hd__nor2_2
XFILLER_137_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput140 _5695_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[6] sky130_fd_sc_hd__buf_2
X_5418_ _5757_/CLK _5418_/D vssd1 vssd1 vccd1 vccd1 _5418_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput151 _3100_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[1] sky130_fd_sc_hd__buf_2
XFILLER_133_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput162 _3096_/X vssd1 vssd1 vccd1 vccd1 o_mem_sel[1] sky130_fd_sc_hd__buf_2
XFILLER_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput173 _3034_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[3] sky130_fd_sc_hd__buf_2
Xoutput184 _5482_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[12] sky130_fd_sc_hd__buf_2
X_5349_ _5716_/CLK _5349_/D vssd1 vssd1 vccd1 vccd1 _5349_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput195 _5478_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3826__A0 _5480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5470__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5067__A _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3294__A1_N _5365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2873__B _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4146__A _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3050__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2981_ _2979_/Y _2840_/A _2840_/C _2980_/Y vssd1 vssd1 vccd1 vccd1 _2981_/X sky130_fd_sc_hd__a211o_1
XFILLER_159_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _5719_/Q vssd1 vssd1 vccd1 vccd1 _4720_/Y sky130_fd_sc_hd__inv_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_304 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4651_ input22/X input14/X _4651_/S vssd1 vssd1 vccd1 vccd1 _4651_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2717__A_N _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3602_ _3602_/A vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__buf_6
Xinput20 i_mem_data[7] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
Xinput31 i_req_data[16] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4582_ _4529_/X _4580_/X _4581_/X _3919_/X vssd1 vssd1 vccd1 vccd1 _5540_/D sky130_fd_sc_hd__o211a_1
Xinput42 i_req_data[26] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 i_req_data[7] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
XFILLER_162_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3533_ _5472_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _3533_/Y sky130_fd_sc_hd__nand2_2
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3464_ _3464_/A vssd1 vssd1 vccd1 vccd1 _5412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_254_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5203_ _5716_/Q _5202_/X _5233_/S vssd1 vssd1 vccd1 vccd1 _5204_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3395_ _3395_/A vssd1 vssd1 vccd1 vccd1 _5377_/D sky130_fd_sc_hd__clkbuf_1
X_5134_ _5133_/X _2743_/Y _5179_/S vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_229_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5343__CLK _5680_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _5060_/Y _5062_/Y _5200_/B _4500_/A vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_270_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4016_ _4011_/X _4012_/X _4014_/X _4015_/X vssd1 vssd1 vccd1 vccd1 _4016_/X sky130_fd_sc_hd__o31a_2
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5493__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3895__A _5319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3587__A2 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4918_ _4653_/X _4912_/Y _4917_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5645_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4503__B _5156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4849_ _4668_/X _4836_/Y _4848_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5616_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3834__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4395__S0 _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3135__A _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3275__A1 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3578__A2 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_304 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2786__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5366__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3180_ _5650_/Q _3147_/X _3149_/X _5570_/Q vssd1 vssd1 vccd1 vccd1 _3180_/X sky130_fd_sc_hd__a22o_1
XFILLER_224_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4575__S _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2884__A _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_226_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3569__A2 _3607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5752_ _5756_/CLK _5752_/D vssd1 vssd1 vccd1 vccd1 _5752_/Q sky130_fd_sc_hd__dfxtp_1
X_2964_ _5403_/Q vssd1 vssd1 vccd1 vccd1 _2964_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2777__B1 _2770_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4703_ _5715_/Q vssd1 vssd1 vccd1 vccd1 _4703_/Y sky130_fd_sc_hd__inv_2
X_2895_ _5361_/Q _5360_/Q vssd1 vssd1 vccd1 vccd1 _3281_/C sky130_fd_sc_hd__and2_1
X_5683_ _5686_/CLK _5683_/D vssd1 vssd1 vccd1 vccd1 _5683_/Q sky130_fd_sc_hd__dfxtp_2
X_4634_ _4634_/A _4634_/B vssd1 vssd1 vccd1 vccd1 _4634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4565_ _4532_/X _4559_/Y _4560_/X _4564_/Y _4529_/X vssd1 vssd1 vccd1 vccd1 _4565_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5709__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3741__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3516_ _3516_/A vssd1 vssd1 vccd1 vccd1 _5437_/D sky130_fd_sc_hd__clkbuf_1
X_4496_ _4496_/A _5132_/A vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_21_i_clk clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5680_/CLK sky130_fd_sc_hd__clkbuf_16
X_3447_ _5403_/Q _3082_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3448_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3378_ _3378_/A vssd1 vssd1 vccd1 vccd1 _5370_/D sky130_fd_sc_hd__clkbuf_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2794__A _5355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5117_ _5765_/A _5125_/A _5116_/Y _5460_/Q vssd1 vssd1 vccd1 vccd1 _5117_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_245_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5048_ _5196_/A _5462_/Q vssd1 vssd1 vccd1 vccd1 _5156_/B sky130_fd_sc_hd__nor2_4
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4206__B1 _4192_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4514__A _5513_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4509__A1 _5532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5389__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3193__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4390__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2688__B _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2940__A0 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input31_A i_req_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_263_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4408__B _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output118_A _5550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4424__A _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4748__A1 _5573_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5239__B _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2680_ _5639_/Q _2655_/X _2657_/X _5671_/Q vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__a22o_1
XFILLER_144_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5173__A1 _5522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3184__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4350_ _4350_/A _4350_/B _4350_/C vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__and3_1
XANTENNA__4920__A1 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3723__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3301_ _5365_/Q _3300_/X _3293_/X _5338_/Q vssd1 vssd1 vccd1 vccd1 _5338_/D sky130_fd_sc_hd__a2bb2o_1
X_4281_ _4281_/A _4281_/B vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__xor2_1
XFILLER_125_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3232_ _5461_/Q _4988_/B vssd1 vssd1 vccd1 vccd1 _3233_/A sky130_fd_sc_hd__and2_1
XFILLER_239_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3163_ _5663_/Q _3137_/X _3139_/X _5583_/Q vssd1 vssd1 vccd1 vccd1 _3163_/X sky130_fd_sc_hd__a22o_1
XFILLER_254_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3094_ _4651_/S vssd1 vssd1 vccd1 vccd1 _3113_/S sky130_fd_sc_hd__buf_2
XANTENNA__2764__D _5567_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3649__S _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3996_ _5055_/A _3996_/B _5055_/C vssd1 vssd1 vccd1 vccd1 _5051_/B sky130_fd_sc_hd__and3_4
XFILLER_210_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5735_ _5738_/CLK _5735_/D vssd1 vssd1 vccd1 vccd1 _5735_/Q sky130_fd_sc_hd__dfxtp_1
X_2947_ _3799_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _5241_/D sky130_fd_sc_hd__nor2_1
XANTENNA__5531__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5666_ _5747_/CLK _5666_/D vssd1 vssd1 vccd1 vccd1 _5666_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_276_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2878_ _5364_/Q _5362_/Q _5363_/Q vssd1 vssd1 vccd1 vccd1 _2879_/A sky130_fd_sc_hd__or3b_1
XANTENNA__4988__B _4988_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4617_ _4617_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4617_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__5164__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5597_ _5598_/CLK _5597_/D vssd1 vssd1 vccd1 vccd1 _5597_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__3175__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3714__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4911__A1 _5643_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5681__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4548_ _4532_/X _4546_/Y _4547_/X _4529_/A vssd1 vssd1 vccd1 vccd1 _4548_/X sky130_fd_sc_hd__a31o_1
XFILLER_150_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _4523_/B _4485_/A vssd1 vssd1 vccd1 vccd1 _4479_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_225_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3132__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2674__D _5592_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2989__B1 _2845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3166__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4902__A1 _5639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3705__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3307__B _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4666__A0 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_1_0_i_clk_A clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4419__A _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5404__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5091__B1 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2881__B _5360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3641__A1 _5618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3469__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3641__B2 _5586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5554__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _5263_/A vssd1 vssd1 vccd1 vccd1 _3893_/A sky130_fd_sc_hd__clkbuf_4
X_2801_ _5676_/Q _5486_/Q vssd1 vssd1 vccd1 vccd1 _2802_/C sky130_fd_sc_hd__nor2_1
XANTENNA__3929__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3781_ _5196_/A _3780_/A _3780_/Y vssd1 vssd1 vccd1 vccd1 _5460_/D sky130_fd_sc_hd__o21a_1
XANTENNA__3993__A _4635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5520_ _5740_/CLK _5520_/D vssd1 vssd1 vccd1 vccd1 _5520_/Q sky130_fd_sc_hd__dfxtp_2
X_2732_ _2747_/B vssd1 vssd1 vccd1 vccd1 _2789_/C sky130_fd_sc_hd__buf_6
XANTENNA__5146__A1 _5145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5451_ _5692_/CLK _5451_/D vssd1 vssd1 vccd1 vccd1 _5451_/Q sky130_fd_sc_hd__dfxtp_1
X_2663_ _2663_/A vssd1 vssd1 vccd1 vccd1 _5325_/A sky130_fd_sc_hd__buf_4
X_4402_ _4419_/A _4418_/A vssd1 vssd1 vccd1 vccd1 _4405_/A sky130_fd_sc_hd__nand2_1
X_5382_ _5404_/CLK _5382_/D vssd1 vssd1 vccd1 vccd1 _5382_/Q sky130_fd_sc_hd__dfxtp_1
X_4333_ _4333_/A vssd1 vssd1 vccd1 vccd1 _4438_/B sky130_fd_sc_hd__clkinv_2
XFILLER_259_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4264_ _4081_/Y _4258_/X _4261_/Y _4263_/X vssd1 vssd1 vccd1 vccd1 _4269_/A sky130_fd_sc_hd__a211oi_1
XFILLER_262_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4657__A0 _5706_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3215_ _5657_/Q _3147_/A _3149_/A _5577_/Q vssd1 vssd1 vccd1 vccd1 _3215_/X sky130_fd_sc_hd__a22o_1
XFILLER_262_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ _4213_/A _4213_/B _4101_/B vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__2775__C _5646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3146_ input1/X input2/X input3/X vssd1 vssd1 vccd1 vccd1 _3147_/A sky130_fd_sc_hd__and3b_4
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3077_ _2835_/B _3089_/A _3074_/X _3076_/Y _3018_/A vssd1 vssd1 vccd1 vccd1 _3077_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2791__B _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3379__S _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3979_ _5772_/A _5737_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3979_/X sky130_fd_sc_hd__mux2_1
X_5718_ _5757_/CLK _5718_/D vssd1 vssd1 vccd1 vccd1 _5718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5137__A1 _5519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5649_ _5667_/CLK _5649_/D vssd1 vssd1 vccd1 vccd1 _5649_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5137__B2 _5499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3699__A1 _5577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3699__B2 _5593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5427__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3143__A _3143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5577__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4673__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3623__A1 _5617_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__B2 _5601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5128__B2 _5460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output185_A _5483_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2901__A3 _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4639__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output62_A _3217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3311__B1 _3310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3000_ input25/X _5420_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _3001_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 i_mem_data[0] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2665__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4583__S _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_214 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _4969_/A vssd1 vssd1 vccd1 vccd1 _4985_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__3614__A1 _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3902_ _5505_/Q _5323_/A _3905_/S vssd1 vssd1 vccd1 vccd1 _3903_/B sky130_fd_sc_hd__mux2_1
X_4882_ _4658_/X _4874_/Y _4881_/X _4862_/X vssd1 vssd1 vccd1 vccd1 _5630_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3833_ _3833_/A vssd1 vssd1 vccd1 vccd1 _5483_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3927__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2831__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3764_ _4527_/C _3760_/Y _4585_/A vssd1 vssd1 vccd1 vccd1 _3764_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_338 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5503_ _5756_/CLK _5503_/D vssd1 vssd1 vccd1 vccd1 _5503_/Q sky130_fd_sc_hd__dfxtp_1
X_2715_ _5572_/Q _2644_/X _2664_/X _5604_/Q vssd1 vssd1 vccd1 vccd1 _2715_/X sky130_fd_sc_hd__a22o_1
X_3695_ _2936_/X _4278_/A _3686_/Y _3694_/X vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__a211o_1
XFILLER_257_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5434_ _5441_/CLK _5434_/D vssd1 vssd1 vccd1 vccd1 _5434_/Q sky130_fd_sc_hd__dfxtp_1
X_2646_ _2681_/A _2682_/A _2761_/B vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__nor3_4
XFILLER_160_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4342__A2 _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5365_ _5757_/CLK _5365_/D vssd1 vssd1 vccd1 vccd1 _5365_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3662__S _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4316_ _4127_/X _4148_/X _4149_/X _4150_/X _4272_/S _4146_/A vssd1 vssd1 vccd1 vccd1
+ _4396_/B sky130_fd_sc_hd__mux4_2
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5296_ _5742_/Q _3843_/B _5295_/X vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_247_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4247_ _4151_/X _4154_/X _4447_/S vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3302__B1 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4178_ _4176_/Y _4140_/Y _4141_/Y _4177_/Y _4447_/S _4146_/A vssd1 vssd1 vccd1 vccd1
+ _4178_/X sky130_fd_sc_hd__mux4_1
XFILLER_274_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3898__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3129_ input3/X input2/X input1/X vssd1 vssd1 vccd1 vccd1 _3130_/A sky130_fd_sc_hd__or3_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_190 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_248_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3081__A2 _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2773__A_N _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4522__A _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_198 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3138__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4318__C1 _4396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4557__C1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3480_ _5420_/Q input25/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3481_/A sky130_fd_sc_hd__mux2_1
XFILLER_182_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3482__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5742__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5263__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5150_ _5749_/Q _3840_/X _5149_/X vssd1 vssd1 vccd1 vccd1 _5150_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_243_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4101_ _4101_/A _4101_/B vssd1 vssd1 vccd1 vccd1 _4102_/B sky130_fd_sc_hd__nor2_1
XFILLER_256_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5081_ _5081_/A _5125_/A vssd1 vssd1 vccd1 vccd1 _5081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_256_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4032_ _4029_/X _4348_/B _4031_/X vssd1 vssd1 vccd1 vccd1 _4032_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_264_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3048__C1 _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4934_ _5652_/Q _4935_/B _4932_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5652_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4796__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4865_ _5623_/Q _4859_/B _4864_/Y _4862_/X vssd1 vssd1 vccd1 vccd1 _5623_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_220_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3816_ _5475_/Q _5379_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3817_/A sky130_fd_sc_hd__mux2_1
X_4796_ _5594_/Q _4784_/B _4795_/Y _4791_/X vssd1 vssd1 vccd1 vccd1 _5594_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3747_ _3747_/A _3747_/B _4112_/B vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__or3_1
XANTENNA__4563__A2 _3956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3678_ _4116_/A _4326_/A vssd1 vssd1 vccd1 vccd1 _3678_/Y sky130_fd_sc_hd__nor2_2
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5417_ _5757_/CLK _5417_/D vssd1 vssd1 vccd1 vccd1 _5417_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput130 _5699_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[10] sky130_fd_sc_hd__buf_2
XANTENNA__2797__A _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput141 _5696_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[7] sky130_fd_sc_hd__buf_2
XANTENNA__3392__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput152 _3102_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[2] sky130_fd_sc_hd__buf_2
Xoutput163 _5721_/Q vssd1 vssd1 vccd1 vccd1 o_mem_we sky130_fd_sc_hd__buf_2
Xoutput174 _3038_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[4] sky130_fd_sc_hd__buf_2
XFILLER_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5348_ _5721_/CLK _5348_/D vssd1 vssd1 vccd1 vccd1 _5348_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput185 _5483_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[13] sky130_fd_sc_hd__buf_2
Xoutput196 _5479_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[9] sky130_fd_sc_hd__buf_2
XFILLER_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5279_ _5736_/Q _5771_/A _5285_/S vssd1 vssd1 vccd1 vccd1 _5280_/B sky130_fd_sc_hd__mux2_1
XFILLER_233_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4517__A _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_285 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4787__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5615__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5067__B _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_266_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_238_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5022__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4778__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4242__A1 _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ _5390_/Q vssd1 vssd1 vccd1 vccd1 _2980_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4242__B2 _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5258__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4650_ _4642_/Y _4646_/X _4649_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5548_/D sky130_fd_sc_hd__o211a_1
Xinput10 i_mem_data[12] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_2
X_3601_ _3599_/B _3601_/B _3601_/C vssd1 vssd1 vccd1 vccd1 _3602_/A sky130_fd_sc_hd__and3b_4
Xinput21 i_mem_data[8] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 i_req_data[17] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5408__D _5408_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4581_ _5768_/A _4581_/B vssd1 vssd1 vccd1 vccd1 _4581_/X sky130_fd_sc_hd__or2_1
Xinput43 i_req_data[27] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
XFILLER_238_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput54 i_req_data[8] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
X_3532_ _3585_/B vssd1 vssd1 vccd1 vccd1 _3532_/X sky130_fd_sc_hd__buf_4
XFILLER_155_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3463_ _5412_/Q input46/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3464_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5202_ _5201_/X _5321_/A _5464_/Q vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4702__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_276_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3394_ _2845_/B _5377_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3395_/A sky130_fd_sc_hd__mux2_1
X_5133_ _5200_/B _5130_/Y _5155_/B _5132_/X vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__a31o_1
XFILLER_269_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5064_ _5231_/S vssd1 vssd1 vccd1 vccd1 _5200_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_270_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4015_ _4306_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _4015_/X sky130_fd_sc_hd__or2_1
XANTENNA__4481__A1 _5530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4056__B _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4233__A1 _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4917_ _5645_/Q _4947_/B vssd1 vssd1 vccd1 vccd1 _4917_/X sky130_fd_sc_hd__or2_1
XFILLER_240_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5168__A _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3992__A0 _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4848_ _5616_/Q _4856_/A vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__or2_1
XFILLER_165_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4779_ _5587_/Q _4781_/A vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__or2_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3744__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4800__A _5683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4395__S1 _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_216_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2786__A1 _5580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3983__A0 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2786__B2 _5660_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_316 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3735__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5721_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_258_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4215__A1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4215__B2 _4096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_222_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5751_ _5756_/CLK _5751_/D vssd1 vssd1 vccd1 vccd1 _5751_/Q sky130_fd_sc_hd__dfxtp_1
X_2963_ _5404_/Q vssd1 vssd1 vccd1 vccd1 _3084_/A sky130_fd_sc_hd__inv_2
XANTENNA__2777__A1 _5550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2777__B2 _2776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4702_ _5558_/Q _4697_/A _4701_/Y _4670_/X vssd1 vssd1 vccd1 vccd1 _5558_/D sky130_fd_sc_hd__o211a_1
XFILLER_147_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5682_ _5686_/CLK _5682_/D vssd1 vssd1 vccd1 vccd1 _5682_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3000__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2894_ _5364_/Q _5363_/Q _5362_/Q vssd1 vssd1 vccd1 vccd1 _3330_/C sky130_fd_sc_hd__nor3_4
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _5775_/A _4633_/B vssd1 vssd1 vccd1 vccd1 _4634_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4564_ _4561_/Y _4563_/X _4634_/A vssd1 vssd1 vccd1 vccd1 _4564_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3515_ _5437_/Q input43/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3516_/A sky130_fd_sc_hd__mux2_1
X_4495_ _4457_/Y _4493_/X _4492_/X _4491_/Y vssd1 vssd1 vccd1 vccd1 _4495_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_143_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3446_ _3446_/A vssd1 vssd1 vccd1 vccd1 _5402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4151__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _3376_/X _5370_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3378_/A sky130_fd_sc_hd__mux2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5460__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5116_ _5746_/Q _3840_/A _5115_/X vssd1 vssd1 vccd1 vccd1 _5116_/Y sky130_fd_sc_hd__a21oi_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4067__A _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5047_ _5047_/A vssd1 vssd1 vccd1 vccd1 _5703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_272_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4206__A1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4206__B2 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_378 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_138_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4509__A2 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3193__A1 _5669_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4390__B1 _4363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3791__D _3791_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4142__A0 _4140_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input24_A i_req_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4445__A1 _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__B2 _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4748__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4424__B _4424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2759__A1 _5552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5239__C _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5333__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3184__A1 _5603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3184__B2 _5619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4920__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3300_ _5366_/Q _3300_/B vssd1 vssd1 vccd1 vccd1 _3300_/X sky130_fd_sc_hd__or2_1
XFILLER_235_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5483__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4280_ _4080_/X _4280_/B vssd1 vssd1 vccd1 vccd1 _4281_/B sky130_fd_sc_hd__and2b_1
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2895__A _5361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3231_ _3419_/S vssd1 vssd1 vccd1 vccd1 _5406_/D sky130_fd_sc_hd__inv_2
XANTENNA__3490__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5271__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3162_ _5550_/Q _3131_/X _3159_/X _3161_/X vssd1 vssd1 vccd1 vccd1 _3162_/X sky130_fd_sc_hd__o22a_1
XFILLER_251_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__B_N _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3093_ _4682_/S vssd1 vssd1 vccd1 vccd1 _4651_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4436__A1 _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2834__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3995_ _5527_/Q _3923_/A _3994_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5527_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3947__A0 _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5734_ _5740_/CLK _5734_/D vssd1 vssd1 vccd1 vccd1 _5734_/Q sky130_fd_sc_hd__dfxtp_1
X_2946_ _2946_/A _3775_/B vssd1 vssd1 vccd1 vccd1 _3772_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5665_ _5665_/CLK _5665_/D vssd1 vssd1 vccd1 vccd1 _5665_/Q sky130_fd_sc_hd__dfxtp_2
X_2877_ _3308_/A vssd1 vssd1 vccd1 vccd1 _2877_/Y sky130_fd_sc_hd__inv_2
XFILLER_276_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4350__A _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4616_ _5772_/A _4581_/B _4612_/Y _4615_/Y _3919_/X vssd1 vssd1 vccd1 vccd1 _5544_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2789__B _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5596_ _5598_/CLK _5596_/D vssd1 vssd1 vccd1 vccd1 _5596_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_276_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3175__A1 _5649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3175__B2 _5569_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4911__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4547_ _4552_/B _4552_/C vssd1 vssd1 vccd1 vccd1 _4547_/X sky130_fd_sc_hd__or2_1
XFILLER_150_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4478_ _4484_/B _4484_/C _4478_/C vssd1 vssd1 vccd1 vccd1 _4482_/B sky130_fd_sc_hd__or3_4
XFILLER_277_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3429_ _5394_/Q _3038_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3430_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4427__A1 _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3132__C input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5356__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3938__A0 _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3575__S _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3166__A1 _5631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4902__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3307__C _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5312__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4666__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2677__B1 _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5030__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2881__C _3304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3641__A2 _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_20_i_clk clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5667_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_204_164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2800_ _2800_/A vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__clkbuf_4
X_3780_ _3780_/A _3780_/B vssd1 vssd1 vccd1 vccd1 _3780_/Y sky130_fd_sc_hd__nand2_1
X_2731_ _2731_/A vssd1 vssd1 vccd1 vccd1 _5311_/A sky130_fd_sc_hd__buf_4
XFILLER_145_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5450_ _5692_/CLK _5450_/D vssd1 vssd1 vccd1 vccd1 _5450_/Q sky130_fd_sc_hd__dfxtp_2
X_2662_ _2653_/X _2658_/X _2661_/X _2791_/B _5562_/Q vssd1 vssd1 vccd1 vccd1 _2663_/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_67_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3157__A1 _5549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4401_ _4491_/A _4401_/B _4600_/B _4490_/B vssd1 vssd1 vccd1 vccd1 _4401_/Y sky130_fd_sc_hd__nor4_1
X_5381_ _5722_/CLK _5381_/D vssd1 vssd1 vccd1 vccd1 _5381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4332_ _4332_/A _4332_/B _4332_/C _4332_/D vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__and4_1
XFILLER_125_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4263_ _3692_/X _4083_/B _4015_/X _4262_/X vssd1 vssd1 vccd1 vccd1 _4263_/X sky130_fd_sc_hd__a22o_1
XFILLER_86_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3214_ _5609_/Q _3133_/A _3135_/A _5625_/Q _3213_/X vssd1 vssd1 vccd1 vccd1 _3214_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_274_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4194_ _4194_/A _4194_/B vssd1 vssd1 vccd1 vccd1 _4213_/A sky130_fd_sc_hd__and2_1
XANTENNA__2775__D _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3145_ _3145_/A vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _3089_/A _3079_/B vssd1 vssd1 vccd1 vccd1 _3076_/Y sky130_fd_sc_hd__nor2_1
XFILLER_199_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5379__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4064__B _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3978_ _5523_/Q _3923_/A _3977_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5523_/D sky130_fd_sc_hd__o211a_1
X_5717_ _5757_/CLK _5717_/D vssd1 vssd1 vccd1 vccd1 _5717_/Q sky130_fd_sc_hd__dfxtp_1
X_2929_ _3307_/A _2946_/A vssd1 vssd1 vccd1 vccd1 _3317_/B sky130_fd_sc_hd__nand2_1
X_5648_ _5667_/CLK _5648_/D vssd1 vssd1 vccd1 vccd1 _5648_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4345__B1 _4340_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5579_ _5675_/CLK _5579_/D vssd1 vssd1 vccd1 vccd1 _5579_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4896__A1 _5636_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3699__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4239__B _4239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2685__D _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3320__A1 _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_250 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__A1 _5529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4255__A _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__A2 _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4179__A3 _4127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4584__A0 _5521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4336__B1 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4887__A1 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4639__A1 _5775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5521__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 i_mem_data[10] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_224_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4950_ _5687_/Q _4950_/B vssd1 vssd1 vccd1 vccd1 _4969_/A sky130_fd_sc_hd__and2_1
XFILLER_17_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3614__A2 _3572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4811__A1 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5671__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3901_ _3901_/A vssd1 vssd1 vccd1 vccd1 _5504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4881_ _5630_/Q _4910_/B vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__or2_1
XFILLER_232_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3832_ _5483_/Q _5387_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3833_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4575__A0 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3763_ _4528_/A vssd1 vssd1 vccd1 vccd1 _4585_/A sky130_fd_sc_hd__inv_2
XFILLER_257_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5502_ _5756_/CLK _5502_/D vssd1 vssd1 vccd1 vccd1 _5502_/Q sky130_fd_sc_hd__dfxtp_1
X_2714_ _2714_/A vssd1 vssd1 vccd1 vccd1 _5315_/A sky130_fd_sc_hd__buf_4
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _5452_/Q _3683_/A _3683_/X _5449_/Q _3693_/X vssd1 vssd1 vccd1 vccd1 _3694_/X
+ sky130_fd_sc_hd__a221o_1
X_5433_ _5441_/CLK _5433_/D vssd1 vssd1 vccd1 vccd1 _5433_/Q sky130_fd_sc_hd__dfxtp_1
X_2645_ _2747_/D _2682_/A _2761_/B _5611_/Q vssd1 vssd1 vccd1 vccd1 _2645_/X sky130_fd_sc_hd__and4b_1
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4878__A1 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5364_ _5716_/CLK _5364_/D vssd1 vssd1 vccd1 vccd1 _5364_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4315_ _4496_/A vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__inv_2
X_5295_ _5327_/B vssd1 vssd1 vccd1 vccd1 _5295_/X sky130_fd_sc_hd__buf_2
XFILLER_273_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4246_ _4347_/A _4471_/S _4220_/X _4245_/X vssd1 vssd1 vccd1 vccd1 _4537_/B sky130_fd_sc_hd__a31o_4
XFILLER_259_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4059__B _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4177_ _4373_/A _4177_/B vssd1 vssd1 vccd1 vccd1 _4177_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3128_ _3128_/A vssd1 vssd1 vccd1 vccd1 _3128_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ _5399_/Q _3060_/B vssd1 vssd1 vccd1 vccd1 _3069_/C sky130_fd_sc_hd__and2_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4566__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4522__B _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3138__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4869__A1 _5625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5151__A1_N _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5544__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5694__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5046__A1 _4482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3601__B _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__A0 _5680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4100_ _4194_/A _4194_/B _4213_/B _4099_/X vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__a211o_2
XFILLER_110_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5080_ _5705_/Q _5235_/S _5078_/X _5079_/Y vssd1 vssd1 vccd1 vccd1 _5705_/D sky130_fd_sc_hd__a22o_1
XFILLER_173_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5285__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3999__A _4045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _4067_/A _4232_/B vssd1 vssd1 vccd1 vccd1 _4031_/X sky130_fd_sc_hd__and2_1
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3296__B1 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5037__A1 _4600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4933_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__buf_6
XANTENNA__4260__A2 _4014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3938__S _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2842__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4864_ _4976_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4864_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5417__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3815_ _5242_/S vssd1 vssd1 vccd1 vccd1 _3834_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__4548__B1 _4529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4795_ _4983_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3746_ _4379_/C vssd1 vssd1 vccd1 vccd1 _4112_/B sky130_fd_sc_hd__clkinv_2
XFILLER_118_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3220__B1 _3149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5567__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3677_ _4030_/A _3751_/B vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__or2_2
XFILLER_133_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5416_ _5757_/CLK _5416_/D vssd1 vssd1 vccd1 vccd1 _5416_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput120 _5552_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[4] sky130_fd_sc_hd__buf_2
Xoutput131 _5700_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[11] sky130_fd_sc_hd__buf_2
Xoutput142 _5697_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[8] sky130_fd_sc_hd__buf_2
Xoutput153 _3104_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[3] sky130_fd_sc_hd__buf_2
XANTENNA__3523__A1 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3241__B_N _5473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5347_ _5692_/CLK _5347_/D vssd1 vssd1 vccd1 vccd1 _5347_/Q sky130_fd_sc_hd__dfxtp_4
Xoutput164 _3017_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_87_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput175 _3043_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[5] sky130_fd_sc_hd__buf_2
Xoutput186 _5484_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[14] sky130_fd_sc_hd__buf_2
Xoutput197 _5067_/B vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[0] sky130_fd_sc_hd__buf_2
X_5278_ _5278_/A vssd1 vssd1 vccd1 vccd1 _5735_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5276__A1 _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4229_ _4229_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _4229_/X sky130_fd_sc_hd__or2_1
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3702__A _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4517__B _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2740__A_N _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4236__C1 _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_253_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4787__B1 _4786_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4533__A _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4539__B1 _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3149__A _3149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3211__B1 _3145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3583__S _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input54_A i_req_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5267__A1 _5539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3278__B1 _3308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3612__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4475__C1 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output210_A _5311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3600_ _3600_/A vssd1 vssd1 vccd1 vccd1 _3600_/X sky130_fd_sc_hd__buf_6
Xinput11 i_mem_data[13] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_2
XFILLER_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 i_mem_data[9] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4580_ _4585_/A _4576_/X _4579_/X vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__a21bo_1
XFILLER_238_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput33 i_req_data[18] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
Xinput44 i_req_data[28] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
X_3531_ _5468_/Q vssd1 vssd1 vccd1 vccd1 _3585_/B sky130_fd_sc_hd__clkbuf_4
Xinput55 i_req_data[9] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5274__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3462_ _3462_/A vssd1 vssd1 vccd1 vccd1 _5411_/D sky130_fd_sc_hd__clkbuf_1
X_5201_ _5200_/B _5198_/Y _5225_/B _5200_/Y vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__a31o_1
XFILLER_130_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3393_ _3393_/A vssd1 vssd1 vccd1 vccd1 _5376_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5132_ _5132_/A _5156_/B vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__and2_1
XFILLER_69_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5063_ _5196_/A _5462_/Q vssd1 vssd1 vccd1 vccd1 _5231_/S sky130_fd_sc_hd__or2_2
XANTENNA__2837__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_270_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4014_ _4278_/A _4278_/B _4278_/C vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4481__A2 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_18_i_clk_A clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_252_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4233__A2 _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4916_ _4646_/X _4912_/Y _4915_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5644_/D sky130_fd_sc_hd__o211a_1
XFILLER_240_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5168__B _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4847_ _4663_/X _4836_/Y _4846_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5615_/D sky130_fd_sc_hd__o211a_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4778_ _4679_/X _4761_/Y _4777_/X _4769_/X vssd1 vssd1 vccd1 vccd1 _5586_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3744__A1 _5639_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3729_ _5636_/Q _3605_/A _3608_/X _5588_/Q vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4800__B _4950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4154__D1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2781__B_N _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5123__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3275__A3 _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_332 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_260_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3680__B1 _4076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5732__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2786__A2 _2635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3735__A1 _5622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3735__B2 _5606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3607__A _3607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5094__A _5515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5033__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3342__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3488__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5750_ _5756_/CLK _5750_/D vssd1 vssd1 vccd1 vccd1 _5750_/Q sky130_fd_sc_hd__dfxtp_1
X_2962_ _5405_/Q vssd1 vssd1 vccd1 vccd1 _2962_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4696__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2777__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4701_ _4722_/A _4974_/A vssd1 vssd1 vccd1 vccd1 _4701_/Y sky130_fd_sc_hd__nand2_1
XFILLER_249_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3974__A1 _5522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5681_ _5686_/CLK _5681_/D vssd1 vssd1 vccd1 vccd1 _5681_/Q sky130_fd_sc_hd__dfxtp_2
X_2893_ _5453_/Q vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__buf_4
XFILLER_249_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4632_ _5774_/A _4511_/X _3919_/A _4631_/X vssd1 vssd1 vccd1 vccd1 _5546_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4901__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4563_ _4635_/A _3956_/A _4562_/Y _5294_/A vssd1 vssd1 vccd1 vccd1 _4563_/X sky130_fd_sc_hd__a211o_1
XFILLER_162_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3514_ _3514_/A vssd1 vssd1 vccd1 vccd1 _5436_/D sky130_fd_sc_hd__clkbuf_1
X_4494_ _4491_/Y _4492_/X _4493_/X _4457_/Y vssd1 vssd1 vccd1 vccd1 _4494_/X sky130_fd_sc_hd__a211o_1
XFILLER_103_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3445_ _5402_/Q _3078_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3446_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3951__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4151__A1 _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5605__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ input27/X _5422_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3376_/X sky130_fd_sc_hd__mux2_1
XFILLER_257_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5517_/Q _3931_/A _5082_/B _5497_/Q _5053_/X vssd1 vssd1 vccd1 vccd1 _5115_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_281_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4348__A _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3252__A _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5046_ _5703_/Q _4482_/B _5135_/S vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5100__B1 _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5755__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3662__A0 _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4083__A _4083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2659__A_N _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4611__C1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5167__A0 _4503_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4390__A1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3193__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4390__B2 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4127__D1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3146__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4142__A1 _4141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4258__A _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_102_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_236_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4445__A2 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A i_mem_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4705__B _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3405__A0 _2845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2759__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4712__A1_N input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2940__S _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3708__A1 _5560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5028__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3337__A _5353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4381__A1 _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3184__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output85_A _3458_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5330__A0 _5329_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3230_ _3768_/S _3346_/B _3458_/C _3345_/A vssd1 vssd1 vccd1 vccd1 _3419_/S sky130_fd_sc_hd__o211ai_4
XANTENNA__2895__B _5360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3161_ _5630_/Q _3143_/X _3145_/X _3160_/X vssd1 vssd1 vccd1 vccd1 _3161_/X sky130_fd_sc_hd__a211o_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_251_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3092_ _5688_/Q _5677_/Q vssd1 vssd1 vccd1 vccd1 _4682_/S sky130_fd_sc_hd__nand2_4
XANTENNA__3644__B1 _3606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4841__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3994_ _3948_/B _3992_/X _3993_/Y _3965_/A vssd1 vssd1 vccd1 vccd1 _3994_/X sky130_fd_sc_hd__a211o_1
XFILLER_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _3795_/B _2945_/B vssd1 vssd1 vccd1 vccd1 _2951_/B sky130_fd_sc_hd__nor2_1
X_5733_ _5740_/CLK _5733_/D vssd1 vssd1 vccd1 vccd1 _5733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2876_ _3317_/A _2949_/B vssd1 vssd1 vccd1 vccd1 _3308_/A sky130_fd_sc_hd__nor2_2
XFILLER_30_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5664_ _5667_/CLK _5664_/D vssd1 vssd1 vccd1 vccd1 _5664_/Q sky130_fd_sc_hd__dfxtp_2
X_4615_ _4621_/B _4614_/Y _4581_/B vssd1 vssd1 vccd1 vccd1 _4615_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_276_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5595_ _5659_/CLK _5595_/D vssd1 vssd1 vccd1 vccd1 _5595_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2789__C _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3175__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4546_ _4552_/B _4552_/C vssd1 vssd1 vccd1 vccd1 _4546_/Y sky130_fd_sc_hd__nand2_1
XFILLER_209_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4477_ _5529_/Q _4458_/A _4476_/Y _3986_/X vssd1 vssd1 vccd1 vccd1 _5529_/D sky130_fd_sc_hd__o211a_1
XFILLER_277_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3428_ _3428_/A vssd1 vssd1 vccd1 vccd1 _5393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_277_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_225_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input9_A i_mem_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3883__A0 _5499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3359_ _3359_/A vssd1 vssd1 vccd1 vccd1 _5362_/D sky130_fd_sc_hd__clkbuf_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5029_ _5029_/A vssd1 vssd1 vccd1 vccd1 _5695_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__A _5598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2989__A2 _2852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5757_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_166_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3166__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3323__C1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2677__B2 _5560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3626__B1 _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output123_A _5555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5091__A2 _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4823__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_251_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3929__A1 _5512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2730_ _5555_/Q _2720_/B _2726_/X _2729_/X vssd1 vssd1 vccd1 vccd1 _2731_/A sky130_fd_sc_hd__o22a_1
XANTENNA__5450__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2661_ _5578_/Q _2644_/A _2686_/A _2659_/X _2660_/X vssd1 vssd1 vccd1 vccd1 _2661_/X
+ sky130_fd_sc_hd__a2111o_1
X_4400_ _4483_/A _4387_/Y _4389_/Y _4399_/X vssd1 vssd1 vccd1 vccd1 _4490_/B sky130_fd_sc_hd__a211o_4
XANTENNA__4354__A1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3157__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4354__B2 _3555_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5380_ _5722_/CLK _5380_/D vssd1 vssd1 vccd1 vccd1 _5380_/Q sky130_fd_sc_hd__dfxtp_1
X_4331_ _2954_/X _4069_/C _4330_/X vssd1 vssd1 vccd1 vccd1 _4332_/D sky130_fd_sc_hd__a21oi_1
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4262_ _5450_/Q _3617_/A _4011_/X _5445_/Q _5452_/Q vssd1 vssd1 vccd1 vccd1 _4262_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _5673_/Q _3137_/A _3139_/A _5593_/Q vssd1 vssd1 vccd1 vccd1 _3213_/X sky130_fd_sc_hd__a22o_1
X_4193_ _4350_/A _4191_/Y _4192_/X _4037_/A _2936_/X vssd1 vssd1 vccd1 vccd1 _4193_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3006__S _3346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ input3/X input2/X input1/X vssd1 vssd1 vccd1 vccd1 _3145_/A sky130_fd_sc_hd__nor3_4
XFILLER_267_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_282_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3075_ _5402_/Q _3075_/B vssd1 vssd1 vccd1 vccd1 _3079_/B sky130_fd_sc_hd__and2_1
XFILLER_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3530__A _4024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4290__B1 _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_332 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3977_ _3990_/A _3977_/B vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__or2_1
XFILLER_210_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5716_ _5716_/CLK _5716_/D vssd1 vssd1 vccd1 vccd1 _5716_/Q sky130_fd_sc_hd__dfxtp_1
X_2928_ _2928_/A _3284_/B vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__nor2_1
XFILLER_148_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5647_ _5747_/CLK _5647_/D vssd1 vssd1 vccd1 vccd1 _5647_/Q sky130_fd_sc_hd__dfxtp_2
X_2859_ _5354_/Q vssd1 vssd1 vccd1 vccd1 _3016_/A sky130_fd_sc_hd__inv_2
XANTENNA__4345__A1 _4171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4345__B2 _4341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5578_ _5674_/CLK _5578_/D vssd1 vssd1 vccd1 vccd1 _5578_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4896__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4529_ _4529_/A vssd1 vssd1 vccd1 vccd1 _4529_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4300__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_273_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4536__A _5515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4805__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5073__A2 _5051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4255__B _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5473__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4271__A _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3318__C _3318_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4887__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3615__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4639__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5297__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3311__A2 _3318_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 i_mem_data[11] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4272__A0 _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4811__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3900_ _5261_/A _3900_/B vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__and2_1
XFILLER_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4880_ _4653_/X _4874_/Y _4879_/X _4862_/X vssd1 vssd1 vccd1 vccd1 _5629_/D sky130_fd_sc_hd__o211a_1
XFILLER_177_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _3831_/A vssd1 vssd1 vccd1 vccd1 _5482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3496__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5277__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4575__A1 _5156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3762_ _5291_/S _3762_/B vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__nand2_1
X_5501_ _5756_/CLK _5501_/D vssd1 vssd1 vccd1 vccd1 _5501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2713_ _2705_/X _2706_/X _2711_/X _2712_/X vssd1 vssd1 vccd1 vccd1 _2714_/A sky130_fd_sc_hd__o31a_1
X_3693_ _5450_/Q _4447_/S _3572_/X _3692_/X vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__a22o_1
XFILLER_257_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4327__A1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5432_ _5441_/CLK _5432_/D vssd1 vssd1 vccd1 vccd1 _5432_/Q sky130_fd_sc_hd__dfxtp_1
X_2644_ _2644_/A vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__buf_6
XFILLER_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4878__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5363_ _5757_/CLK _5363_/D vssd1 vssd1 vccd1 vccd1 _5363_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3525__A _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4314_ _4294_/Y _4298_/X _4313_/Y _4093_/Y _4333_/A vssd1 vssd1 vccd1 vccd1 _4496_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_259_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5294_ _5294_/A _5294_/B vssd1 vssd1 vccd1 vccd1 _5327_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5346__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4245_ _4355_/A _4225_/Y _4236_/X _4238_/Y _4244_/Y vssd1 vssd1 vccd1 vccd1 _4245_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_113_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4176_ _4466_/A _4059_/B _4373_/A vssd1 vssd1 vccd1 vccd1 _4176_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3127_ _5711_/Q _5719_/Q _4651_/S vssd1 vssd1 vccd1 vccd1 _3128_/A sky130_fd_sc_hd__mux2_1
XFILLER_215_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5496__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3058_ _3343_/C _3056_/X _3057_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3058_/X sky130_fd_sc_hd__o211a_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4566__A1 _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4318__A1 _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4869__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3601__C _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__A1 _5681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4713__B _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4557__A1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_329 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output190_A _5473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5369__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_284_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4030_ _4030_/A _4063_/A vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__and2_1
XFILLER_256_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4493__B1 _4457_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3048__A1 _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4932_ _4970_/A _4935_/B vssd1 vssd1 vccd1 vccd1 _4932_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4796__A1 _5594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3453__D1 _3346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4863_ _5622_/Q _4859_/B _4861_/Y _4862_/X vssd1 vssd1 vccd1 vccd1 _5622_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4548__A1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _3814_/A vssd1 vssd1 vccd1 vccd1 _5474_/D sky130_fd_sc_hd__clkbuf_1
X_4794_ _5593_/Q _4784_/B _4793_/Y _4791_/X vssd1 vssd1 vccd1 vccd1 _5593_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3745_ _5559_/Q _3596_/X _3742_/X _3744_/X vssd1 vssd1 vccd1 vccd1 _4379_/C sky130_fd_sc_hd__o22a_4
XANTENNA__3220__A1 _5658_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3220__B2 _5578_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3676_ _4466_/A _5444_/Q vssd1 vssd1 vccd1 vccd1 _3751_/B sky130_fd_sc_hd__nor2_2
XFILLER_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_14_i_clk_A clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5415_ _5757_/CLK _5415_/D vssd1 vssd1 vccd1 vccd1 _5415_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput110 _5548_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[0] sky130_fd_sc_hd__buf_2
Xoutput121 _5553_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[5] sky130_fd_sc_hd__buf_2
Xoutput132 _5701_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[12] sky130_fd_sc_hd__buf_2
Xoutput143 _5698_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[9] sky130_fd_sc_hd__buf_2
Xoutput154 _3106_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[4] sky130_fd_sc_hd__buf_2
XFILLER_217_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _5738_/CLK _5346_/D vssd1 vssd1 vccd1 vccd1 _5346_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput165 _3068_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[10] sky130_fd_sc_hd__buf_2
Xoutput176 _3048_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[6] sky130_fd_sc_hd__buf_2
Xoutput187 _5485_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[15] sky130_fd_sc_hd__buf_2
XFILLER_87_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput198 _5317_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[10] sky130_fd_sc_hd__buf_2
X_5277_ _5292_/A _5277_/B vssd1 vssd1 vccd1 vccd1 _5278_/A sky130_fd_sc_hd__and2_1
XFILLER_247_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4228_ _4303_/A _4228_/B vssd1 vssd1 vccd1 vccd1 _4229_/B sky130_fd_sc_hd__nand2_1
XFILLER_247_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4159_ _4468_/A _4138_/Y _4147_/X _4158_/Y _4372_/B vssd1 vssd1 vccd1 vccd1 _4159_/X
+ sky130_fd_sc_hd__a311o_2
XFILLER_228_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_255_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4787__A1 _5590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4814__A _5602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3995__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4533__B _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4539__A1 _4536_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3211__A1 _5640_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5511__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5661__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input47_A i_req_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3278__A1 _3307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4475__B1 _4289_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3612__B _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4227__A0 _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4778__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output203_A _2650_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4724__A _5681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3202__A1 _5558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 i_mem_data[14] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
Xinput23 i_mem_exception vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__buf_4
Xinput34 i_req_data[19] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 i_req_data[29] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_3530_ _4024_/A vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__buf_6
Xinput56 i_req_data_valid vssd1 vssd1 vccd1 vccd1 _3346_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__2898__B _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3461_ _5411_/Q input35/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3462_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _5200_/A _5200_/B vssd1 vssd1 vccd1 vccd1 _5200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4702__A1 _5558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3392_ _2850_/B _5376_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3393_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _5131_/A _5131_/B _5131_/C vssd1 vssd1 vccd1 vccd1 _5155_/B sky130_fd_sc_hd__or3_2
XFILLER_257_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5062_ _5071_/B _5062_/B vssd1 vssd1 vccd1 vccd1 _5062_/Y sky130_fd_sc_hd__nand2_1
XFILLER_284_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4013_ _4274_/A _4281_/A vssd1 vssd1 vccd1 vccd1 _4278_/C sky130_fd_sc_hd__xnor2_1
XFILLER_203_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3674__D1 _3683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_252_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4634__A _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4915_ _5644_/Q _4947_/B vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__or2_1
XFILLER_240_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _5615_/Q _4872_/B vssd1 vssd1 vccd1 vccd1 _4846_/X sky130_fd_sc_hd__or2_1
XFILLER_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5194__B2 _5504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _5586_/Q _4781_/A vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__or2_1
XANTENNA__3744__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3728_ _5572_/Q _3607_/X _3598_/A _5604_/Q vssd1 vssd1 vccd1 vccd1 _3728_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5684__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2952__A0 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3659_ _5631_/Q _3605_/A _3606_/A _3658_/X vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__a211o_1
XFILLER_161_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5329_ _5329_/A vssd1 vssd1 vccd1 vccd1 _5329_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5185__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3196__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3735__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4696__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5407__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4448__B1 _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4438__B _4438_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_240_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5557__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4454__A _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2961_ _5444_/Q _3780_/A _2960_/X vssd1 vssd1 vccd1 vccd1 _5444_/D sky130_fd_sc_hd__o21ba_1
XFILLER_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ input8/X _4689_/X _4690_/X _4699_/Y vssd1 vssd1 vccd1 vccd1 _4974_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_187_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5680_ _5680_/CLK _5680_/D vssd1 vssd1 vccd1 vccd1 _5680_/Q sky130_fd_sc_hd__dfxtp_2
X_2892_ _2892_/A vssd1 vssd1 vccd1 vccd1 _5454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4631_ _4585_/A _4627_/X _4630_/Y _4529_/X vssd1 vssd1 vccd1 vccd1 _4631_/X sky130_fd_sc_hd__a211o_1
XFILLER_187_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4901__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _4635_/A _5132_/A vssd1 vssd1 vccd1 vccd1 _4562_/Y sky130_fd_sc_hd__nor2_1
X_3513_ _5436_/Q input42/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3514_/A sky130_fd_sc_hd__mux2_1
X_4493_ _4484_/B _4484_/C _4478_/C _4457_/D vssd1 vssd1 vccd1 vccd1 _4493_/X sky130_fd_sc_hd__o31a_1
XFILLER_265_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3444_ _3444_/A vssd1 vssd1 vccd1 vccd1 _5401_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2848__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4151__A2 _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3375_ _3375_/A vssd1 vssd1 vccd1 vccd1 _5369_/D sky130_fd_sc_hd__clkbuf_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3533__A _5472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5517_/Q vssd1 vssd1 vccd1 vccd1 _5114_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_257_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3252__B _3252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5100__A1 _4536_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5045_ _5045_/A vssd1 vssd1 vccd1 vccd1 _5702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_150_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3662__A1 _4024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4083__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4829_ _5608_/Q _4822_/B _4828_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5608_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3178__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4390__A2 _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5345__D _5345_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3146__C input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4678__A0 _5710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5134__S _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3350__A0 _2826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_124_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_105 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3653__A1 _5566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3653__B2 _5582_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4274__A _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4602__B1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2835__D_N _2826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5158__A1 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3169__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3708__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3337__B _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output78_A _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5330__A1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5044__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3160_ _5646_/Q _3147_/X _3149_/X _5566_/Q vssd1 vssd1 vccd1 vccd1 _3160_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3892__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3091_ _5775_/A _3010_/X _3090_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3091_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3644__A1 _5666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3499__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_196 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3993_ _4635_/B _3993_/B vssd1 vssd1 vccd1 vccd1 _3993_/Y sky130_fd_sc_hd__nor2_1
X_5732_ _5740_/CLK _5732_/D vssd1 vssd1 vccd1 vccd1 _5732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_328 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2944_ _2938_/B _3284_/B _5241_/C vssd1 vssd1 vccd1 vccd1 _3791_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__4912__A _5686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5149__A1 _5520_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5663_ _5747_/CLK _5663_/D vssd1 vssd1 vccd1 vccd1 _5663_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5149__B2 _5500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2875_ _5360_/Q _5361_/Q vssd1 vssd1 vccd1 vccd1 _2949_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__3528__A _3528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4614_ _5772_/A _4605_/A _4634_/A vssd1 vssd1 vccd1 vccd1 _4614_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_190_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5594_ _5675_/CLK _5594_/D vssd1 vssd1 vccd1 vccd1 _5594_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2789__D _5596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3247__B _3843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4545_ _4542_/Y _4544_/X _4532_/X vssd1 vssd1 vccd1 vccd1 _4545_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4476_ _3935_/A _4485_/A _4458_/A _4475_/X vssd1 vssd1 vccd1 vccd1 _4476_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_145_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3427_ _5393_/Q _3034_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3428_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5722__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3004_/B _5362_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3359_/A sky130_fd_sc_hd__mux2_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3883__A1 _5311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _5367_/Q _3297_/B vssd1 vssd1 vccd1 vccd1 _3300_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5085__B1 _5460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5028_ _5695_/Q _4361_/A _5030_/S vssd1 vssd1 vccd1 vccd1 _5029_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4806__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_54_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_241_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3399__A0 _2840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4822__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3323__B1 _3335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_282_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5076__B1 _4514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3087__C1 _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3626__B2 _5553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output116_A _5563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_368 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2733_/A _2747_/B _5658_/Q _2747_/D vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__and4b_1
XFILLER_172_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4354__A2 _4203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5745__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ _2904_/X _4028_/X _4033_/X _5445_/Q _4329_/X vssd1 vssd1 vccd1 vccd1 _4330_/X
+ sky130_fd_sc_hd__a221o_1
X_4261_ _4259_/Y _4260_/Y _4081_/Y vssd1 vssd1 vccd1 vccd1 _4261_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_140_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_219 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3212_ _5560_/Q _3131_/A _3209_/X _3211_/X vssd1 vssd1 vccd1 vccd1 _3212_/X sky130_fd_sc_hd__o22a_2
XFILLER_262_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4192_ _4192_/A _4192_/B _4192_/C vssd1 vssd1 vccd1 vccd1 _4192_/X sky130_fd_sc_hd__or3_1
XFILLER_274_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3143_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3143_/X sky130_fd_sc_hd__buf_4
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4907__A _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3074_ _5402_/Q _3075_/B vssd1 vssd1 vccd1 vccd1 _3074_/X sky130_fd_sc_hd__or2_1
XANTENNA__3078__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4642__A _5680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3976_ _3975_/X _5319_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3977_/B sky130_fd_sc_hd__mux2_1
XFILLER_210_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5715_ _5716_/CLK _5715_/D vssd1 vssd1 vccd1 vccd1 _5715_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4361__B _5132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2927_ _2946_/A _3775_/B _3330_/C _5241_/A vssd1 vssd1 vccd1 vccd1 _3791_/B sky130_fd_sc_hd__a31o_1
XFILLER_148_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5646_ _5653_/CLK _5646_/D vssd1 vssd1 vccd1 vccd1 _5646_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2858_ _2830_/Y _2853_/Y _3004_/B _2857_/Y vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4345__A2 _4339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3002__C1 _3001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5577_ _5675_/CLK _5577_/D vssd1 vssd1 vccd1 vccd1 _5577_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_163_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2789_ _2774_/C _2789_/B _2789_/C _5596_/Q vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__and4b_1
X_4528_ _4528_/A _4528_/B _4528_/C vssd1 vssd1 vccd1 vccd1 _4528_/X sky130_fd_sc_hd__and3_1
XANTENNA__4750__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_37 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4459_ _5067_/B _4289_/C _4401_/Y _4457_/Y _4458_/Y vssd1 vssd1 vccd1 vccd1 _4459_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2667__B_N _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4817__A _5603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_364 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2816__C1 _5353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__A _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4271__B _4271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3792__B1 _3791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4336__A2 _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4727__A _5564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__B1 _5460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4272__A1 _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3777__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3830_ _5482_/Q _5386_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3831_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5221__A0 _4457_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3761_ _3761_/A _3267_/B vssd1 vssd1 vccd1 vccd1 _3762_/B sky130_fd_sc_hd__or2b_1
X_5500_ _5740_/CLK _5500_/D vssd1 vssd1 vccd1 vccd1 _5500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2712_ _5557_/Q _2720_/B vssd1 vssd1 vccd1 vccd1 _2712_/X sky130_fd_sc_hd__or2_1
XFILLER_72_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4980__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3692_ _5446_/Q _4160_/A vssd1 vssd1 vccd1 vccd1 _3692_/X sky130_fd_sc_hd__or2_2
XFILLER_257_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5431_ _5441_/CLK _5431_/D vssd1 vssd1 vccd1 vccd1 _5431_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4327__A2 _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2643_ _2681_/A _2761_/B _5346_/Q vssd1 vssd1 vccd1 vccd1 _2644_/A sky130_fd_sc_hd__nor3b_1
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5362_ _5716_/CLK _5362_/D vssd1 vssd1 vccd1 vccd1 _5362_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4732__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4313_ _4347_/A _4428_/B _4305_/Y _4309_/X _4312_/X vssd1 vssd1 vccd1 vccd1 _4313_/Y
+ sky130_fd_sc_hd__a221oi_2
XANTENNA__3525__B _5331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5293_ _5293_/A vssd1 vssd1 vccd1 vccd1 _5740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_273_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5716_/CLK sky130_fd_sc_hd__clkbuf_16
X_4244_ _4171_/A _4240_/X _4243_/Y vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_259_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2856__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4175_ _4468_/A _4175_/B vssd1 vssd1 vccd1 vccd1 _4175_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3541__A _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_255_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_10_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3057_ _5768_/A _3063_/B vssd1 vssd1 vccd1 vccd1 _3057_/X sky130_fd_sc_hd__or2_1
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_230_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5187__B _5187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4566__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3959_ _5539_/Q _5732_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3959_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4971__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_224 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_176_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5629_ _5653_/CLK _5629_/D vssd1 vssd1 vccd1 vccd1 _5629_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_191_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3526__B1 _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4723__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4547__A _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5440__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__A1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_194 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4962__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output183_A _5481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4714__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output60_A _3207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_264_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4245__A1 _4355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4931_ _4931_/A vssd1 vssd1 vccd1 vccd1 _4935_/B sky130_fd_sc_hd__buf_4
XFILLER_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4796__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3453__C1 _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4862_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__buf_4
XFILLER_268_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3813_ _5474_/Q _5378_/Q _3813_/S vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__mux2_1
XFILLER_268_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4793_ _4981_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4793_/Y sky130_fd_sc_hd__nand2_1
X_3744_ _5639_/Q _3605_/X _3606_/X _3743_/X vssd1 vssd1 vccd1 vccd1 _3744_/X sky130_fd_sc_hd__a211o_1
XFILLER_158_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4953__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3220__A2 _3147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3675_ _4454_/B _4303_/A _3662_/X _3674_/X _3617_/A vssd1 vssd1 vccd1 vccd1 _3675_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_137_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3536__A _5471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5414_ _5757_/CLK _5414_/D vssd1 vssd1 vccd1 vccd1 _5414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput100 _5775_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[15] sky130_fd_sc_hd__buf_2
Xoutput111 _5558_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[10] sky130_fd_sc_hd__buf_2
XFILLER_279_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput122 _5554_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[6] sky130_fd_sc_hd__buf_2
Xoutput133 _5702_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput144 _3098_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[0] sky130_fd_sc_hd__buf_2
X_5345_ _5738_/CLK _5345_/D vssd1 vssd1 vccd1 vccd1 _5345_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput155 _3108_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[5] sky130_fd_sc_hd__buf_2
Xoutput166 _3073_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[11] sky130_fd_sc_hd__buf_2
Xoutput177 _3052_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[7] sky130_fd_sc_hd__buf_2
Xoutput188 _5471_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[1] sky130_fd_sc_hd__buf_2
XANTENNA__5463__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput199 _5319_/A vssd1 vssd1 vccd1 vccd1 sr_bus_data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5276_ _5735_/Q _5770_/A _5285_/S vssd1 vssd1 vccd1 vccd1 _5277_/B sky130_fd_sc_hd__mux2_1
X_4227_ _4132_/B _4161_/B _4302_/S vssd1 vssd1 vccd1 vccd1 _4228_/B sky130_fd_sc_hd__mux2_1
X_4158_ _4347_/B _4347_/C _4372_/A vssd1 vssd1 vccd1 vccd1 _4158_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_262_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3109_ _5710_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3110_/A sky130_fd_sc_hd__and2_1
XFILLER_228_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4089_ _4089_/A _4352_/A vssd1 vssd1 vccd1 vccd1 _4090_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4236__A1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4814__B _4819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4787__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5198__A _5198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4533__C _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4944__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4830__A _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3211__A2 _3143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3142__A_N input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_219_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4227__A1 _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4778__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4724__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4443__C _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5336__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 i_mem_data[15] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_2
XANTENNA__3202__A2 _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 i_req_data[0] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
Xinput35 i_req_data[1] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 i_req_data[2] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput57 i_rst vssd1 vssd1 vccd1 vccd1 _5300_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_182_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3460_ _3460_/A vssd1 vssd1 vccd1 vccd1 _5410_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5486__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3391_ _3391_/A vssd1 vssd1 vccd1 vccd1 _5375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_184_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5130_ _5131_/A _5131_/B _5131_/C vssd1 vssd1 vccd1 vccd1 _5130_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3910__B1 _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5061_ _5050_/X _5058_/X _3759_/X vssd1 vssd1 vccd1 vccd1 _5062_/B sky130_fd_sc_hd__o21ai_1
XFILLER_96_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4012_ _4229_/A _4281_/A vssd1 vssd1 vccd1 vccd1 _4012_/X sky130_fd_sc_hd__and2_1
XANTENNA__3674__C1 _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4218__A1 _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4915__A _5644_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3241__D _5471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4914_ _4931_/A vssd1 vssd1 vccd1 vccd1 _4947_/B sky130_fd_sc_hd__buf_4
XFILLER_279_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4845_ _4658_/X _4836_/Y _4844_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5614_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3729__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4926__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4776_ _4674_/X _4761_/Y _4775_/X _4769_/X vssd1 vssd1 vccd1 vccd1 _5585_/D sky130_fd_sc_hd__o211a_1
X_3727_ _5668_/Q _3600_/X _3602_/X _5652_/Q vssd1 vssd1 vccd1 vccd1 _3727_/X sky130_fd_sc_hd__a22o_1
X_3658_ _5567_/Q _3607_/A _3608_/A _5583_/Q vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__a22o_1
XFILLER_228_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4154__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3589_ _4124_/A _4045_/A _3619_/B _4379_/B vssd1 vssd1 vccd1 vccd1 _3590_/D sky130_fd_sc_hd__a211o_1
XFILLER_161_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5328_ _2650_/Y _5319_/B _5327_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5756_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_275_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5259_ _5259_/A vssd1 vssd1 vccd1 vccd1 _5729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_228_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3680__A2 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5359__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4560__A _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3196__A1 _5637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4448__A1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3115__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4735__A _5568_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5330__S _5720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4454__B _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3959__A0 _5539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2960_ _2877_/Y _2889_/B _2923_/B _3799_/A _3337_/B vssd1 vssd1 vccd1 vccd1 _2960_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4620__A1 _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _4466_/A _3283_/A _3337_/B vssd1 vssd1 vccd1 vccd1 _2892_/A sky130_fd_sc_hd__mux2_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4630_ _5253_/S _3762_/B _4629_/B _4629_/A _4633_/B vssd1 vssd1 vccd1 vccd1 _4630_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_8_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3187__A1 _5555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4561_ _5518_/Q _4599_/B vssd1 vssd1 vccd1 vccd1 _4561_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_162_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3512_ _3512_/A vssd1 vssd1 vccd1 vccd1 _5435_/D sky130_fd_sc_hd__clkbuf_1
X_4492_ _4491_/A _4491_/B _4491_/C vssd1 vssd1 vccd1 vccd1 _4492_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3443_ _5401_/Q _3073_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3444_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3373_/X _5369_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3375_/A sky130_fd_sc_hd__mux2_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5708_/Q _5235_/S _5111_/X _5112_/Y vssd1 vssd1 vccd1 vccd1 _5708_/D sky130_fd_sc_hd__a22o_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5702_/Q _4457_/D _5135_/S vssd1 vssd1 vccd1 vccd1 _5045_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5501__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_225_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4611__A1 _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5651__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _4978_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4828_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3178__A1 _5666_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3178__B2 _5586_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4759_ _4985_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4127__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5324__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3350__A1 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3653__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4274__B _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2803__A _5720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3169__A1 _5600_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3877__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5524__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3090_ _2850_/C _3027_/X _3018_/A _3089_/Y vssd1 vssd1 vccd1 vccd1 _3090_/X sky130_fd_sc_hd__a211o_1
XFILLER_181_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5164__A1_N _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3644__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4841__A1 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5674__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3992_ _5775_/A _5740_/Q _5329_/A vssd1 vssd1 vccd1 vccd1 _3992_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5731_ _5740_/CLK _5731_/D vssd1 vssd1 vccd1 vccd1 _5731_/Q sky130_fd_sc_hd__dfxtp_1
X_2943_ _3799_/A _2946_/A _2943_/C vssd1 vssd1 vccd1 vccd1 _5241_/C sky130_fd_sc_hd__and3b_1
XFILLER_200_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4912__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5662_ _5667_/CLK _5662_/D vssd1 vssd1 vccd1 vccd1 _5662_/Q sky130_fd_sc_hd__dfxtp_4
X_2874_ _5364_/Q _5363_/Q _5362_/Q vssd1 vssd1 vccd1 vccd1 _3317_/A sky130_fd_sc_hd__or3b_4
XFILLER_175_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4613_ _5772_/A _5771_/A _4613_/C vssd1 vssd1 vccd1 vccd1 _4621_/B sky130_fd_sc_hd__and3_1
X_5593_ _5659_/CLK _5593_/D vssd1 vssd1 vccd1 vccd1 _5593_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4544_ _4600_/A _3948_/A _4543_/Y _5294_/A vssd1 vssd1 vccd1 vccd1 _4544_/X sky130_fd_sc_hd__a211o_1
XFILLER_128_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5306__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4475_ _4462_/X _4465_/Y _4474_/X _4289_/C _4333_/A vssd1 vssd1 vccd1 vccd1 _4475_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_143_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5235__S _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3544__A _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3426_ _3426_/A vssd1 vssd1 vccd1 vccd1 _5392_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5117__A1_N _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3357_/A vssd1 vssd1 vccd1 vccd1 _5361_/D sky130_fd_sc_hd__clkbuf_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _3791_/A _3292_/D vssd1 vssd1 vccd1 vccd1 _3297_/B sky130_fd_sc_hd__nor2_1
X_5027_ _5027_/A vssd1 vssd1 vccd1 vccd1 _5694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_245_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4375__A _4396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_364 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4596__B1 _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4822__B _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_221_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5547__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3454__A _3523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4269__B _4269_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5697__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input22_A i_mem_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4823__A1 _5605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2834__A0 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4339__A0 _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4260_ _4012_/X _4014_/X _4350_/A vssd1 vssd1 vccd1 vccd1 _4260_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3314__A1 _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3211_ _5640_/Q _3143_/A _3145_/A _3210_/X vssd1 vssd1 vccd1 vccd1 _3211_/X sky130_fd_sc_hd__a211o_1
XFILLER_262_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4191_ _4192_/A _4192_/B _4192_/C vssd1 vssd1 vccd1 vccd1 _4191_/Y sky130_fd_sc_hd__o21ai_1
X_3142_ input2/X input1/X input3/X vssd1 vssd1 vccd1 vccd1 _3143_/A sky130_fd_sc_hd__and3b_4
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4907__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2708__A _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3073_ _5771_/A _3063_/B _3071_/Y _3072_/X _3016_/A vssd1 vssd1 vccd1 vccd1 _3073_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_227_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4923__A _5648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4578__B1 _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4642__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3975_ _5771_/A _5736_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3975_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2926_ _5359_/Q _3277_/A _3775_/A _3775_/C vssd1 vssd1 vccd1 vccd1 _5241_/A sky130_fd_sc_hd__and4_1
X_5714_ _5716_/CLK _5714_/D vssd1 vssd1 vccd1 vccd1 _5714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4361__C _4543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5645_ _5653_/CLK _5645_/D vssd1 vssd1 vccd1 vccd1 _5645_/Q sky130_fd_sc_hd__dfxtp_4
X_2857_ _3003_/A _3003_/B vssd1 vssd1 vccd1 vccd1 _2857_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3002__B1 _2830_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5576_ _5675_/CLK _5576_/D vssd1 vssd1 vccd1 vccd1 _5576_/Q sky130_fd_sc_hd__dfxtp_2
X_2788_ _2774_/C _2789_/C _2789_/B _5564_/Q vssd1 vssd1 vccd1 vccd1 _2788_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__3553__A1 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4527_ _5081_/A _4533_/C _4527_/C vssd1 vssd1 vccd1 vccd1 _4528_/C sky130_fd_sc_hd__nand3_1
XFILLER_116_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4458_ _4458_/A vssd1 vssd1 vccd1 vccd1 _4458_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3305__A1 _3330_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_155 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3409_ _2966_/A _5384_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3410_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4389_ _4389_/A _4389_/B vssd1 vssd1 vccd1 vccd1 _4389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4817__B _4819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5058__A1 _5051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_218_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4805__A1 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4708__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__B _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3883__S _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5297__A1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4727__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3123__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2807__A0 _5684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5712__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3760_ _4619_/B _3757_/X _3759_/X vssd1 vssd1 vccd1 vccd1 _3760_/Y sky130_fd_sc_hd__o21ai_1
X_2711_ _5621_/Q _2652_/X _2709_/X _2710_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2711_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3691_ _3691_/A _3691_/B vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__nor2_2
XANTENNA__3793__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5430_ _5441_/CLK _5430_/D vssd1 vssd1 vccd1 vccd1 _5430_/Q sky130_fd_sc_hd__dfxtp_1
X_2642_ _5595_/Q _2635_/Y _2636_/X _2638_/X _2641_/X vssd1 vssd1 vccd1 vccd1 _2642_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_65_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5361_ _5724_/CLK _5361_/D vssd1 vssd1 vccd1 vccd1 _5361_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_160_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2710__B _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3094__A _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4312_ _2954_/X _4071_/C _4310_/X _4311_/X vssd1 vssd1 vccd1 vccd1 _4312_/X sky130_fd_sc_hd__a211o_1
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _5292_/A _5292_/B vssd1 vssd1 vccd1 vccd1 _5293_/A sky130_fd_sc_hd__and2_1
XFILLER_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5288__A1 _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4243_ _4084_/B _4241_/X _4242_/X vssd1 vssd1 vccd1 vccd1 _4243_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3299__B1 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4174_ _4454_/A _4124_/B _4248_/C _4471_/S _4173_/X vssd1 vssd1 vccd1 vccd1 _4175_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3541__B _4301_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _5710_/Q _5718_/Q _4651_/S vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__mux2_1
XFILLER_255_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3056_ _3055_/Y _2845_/C _3089_/A vssd1 vssd1 vccd1 vccd1 _3056_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3968__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4263__A2 _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_270_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4372__B _4372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5392__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3269__A _5472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3223__B1 _3139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3958_ _5518_/Q _3923_/X _3957_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5518_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2909_ _3281_/B vssd1 vssd1 vccd1 vccd1 _3775_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_176_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3889_ _5501_/Q _5315_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3890_/B sky130_fd_sc_hd__mux2_1
XFILLER_176_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5628_ _5650_/CLK _5628_/D vssd1 vssd1 vccd1 vccd1 _5628_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3526__A1 _5347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5559_ _5675_/CLK _5559_/D vssd1 vssd1 vccd1 vccd1 _5559_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_191_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5279__A1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4828__A _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3878__S _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4254__A2 _4251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5735__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2804__A3 _5683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5203__A1 _5202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3214__B1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2789__A_N _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_326 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_110_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3788__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_252_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4930_ _4684_/X _4912_/Y _4929_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5651_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4650__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4861_ _4974_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4861_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3089__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3812_ _3812_/A vssd1 vssd1 vccd1 vccd1 _5473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3205__B1 _3149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4792_ _5592_/Q _4784_/B _4790_/Y _4791_/X vssd1 vssd1 vccd1 vccd1 _5592_/D sky130_fd_sc_hd__o211a_1
XFILLER_268_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3743_ _5575_/Q _3607_/X _3608_/X _5591_/Q vssd1 vssd1 vccd1 vccd1 _3743_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3239__D _5470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3674_ _4449_/S _4281_/A _4303_/A _4304_/S _3683_/A vssd1 vssd1 vccd1 vccd1 _3674_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_284_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5413_ _5757_/CLK _5413_/D vssd1 vssd1 vccd1 vccd1 _5413_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput101 _5761_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[1] sky130_fd_sc_hd__buf_2
XFILLER_173_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput112 _5559_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[11] sky130_fd_sc_hd__buf_2
XFILLER_217_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput123 _5555_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[7] sky130_fd_sc_hd__buf_2
XANTENNA__4181__A1 _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 _5703_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[14] sky130_fd_sc_hd__buf_2
X_5344_ _5738_/CLK _5344_/D vssd1 vssd1 vccd1 vccd1 _5344_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput145 _3118_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[10] sky130_fd_sc_hd__buf_2
XANTENNA__5608__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput156 _3110_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[6] sky130_fd_sc_hd__buf_2
Xoutput167 _3078_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[12] sky130_fd_sc_hd__buf_2
Xoutput178 _3058_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[8] sky130_fd_sc_hd__buf_2
Xoutput189 _5472_/Q vssd1 vssd1 vccd1 vccd1 sr_bus_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_141_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5275_ _5275_/A vssd1 vssd1 vccd1 vccd1 _5734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_275_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _3726_/Y _3740_/X _4272_/S vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5130__B1 _5131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4157_ _4469_/D _4198_/C _4396_/A vssd1 vssd1 vccd1 vccd1 _4347_/C sky130_fd_sc_hd__a21o_1
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _3108_/A vssd1 vssd1 vccd1 vccd1 _3108_/X sky130_fd_sc_hd__clkbuf_1
X_4088_ _4348_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__xor2_1
XFILLER_270_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3039_ _5395_/Q _5394_/Q _3039_/C vssd1 vssd1 vccd1 vccd1 _3045_/B sky130_fd_sc_hd__and3_1
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3995__A1 _5527_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4533__D _5760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4830__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2955__C1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4558__A _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5121__B1 _4499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4880__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_234_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2806__A _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3401__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A0 _4600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3738__A1 _5558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput14 i_mem_data[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
Xinput25 i_req_data[10] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 i_req_data[20] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
Xinput47 i_req_data[30] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4148__D1 _4128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2961__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4163__A1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4163__B2 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3390_ _2840_/A _5375_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3391_/A sky130_fd_sc_hd__mux2_1
XFILLER_254_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_254 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5112__B1 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5060_ _5156_/B _5060_/B vssd1 vssd1 vccd1 vccd1 _5060_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4011_ _4306_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _4011_/X sky130_fd_sc_hd__and2_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3674__B1 _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4871__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4218__A2 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4915__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ _5686_/Q _4950_/B vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__and2_4
XFILLER_178_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4931__A _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4844_ _5614_/Q _4872_/B vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__or2_1
XANTENNA__3729__A1 _5636_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3729__B2 _5588_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4775_ _5585_/Q _4781_/A vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__or2_1
XANTENNA__3547__A _5475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4142__S _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3726_ _3732_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5430__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3657_ _5663_/Q _3600_/A _3602_/A _5647_/Q _3656_/X vssd1 vssd1 vccd1 vccd1 _3657_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5762__A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4154__A1 _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3588_ _5481_/Q _5319_/A _3588_/S vssd1 vssd1 vccd1 vccd1 _4379_/B sky130_fd_sc_hd__mux2_8
XFILLER_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5580__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5327_ _5756_/Q _5327_/B vssd1 vssd1 vccd1 vccd1 _5327_/X sky130_fd_sc_hd__or2_1
XFILLER_275_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4097__B _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ _5261_/A _5258_/B vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__and2_1
X_4209_ _4503_/A vssd1 vssd1 vccd1 vccd1 _4362_/A sky130_fd_sc_hd__clkinv_2
XFILLER_275_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5189_ _5188_/X _5319_/A _5464_/Q vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3665__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4317__S _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3417__A0 _2850_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3968__A1 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4393__A1 _3678_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3196__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_137_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_1_0_i_clk clkbuf_2_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_i_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input52_A i_req_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4288__A _4500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4448__A2 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3656__B1 _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4853__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4227__S _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4751__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2890_ _2928_/A _3799_/B _3799_/A vssd1 vssd1 vccd1 vccd1 _3283_/A sky130_fd_sc_hd__a21oi_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5453__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3187__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ _5766_/A _4560_/B vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__or2_1
XFILLER_128_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3511_ _5435_/Q input41/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3512_/A sky130_fd_sc_hd__mux2_1
X_4491_ _4491_/A _4491_/B _4491_/C vssd1 vssd1 vccd1 vccd1 _4491_/Y sky130_fd_sc_hd__nand3_1
X_3442_ _3442_/A vssd1 vssd1 vccd1 vccd1 _5400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4198__A _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3373_ input26/X _5421_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3373_/X sky130_fd_sc_hd__mux2_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _3790_/X _3948_/A _5235_/S vssd1 vssd1 vccd1 vccd1 _5112_/Y sky130_fd_sc_hd__a21oi_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5043_/A vssd1 vssd1 vccd1 vccd1 _5701_/D sky130_fd_sc_hd__clkbuf_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__A2 _5200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3976__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3132__A_N input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _5607_/Q _4822_/B _4826_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5607_/D sky130_fd_sc_hd__o211a_1
XFILLER_138_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3277__A _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3178__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4758_ _5578_/Q _4747_/B _4757_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5578_/D sky130_fd_sc_hd__o211a_1
X_3709_ _4059_/B vssd1 vssd1 vccd1 vccd1 _4000_/B sky130_fd_sc_hd__inv_2
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4689_ _4689_/A vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4127__A1 _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_255_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3886__A0 _5500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4836__A _5684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3638__B1 _3608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5476__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3886__S _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3169__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_251_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3629__B1 _3608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3650__A _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4841__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3991_ _5526_/Q _3923_/A _3990_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5526_/D sky130_fd_sc_hd__o211a_1
X_5730_ _5740_/CLK _5730_/D vssd1 vssd1 vccd1 vccd1 _5730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2942_ _5447_/Q vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5661_ _5674_/CLK _5661_/D vssd1 vssd1 vccd1 vccd1 _5661_/Q sky130_fd_sc_hd__dfxtp_4
X_2873_ _3281_/A _3277_/A vssd1 vssd1 vccd1 vccd1 _2949_/A sky130_fd_sc_hd__nand2_1
XFILLER_230_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4357__A1 _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4612_ _5198_/A _4611_/X _4532_/X vssd1 vssd1 vccd1 vccd1 _4612_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_276_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5592_ _5659_/CLK _5592_/D vssd1 vssd1 vccd1 vccd1 _5592_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4543_ _4600_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4543_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4474_ _4474_/A _4474_/B _4473_/X vssd1 vssd1 vccd1 vccd1 _4474_/X sky130_fd_sc_hd__or3b_2
XFILLER_143_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5349__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3425_ _5392_/Q _3029_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3426_/A sky130_fd_sc_hd__mux2_1
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3332__A2 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _2829_/B _5361_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3357_/A sky130_fd_sc_hd__mux2_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3310_/A _3802_/B _3287_/C _3287_/D vssd1 vssd1 vccd1 vccd1 _3292_/D sky130_fd_sc_hd__nor4_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3560__A _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5499__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5026_ _5694_/Q _5132_/A _5030_/S vssd1 vssd1 vccd1 vccd1 _5027_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4293__B1 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2904__A _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_186_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3020__A1 _2840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3859__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4520__A1 _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3087__A1 _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A i_mem_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4823__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4240__S _4240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output83_A _4987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2770__B1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3210_ _5656_/Q _3147_/A _3149_/A _5576_/Q vssd1 vssd1 vccd1 vccd1 _3210_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3314__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4190_ _4025_/Y _4036_/Y _4040_/X vssd1 vssd1 vccd1 vccd1 _4192_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__5641__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3141_ _5596_/Q _3133_/X _3135_/X _5612_/Q _3140_/X vssd1 vssd1 vccd1 vccd1 _3141_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_121_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_227_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_267_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3072_ _2967_/A _3027_/X _3018_/A vssd1 vssd1 vccd1 vccd1 _3072_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3078__A1 _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4923__B _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4578__A1 _5539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2695__A_N _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ _5522_/Q _3923_/A _3973_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5522_/D sky130_fd_sc_hd__o211a_1
X_5713_ _5716_/CLK _5713_/D vssd1 vssd1 vccd1 vccd1 _5713_/Q sky130_fd_sc_hd__dfxtp_1
X_2925_ _3281_/A _3277_/A vssd1 vssd1 vccd1 vccd1 _3775_/B sky130_fd_sc_hd__nor2_2
XFILLER_148_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4361__D _4499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5644_ _5650_/CLK _5644_/D vssd1 vssd1 vccd1 vccd1 _5644_/Q sky130_fd_sc_hd__dfxtp_4
X_2856_ input51/X _5415_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _3003_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5575_ _5675_/CLK _5575_/D vssd1 vssd1 vccd1 vccd1 _5575_/Q sky130_fd_sc_hd__dfxtp_2
X_2787_ _5628_/Q _2655_/X _2761_/X _5644_/Q vssd1 vssd1 vccd1 vccd1 _2787_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3555__A _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3553__A2 _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4526_ _4533_/C _4527_/C _5081_/A vssd1 vssd1 vccd1 vccd1 _4528_/B sky130_fd_sc_hd__a21o_1
XANTENNA__4750__A1 _5574_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4457_ _4484_/B _4484_/C _4478_/C _4457_/D vssd1 vssd1 vccd1 vccd1 _4457_/Y sky130_fd_sc_hd__nor4_2
XFILLER_171_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_131_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5770__A _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3305__A2 _2943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3408_ _3408_/A vssd1 vssd1 vccd1 vccd1 _5383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4388_ _4108_/C _4009_/Y _4041_/X _4322_/A vssd1 vssd1 vccd1 vccd1 _4389_/B sky130_fd_sc_hd__a31o_1
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input7_A i_mem_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4386__A _4386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3339_ _4987_/A vssd1 vssd1 vccd1 vccd1 _3340_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_258_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4266__B1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4805__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5009_ _5032_/A vssd1 vssd1 vccd1 vccd1 _5233_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2816__A1 _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5514__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3792__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5664__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4995__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5297__A2 _2785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_167 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_249_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_224_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output121_A _5553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2807__A1 _5685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_162 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2710_ _2727_/C _2775_/B _5653_/Q _2775_/D vssd1 vssd1 vccd1 vccd1 _2710_/X sky130_fd_sc_hd__and4b_1
XFILLER_185_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4980__A1 _5672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3690_ _5455_/Q _5454_/Q _3690_/C _3690_/D vssd1 vssd1 vccd1 vccd1 _3691_/B sky130_fd_sc_hd__or4_1
XFILLER_185_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2641_ _5675_/Q _2747_/D _2733_/A _2747_/B vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__and4_1
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4732__A1 _4658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5360_ _5716_/CLK _5360_/D vssd1 vssd1 vccd1 vccd1 _5360_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_160_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4311_ _2904_/X _4036_/A _4034_/X _5445_/Q vssd1 vssd1 vccd1 vccd1 _4311_/X sky130_fd_sc_hd__a22o_1
XFILLER_153_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _5740_/Q _5775_/A _5291_/S vssd1 vssd1 vccd1 vccd1 _5292_/B sky130_fd_sc_hd__mux2_1
X_4242_ _5445_/Q _4010_/X _4239_/A _5449_/Q vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__a22o_1
XFILLER_259_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3299__A1 _5365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4173_ _4149_/X _4150_/X _4151_/X _4154_/X _4447_/S _4146_/A vssd1 vssd1 vccd1 vccd1
+ _4173_/X sky130_fd_sc_hd__mux4_1
XFILLER_255_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3124_ _3124_/A vssd1 vssd1 vccd1 vccd1 _3124_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3055_ _3060_/B _3055_/B vssd1 vssd1 vccd1 vccd1 _3055_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5537__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4145__S _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3269__B _5473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3223__A1 _5675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _3948_/B _3955_/X _3956_/Y _3965_/A vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3223__B2 _5595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3984__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5765__A _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2908_ _5364_/Q _5363_/Q _5362_/Q vssd1 vssd1 vccd1 vccd1 _3281_/B sky130_fd_sc_hd__nor3b_1
XANTENNA__4971__A1 _5668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3888_ _3888_/A vssd1 vssd1 vccd1 vccd1 _5500_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5687__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2982__B1 _2840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5627_ _5658_/CLK _5627_/D vssd1 vssd1 vccd1 vccd1 _5627_/Q sky130_fd_sc_hd__dfxtp_2
X_2839_ input37/X _5431_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2840_/D sky130_fd_sc_hd__mux2_2
XFILLER_191_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4184__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3526__A2 _5469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4723__A1 _5563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5558_ _5675_/CLK _5558_/D vssd1 vssd1 vccd1 vccd1 _5558_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_191_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2710__A_N _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4509_ _5532_/Q _4458_/A _4507_/Y _4508_/Y _4487_/X vssd1 vssd1 vccd1 vccd1 _5532_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_104_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5489_ _5722_/CLK _5489_/D vssd1 vssd1 vccd1 vccd1 _5489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4828__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3732__B _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4844__A _5614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3214__A1 _5609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3214__B2 _5625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4962__A1 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4714__A1 _5561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output169_A _3087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_338 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3150__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4325__S0 _4302_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4245__A3 _4236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4860_ _5621_/Q _4859_/B _4859_/Y _4840_/X vssd1 vssd1 vccd1 vccd1 _5621_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4192__C _4192_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3811_ _5473_/Q _5377_/Q _3813_/S vssd1 vssd1 vccd1 vccd1 _3812_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3205__B2 _5575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4791_ _5331_/A vssd1 vssd1 vccd1 vccd1 _4791_/X sky130_fd_sc_hd__buf_4
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3742_ _5623_/Q _3597_/X _3598_/X _5607_/Q _3741_/X vssd1 vssd1 vccd1 vccd1 _3742_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4953__A1 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3673_ _3673_/A _3673_/B _4076_/A vssd1 vssd1 vccd1 vccd1 _3683_/A sky130_fd_sc_hd__nand3_2
XFILLER_185_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5412_ _5757_/CLK _5412_/D vssd1 vssd1 vccd1 vccd1 _5412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput102 _5762_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[2] sky130_fd_sc_hd__buf_2
XANTENNA__2716__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 _5560_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[12] sky130_fd_sc_hd__buf_2
Xoutput124 _5556_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[8] sky130_fd_sc_hd__buf_2
X_5343_ _5680_/CLK _5343_/D vssd1 vssd1 vccd1 vccd1 _5343_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput135 _5690_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[1] sky130_fd_sc_hd__buf_2
XANTENNA__4929__A _5651_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput146 _3120_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[11] sky130_fd_sc_hd__buf_2
Xoutput157 _3112_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[7] sky130_fd_sc_hd__buf_2
XFILLER_99_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput168 _3082_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[13] sky130_fd_sc_hd__buf_2
Xoutput179 _3064_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[9] sky130_fd_sc_hd__buf_2
X_5274_ _5292_/A _5274_/B vssd1 vssd1 vccd1 vccd1 _5275_/A sky130_fd_sc_hd__and2_1
XFILLER_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4225_ _4454_/A _4223_/X _4224_/X _4271_/A vssd1 vssd1 vccd1 vccd1 _4225_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_87_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3141__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4156_ _4306_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4396_/A sky130_fd_sc_hd__xnor2_4
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3239__A_N _5478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3979__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4316__S0 _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3107_ _5709_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3108_/A sky130_fd_sc_hd__and2_1
XANTENNA__4664__A _5551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4087_ _4087_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__xor2_1
XFILLER_255_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3038_ _4552_/B _3010_/X _3036_/Y _3037_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3038_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_102_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4989_ _5235_/S vssd1 vssd1 vccd1 vccd1 _5032_/A sky130_fd_sc_hd__inv_2
XFILLER_211_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4944__A1 _5657_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4839__A _5612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5121__B2 _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5702__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4475__A3 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3889__S _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4632__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2756__A_N _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3199__B1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3918__A _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3738__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4513__S _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 i_mem_data[2] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
Xinput26 i_req_data[11] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 i_req_data[21] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 i_req_data[31] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4148__C1 _4128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4749__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2713__A3 _2711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3910__A2 _3843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_269_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5382__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3123__A0 _5709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4010_ _4024_/A _4024_/B vssd1 vssd1 vccd1 vccd1 _4010_/X sky130_fd_sc_hd__and2_1
XFILLER_284_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3674__A1 _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4484__A _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2882__C1 _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4912_ _5686_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4912_/Y sky130_fd_sc_hd__nand2_8
XFILLER_252_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5179__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4843_ _4653_/X _4836_/Y _4842_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5613_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2732__A _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3729__A2 _3605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4926__A1 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4774_ _4668_/X _4761_/Y _4773_/X _4769_/X vssd1 vssd1 vccd1 vccd1 _5584_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2937__B1 _3799_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3725_ _5557_/Q _3596_/X _3722_/X _3724_/X vssd1 vssd1 vccd1 vccd1 _4130_/B sky130_fd_sc_hd__o22a_4
XFILLER_106_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3656_ _5615_/Q _3597_/A _3598_/A _5599_/Q vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__a22o_1
XFILLER_228_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4154__A2 _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4659__A _5550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3587_ _5479_/Q _3532_/X _3584_/X _4006_/A _4006_/B vssd1 vssd1 vccd1 vccd1 _3619_/B
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5725__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3362__A0 _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5326_ _5755_/Q _5295_/X _5325_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5755_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5103__A1 _5707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5257_ _5729_/Q _4552_/B _5285_/S vssd1 vssd1 vccd1 vccd1 _5258_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4097__C _4192_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_57_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4208_ _4193_/X _4208_/B _4208_/C vssd1 vssd1 vccd1 vccd1 _4503_/A sky130_fd_sc_hd__and3b_4
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3665__A1 _5661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5188_ _4600_/B _5187_/Y _5231_/S vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3665__B2 _5645_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _4229_/A _4139_/B vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__2907__A _3304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4614__B1 _4634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3148__C_N input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4569__A _5519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4288__B _5015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A i_req_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3656__A1 _5615_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3656__B2 _5599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4454__D _4454_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output201_A _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4751__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__A _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_175_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5748__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3510_ _3510_/A vssd1 vssd1 vccd1 vccd1 _5434_/D sky130_fd_sc_hd__clkbuf_1
X_4490_ _4600_/B _4490_/B vssd1 vssd1 vccd1 vccd1 _4491_/C sky130_fd_sc_hd__xor2_1
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3441_ _5400_/Q _3068_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3442_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4479__A _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3372_/A vssd1 vssd1 vccd1 vccd1 _5368_/D sky130_fd_sc_hd__clkbuf_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4198__B _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _4543_/B _5156_/B _5108_/Y _5110_/X _3790_/X vssd1 vssd1 vccd1 vccd1 _5111_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5701_/Q _4617_/Y _5135_/S vssd1 vssd1 vccd1 vccd1 _5043_/A sky130_fd_sc_hd__mux2_1
XFILLER_257_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2727__A _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_280_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4072__A1 _4071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4826_ _4976_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4983_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_239_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3992__S _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3583__A0 _5482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5773__A _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3708_ _5560_/Q _3596_/X _3705_/X _3707_/X vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__o22a_4
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4780__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4688_ _5677_/Q _4690_/A vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4127__A2 _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3639_ _5635_/Q _3605_/A _3606_/A _3638_/X vssd1 vssd1 vccd1 vccd1 _3639_/X sky130_fd_sc_hd__a211o_1
XFILLER_255_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3293__A _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3886__A1 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5309_ _5747_/Q _5327_/B vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__or2_1
XANTENNA__5088__B1 _5086_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3638__A1 _5571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3638__B2 _5587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2637__A _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_231_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4852__A _5618_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3023__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3574__A0 _5485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3915__B _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3407__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3326__B1 _3325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5079__B1 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_239_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3629__A1 _5568_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3629__B2 _5584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5420__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _3990_/A _3990_/B vssd1 vssd1 vccd1 vccd1 _3990_/X sky130_fd_sc_hd__or2_1
XFILLER_222_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2941_ _2941_/A vssd1 vssd1 vccd1 vccd1 _5445_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3801__A1 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5069__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5570__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5003__A0 _5684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5660_ _5747_/CLK _5660_/D vssd1 vssd1 vccd1 vccd1 _5660_/Q sky130_fd_sc_hd__dfxtp_4
X_2872_ _5358_/Q vssd1 vssd1 vccd1 vccd1 _3277_/A sky130_fd_sc_hd__buf_4
XANTENNA__3097__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4611_ _4626_/S _5200_/A _4610_/Y _5294_/A vssd1 vssd1 vccd1 vccd1 _4611_/X sky130_fd_sc_hd__a211o_1
X_5591_ _5658_/CLK _5591_/D vssd1 vssd1 vccd1 vccd1 _5591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4542_ _5516_/Q _4599_/B vssd1 vssd1 vccd1 vccd1 _4542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5306__A1 _2760_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4473_ _4468_/A _3556_/X _3615_/X _4468_/X _4472_/Y vssd1 vssd1 vccd1 vccd1 _4473_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4002__A _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3424_ _3424_/A vssd1 vssd1 vccd1 vccd1 _5391_/D sky130_fd_sc_hd__clkbuf_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4937__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3355_ _3355_/A vssd1 vssd1 vccd1 vccd1 _5360_/D sky130_fd_sc_hd__clkbuf_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3800_/C _3791_/B _3309_/A _3285_/X vssd1 vssd1 vccd1 vccd1 _3287_/D sky130_fd_sc_hd__or4b_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3560__B _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5025_ _5025_/A vssd1 vssd1 vccd1 vccd1 _5693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5768__A _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2891__S _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4596__A2 _4595_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3288__A _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4809_ _4663_/X _4799_/Y _4808_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _5599_/D sky130_fd_sc_hd__o211a_2
XFILLER_166_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2920__A _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3859__A1 _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3751__A _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5443__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_236_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4284__A1 _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3087__A2 _3063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4284__B2 _5453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5593__CLK _5659_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output199_A _5319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2770__A1 _5566_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2770__B2 _5598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output76_A _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4757__A _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3661__A _4301_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _5660_/Q _3137_/X _3139_/X _5580_/Q vssd1 vssd1 vccd1 vccd1 _3140_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3071_ _3085_/A _3075_/B _3071_/C vssd1 vssd1 vccd1 vccd1 _3071_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4275__A1 _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_282_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_250_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2724__B _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3973_ _3990_/A _3973_/B vssd1 vssd1 vccd1 vccd1 _3973_/X sky130_fd_sc_hd__or2_1
XANTENNA__3786__B1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5712_ _5716_/CLK _5712_/D vssd1 vssd1 vccd1 vccd1 _5712_/Q sky130_fd_sc_hd__dfxtp_1
X_2924_ _5361_/Q _5360_/Q vssd1 vssd1 vccd1 vccd1 _2946_/A sky130_fd_sc_hd__nor2_2
XFILLER_210_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_224 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5643_ _5658_/CLK _5643_/D vssd1 vssd1 vccd1 vccd1 _5643_/Q sky130_fd_sc_hd__dfxtp_2
X_2855_ input52/X _5416_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _3003_/A sky130_fd_sc_hd__mux2_2
X_5574_ _5675_/CLK _5574_/D vssd1 vssd1 vccd1 vccd1 _5574_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_163_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3002__A2 _2850_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2786_ _5580_/Q _2635_/Y _2657_/X _5660_/Q vssd1 vssd1 vccd1 vccd1 _2786_/X sky130_fd_sc_hd__a22o_1
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4525_ _5229_/S _4522_/X _4523_/Y _4524_/X vssd1 vssd1 vccd1 vccd1 _4525_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4750__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5466__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4456_ _4350_/A _4406_/Y _4440_/X _4443_/X _4455_/X vssd1 vssd1 vccd1 vccd1 _4457_/D
+ sky130_fd_sc_hd__a311o_4
XFILLER_171_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3407_ _2850_/A _5383_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3408_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3305__A3 _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4387_ _4387_/A _4387_/B vssd1 vssd1 vccd1 vccd1 _4387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3338_ _3795_/A _3318_/C _3310_/X _3337_/X vssd1 vssd1 vccd1 vccd1 _5353_/D sky130_fd_sc_hd__o31a_1
XANTENNA__4386__B _4386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4266__A1 _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3269_ _5472_/Q _5473_/Q _3860_/B vssd1 vssd1 vccd1 vccd1 _3838_/C sky130_fd_sc_hd__nor3b_1
XFILLER_252_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5008_/A vssd1 vssd1 vccd1 vccd1 _5686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_233_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3777__A0 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3529__A0 _5473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3746__A _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2650__A _4635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5724_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4577__A _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4257__A1 _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4257__B2 _4171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2807__A2 _5686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output114_A _5561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5339__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3768__A0 _5408_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4980__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5489__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2640_ _5346_/Q vssd1 vssd1 vccd1 vccd1 _2733_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4732__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2710__D _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4310_ _2919_/X _4034_/A _4333_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__a211o_1
XFILLER_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _5290_/A vssd1 vssd1 vccd1 vccd1 _5739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_273_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4241_ _5450_/Q _4326_/A _3692_/X _4024_/B _5452_/Q vssd1 vssd1 vccd1 vccd1 _4241_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_259_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4487__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3299__A2 _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ _4396_/A vssd1 vssd1 vccd1 vccd1 _4471_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _5709_/Q _5717_/Q _4651_/S vssd1 vssd1 vccd1 vccd1 _3124_/A sky130_fd_sc_hd__mux2_1
XFILLER_222_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3054_ _5397_/Q _3053_/C _5398_/Q vssd1 vssd1 vccd1 vccd1 _3055_/B sky130_fd_sc_hd__a21oi_1
XFILLER_208_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_222_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4950__A _5687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3956_ _3956_/A _3993_/B vssd1 vssd1 vccd1 vccd1 _3956_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3223__A2 _3137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2907_ _3304_/A _2922_/A vssd1 vssd1 vccd1 vccd1 _2957_/B sky130_fd_sc_hd__nor2_1
XFILLER_188_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3887_ _3893_/A _3887_/B vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__and2_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4971__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3566__A _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5257__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5626_ _5658_/CLK _5626_/D vssd1 vssd1 vccd1 vccd1 _5626_/Q sky130_fd_sc_hd__dfxtp_1
X_2838_ input31/X _5426_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2840_/C sky130_fd_sc_hd__mux2_2
XFILLER_176_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2719__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4184__B1 _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3526__A3 _3761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5557_ _5675_/CLK _5557_/D vssd1 vssd1 vccd1 vccd1 _5557_/Q sky130_fd_sc_hd__dfxtp_4
X_2769_ _5662_/Q _2774_/C _2789_/B _2789_/C vssd1 vssd1 vccd1 vccd1 _2769_/X sky130_fd_sc_hd__and4_1
X_4508_ _3948_/A _4485_/A _4458_/A vssd1 vssd1 vccd1 vccd1 _4508_/Y sky130_fd_sc_hd__o21ai_1
X_5488_ _5722_/CLK _5488_/D vssd1 vssd1 vccd1 vccd1 _5488_/Q sky130_fd_sc_hd__dfxtp_1
X_4439_ _4055_/B _4403_/X _4052_/A vssd1 vssd1 vccd1 vccd1 _4440_/B sky130_fd_sc_hd__o21a_1
XANTENNA__3505__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4844__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3998__B1 _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2670__B1 _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3214__A2 _3133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5631__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4962__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5167__S _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3922__B1 _3851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3415__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2685__A_N _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4457__D _4457_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3150__A1 _5644_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3150__B2 _5564_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4325__S1 _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4650__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3810_ _3810_/A vssd1 vssd1 vccd1 vccd1 _5472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4938__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4790_ _4978_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4790_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3205__A2 _3147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3741_ _5671_/Q _3600_/X _3602_/X _5655_/Q vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__a22o_1
XFILLER_220_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4953__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5077__S _5077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3672_ _3561_/X _3564_/X _3569_/X _3596_/A _5548_/Q vssd1 vssd1 vccd1 vccd1 _4076_/A
+ sky130_fd_sc_hd__o32ai_4
XFILLER_173_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5411_ _5757_/CLK _5411_/D vssd1 vssd1 vccd1 vccd1 _5411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput103 _5763_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[3] sky130_fd_sc_hd__buf_2
XANTENNA__2716__A1 _5636_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5342_ _5686_/CLK _5342_/D vssd1 vssd1 vccd1 vccd1 _5342_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2716__B2 _5668_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput114 _5561_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[13] sky130_fd_sc_hd__buf_2
Xoutput125 _5557_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[9] sky130_fd_sc_hd__buf_2
Xoutput136 _5691_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[2] sky130_fd_sc_hd__buf_2
XANTENNA__4929__B _4931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput147 _3122_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[12] sky130_fd_sc_hd__buf_2
Xoutput158 _3114_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[8] sky130_fd_sc_hd__buf_2
X_5273_ _5734_/Q _4590_/B _5285_/S vssd1 vssd1 vccd1 vccd1 _5274_/B sky130_fd_sc_hd__mux2_1
Xoutput169 _3087_/X vssd1 vssd1 vccd1 vccd1 o_req_addr[14] sky130_fd_sc_hd__buf_2
XFILLER_217_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4224_ _4276_/A _4307_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__or3b_1
XANTENNA__4010__A _4024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_233_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3141__A1 _5596_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3141__B2 _5612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5504__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4155_ _4248_/C _4154_/X _4449_/S vssd1 vssd1 vccd1 vccd1 _4198_/C sky130_fd_sc_hd__mux2_1
XANTENNA__4945__A _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3106_ _3106_/A vssd1 vssd1 vccd1 vccd1 _3106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_228_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _4240_/S _4239_/B _4239_/A vssd1 vssd1 vccd1 vccd1 _4090_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__4316__S1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3037_ _2840_/B _3027_/X _3343_/C vssd1 vssd1 vccd1 vccd1 _3037_/X sky130_fd_sc_hd__a21o_1
XFILLER_255_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4680__A _5554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4988_ _5263_/A _4988_/B vssd1 vssd1 vccd1 vccd1 _5235_/S sky130_fd_sc_hd__nand2_4
XFILLER_23_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4944__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3939_ _4523_/B _3948_/B vssd1 vssd1 vccd1 vccd1 _3939_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2955__A1 _3308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2955__B2 _3307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4157__B1 _4396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5609_ _5675_/CLK _5609_/D vssd1 vssd1 vccd1 vccd1 _5609_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_124_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4839__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4880__A1 _4653_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2891__A0 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4632__A1 _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4590__A _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3199__A1 _5606_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3199__B2 _5622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 i_mem_data[3] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
XFILLER_167_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 i_req_data[12] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_167_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput38 i_req_data[22] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4148__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput49 i_req_data[3] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output181_A _5470_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4749__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5527__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5112__A2 _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3674__A2 _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__A1 _5626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5677__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2882__B1 _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4623__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4911_ _5643_/Q _4897_/B _4910_/Y _4908_/X vssd1 vssd1 vccd1 vccd1 _5643_/D sky130_fd_sc_hd__o211a_1
XFILLER_252_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2700__A_N _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4842_ _5613_/Q _4872_/B vssd1 vssd1 vccd1 vccd1 _4842_/X sky130_fd_sc_hd__or2_1
X_4773_ _5584_/Q _4781_/A vssd1 vssd1 vccd1 vccd1 _4773_/X sky130_fd_sc_hd__or2_1
XANTENNA__4926__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _5637_/Q _3605_/X _3606_/X _3723_/X vssd1 vssd1 vccd1 vccd1 _3724_/X sky130_fd_sc_hd__a211o_1
XFILLER_146_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4005__A _4108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3655_ _5550_/Q _3596_/X _3652_/X _3654_/X vssd1 vssd1 vccd1 vccd1 _4083_/B sky130_fd_sc_hd__o22a_4
XFILLER_228_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3586_ _2715_/X _2716_/X _2719_/X _2720_/X _3588_/S vssd1 vssd1 vccd1 vccd1 _4006_/B
+ sky130_fd_sc_hd__o311a_2
X_5325_ _5325_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__or2_1
XANTENNA__5103__A2 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5256_ _5291_/S vssd1 vssd1 vccd1 vccd1 _5285_/S sky130_fd_sc_hd__clkbuf_4
X_4207_ _4199_/Y _4202_/Y _4271_/B _4454_/D _4206_/Y vssd1 vssd1 vccd1 vccd1 _4208_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4675__A _5553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5187_ _5192_/A _5187_/B vssd1 vssd1 vccd1 vccd1 _5187_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_228_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5270__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3665__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _4300_/S _4138_/B vssd1 vssd1 vccd1 vccd1 _4138_/Y sky130_fd_sc_hd__nand2_1
XFILLER_228_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4069_ _4467_/A _4232_/B _4069_/C vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__or3_1
XFILLER_260_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4614__A1 _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2923__A _3284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_269_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4550__A0 _5307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4302__A0 _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input38_A i_req_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4585__A _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4853__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3656__A2 _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2723__A_N _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5030__A1 _5156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5318__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3664__A _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3440_ _3440_/A vssd1 vssd1 vccd1 vccd1 _5399_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4479__B _4485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4541__B1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3371_ _3001_/D _5368_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5200_/B _5131_/A vssd1 vssd1 vccd1 vccd1 _5110_/X sky130_fd_sc_hd__and2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A vssd1 vssd1 vccd1 vccd1 _5700_/D sky130_fd_sc_hd__clkbuf_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2727__B _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_280_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4072__A2 _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2743__A _3956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3280__B1 _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4216__A1_N _3750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3558__B _4372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4825_ _5606_/Q _4822_/B _4824_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5606_/D sky130_fd_sc_hd__o211a_1
XFILLER_166_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _5577_/Q _4747_/B _4755_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5577_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3583__A1 _5321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3707_ _5640_/Q _3605_/X _3606_/X _3706_/X vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__a211o_1
X_4687_ _4687_/A vssd1 vssd1 vccd1 vccd1 _4697_/A sky130_fd_sc_hd__buf_2
X_3638_ _5571_/Q _3607_/A _3608_/A _5587_/Q vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__a22o_1
XFILLER_108_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3569_ _5564_/Q _3607_/A _3606_/A _3567_/X _3568_/X vssd1 vssd1 vccd1 vccd1 _3569_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2689__A3 _2687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5308_ _5746_/Q _5295_/X _5307_/X _4979_/X vssd1 vssd1 vccd1 vccd1 _5746_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5088__A1 _5060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2746__A_N _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5239_ _5509_/Q _5263_/A _5253_/S vssd1 vssd1 vccd1 vccd1 _5240_/A sky130_fd_sc_hd__and3_1
XANTENNA__3513__S _3517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3638__A2 _3607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__A1 _5611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3740__C _4105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4852__B _4856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5260__A1 _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3271__B1 _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5372__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4692__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3574__A1 _2650_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3326__A1 _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_239_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2764__B_N _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3629__A2 _3607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3423__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_247_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4762__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5715__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2940_ _2936_/X _2939_/X _3337_/B vssd1 vssd1 vccd1 vccd1 _2941_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3801__A2 _2937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2871_ _5359_/Q vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__inv_2
XFILLER_200_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4610_ _4626_/S _5321_/A vssd1 vssd1 vccd1 vccd1 _4610_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5590_ _5623_/CLK _5590_/D vssd1 vssd1 vccd1 vccd1 _5590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4541_ _5763_/A _4511_/X _3919_/X _4540_/X vssd1 vssd1 vccd1 vccd1 _5535_/D sky130_fd_sc_hd__o211a_1
XFILLER_128_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4472_ _4468_/A _4471_/X _3556_/X vssd1 vssd1 vccd1 vccd1 _4472_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_209_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3423_ _5391_/Q _3023_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3424_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4002__B _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3354_ _2829_/A _5360_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3355_/A sky130_fd_sc_hd__mux2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4937__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _5361_/Q _3317_/A _2945_/B _3780_/B _2938_/X vssd1 vssd1 vccd1 vccd1 _3285_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5114__A _5517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5024_ _5693_/Q _4499_/B _5030_/S vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__mux2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3138__C_N input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5395__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3288__B _3292_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_264 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4808_ _5599_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4808_/X sky130_fd_sc_hd__or2_1
XANTENNA__3005__B1 _3004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4739_ _5570_/Q _4743_/A vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__or2_1
XFILLER_266_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4505__B1 _4504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3859__A2 _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3751__B _3751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5738__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_244_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3244__B1 _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_125_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2770__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4757__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output69_A _3157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3070_ _5400_/Q _3069_/C _5401_/Q vssd1 vssd1 vccd1 vccd1 _3071_/C sky130_fd_sc_hd__a21oi_1
XFILLER_94_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4773__A _5584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4432__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3972_ _3971_/X _5317_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2724__C _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3786__A1 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5711_ _5757_/CLK _5711_/D vssd1 vssd1 vccd1 vccd1 _5711_/Q sky130_fd_sc_hd__dfxtp_1
X_2923_ _3284_/B _2923_/B vssd1 vssd1 vccd1 vccd1 _3800_/C sky130_fd_sc_hd__nor2_1
XFILLER_188_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5642_ _5658_/CLK _5642_/D vssd1 vssd1 vccd1 vccd1 _5642_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2854_ input50/X _5414_/Q _3768_/S vssd1 vssd1 vccd1 vccd1 _3004_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2740__B _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5573_ _5675_/CLK _5573_/D vssd1 vssd1 vccd1 vccd1 _5573_/Q sky130_fd_sc_hd__dfxtp_4
X_2785_ _3935_/A vssd1 vssd1 vccd1 vccd1 _2785_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__5109__A _5109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3555__C _3555_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4013__A _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4524_ _5514_/Q _5459_/Q vssd1 vssd1 vccd1 vccd1 _4524_/X sky130_fd_sc_hd__and2_1
XFILLER_156_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_236_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4455_ _4455_/A _4455_/B _4454_/X vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__or3b_1
X_3406_ _3406_/A vssd1 vssd1 vccd1 vccd1 _5382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_277_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4386_ _4386_/A _4386_/B _4386_/C vssd1 vssd1 vccd1 vccd1 _4387_/B sky130_fd_sc_hd__and3_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3337_ _5353_/Q _3337_/B vssd1 vssd1 vccd1 vccd1 _3337_/X sky130_fd_sc_hd__or2_1
XFILLER_252_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_258_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _5471_/Q vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__inv_2
XANTENNA__4266__A2 _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _5686_/Q _5340_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _5008_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3199_ _5606_/Q _3133_/A _3135_/A _5622_/Q _3198_/X vssd1 vssd1 vccd1 vccd1 _3199_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4671__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3226__B1 _3145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3777__A1 _3775_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3529__A1 _2768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5410__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_107_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3762__A _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4577__B _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3701__A1 _5561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5560__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A i_mem_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4593__A _5522_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__A3 _5687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4193__A1 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4193__B2 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4768__A _5582_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4240_ _4239_/A _4239_/X _4240_/S vssd1 vssd1 vccd1 vccd1 _4240_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4171_ _4171_/A _4171_/B _4171_/C vssd1 vssd1 vccd1 vccd1 _4171_/X sky130_fd_sc_hd__or3_1
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _3122_/A vssd1 vssd1 vccd1 vccd1 _3122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3053_ _5398_/Q _5397_/Q _3053_/C vssd1 vssd1 vccd1 vccd1 _3060_/B sky130_fd_sc_hd__and3_1
XFILLER_67_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2735__B _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_284 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2957__A_N _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4008__A _4108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3208__B1 _3139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4950__B _4950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3955_ _5766_/A _5731_/Q _5329_/A vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3847__A _5263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2906_ _3317_/A _2922_/A vssd1 vssd1 vccd1 vccd1 _3283_/B sky130_fd_sc_hd__nor2_2
XANTENNA__5433__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3886_ _5500_/Q _5313_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3887_/B sky130_fd_sc_hd__mux2_1
XFILLER_176_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4708__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3566__B _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5625_ _5658_/CLK _5625_/D vssd1 vssd1 vccd1 vccd1 _5625_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_136_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2982__A2 _2850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2837_ input36/X _5430_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2840_/B sky130_fd_sc_hd__mux2_2
XFILLER_247_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4184__A1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4184__B2 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5556_ _5675_/CLK _5556_/D vssd1 vssd1 vccd1 vccd1 _5556_/Q sky130_fd_sc_hd__dfxtp_4
X_2768_ _3943_/A vssd1 vssd1 vccd1 vccd1 _2768_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_247_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4507_ _4507_/A _4507_/B vssd1 vssd1 vccd1 vccd1 _4507_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5583__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2699_ _5574_/Q _2644_/X _2695_/X _2697_/X _2698_/X vssd1 vssd1 vccd1 vccd1 _2699_/X
+ sky130_fd_sc_hd__a2111o_1
X_5487_ _5754_/CLK _5487_/D vssd1 vssd1 vccd1 vccd1 _5487_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5273__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _4438_/A _4438_/B vssd1 vssd1 vccd1 vccd1 _4478_/C sky130_fd_sc_hd__nor2_1
XFILLER_116_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4369_ _4370_/B _4387_/A _4370_/A vssd1 vssd1 vccd1 vccd1 _4371_/B sky130_fd_sc_hd__o21ai_1
XFILLER_258_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_342 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_258_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_246_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3521__S _3523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2670__B2 _5561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_127_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3922__A1 _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3150__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3431__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3989__A1 _5325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4650__A2 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2661__A1 _5578_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5456__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ _3747_/A _3747_/B _4105_/B vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__or3_1
XFILLER_158_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3610__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_150 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _4274_/A vssd1 vssd1 vccd1 vccd1 _4304_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_158_386 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4166__A1 _4171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5410_ _5757_/CLK _5410_/D vssd1 vssd1 vccd1 vccd1 _5410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput104 _5764_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[4] sky130_fd_sc_hd__buf_2
XANTENNA__2716__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput115 _5562_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[14] sky130_fd_sc_hd__buf_2
XFILLER_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5341_ _5680_/CLK _5341_/D vssd1 vssd1 vccd1 vccd1 _5341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput126 _5742_/Q vssd1 vssd1 vccd1 vccd1 o_c_data_page sky130_fd_sc_hd__buf_2
Xoutput137 _5692_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[3] sky130_fd_sc_hd__buf_2
Xoutput148 _3124_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[13] sky130_fd_sc_hd__buf_2
Xoutput159 _3116_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[9] sky130_fd_sc_hd__buf_2
X_5272_ _5272_/A vssd1 vssd1 vccd1 vccd1 _5733_/D sky130_fd_sc_hd__clkbuf_1
X_4223_ _4221_/X _4222_/X _4304_/S vssd1 vssd1 vccd1 vccd1 _4223_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4010__B _4024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4154_ _4132_/A _4281_/A _3613_/X _4469_/C _4469_/B vssd1 vssd1 vccd1 vccd1 _4154_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3141__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4945__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3105_ _5708_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3106_/A sky130_fd_sc_hd__and2_1
X_4085_ _4085_/A vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_233_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3036_ _3085_/A _3036_/B vssd1 vssd1 vccd1 vccd1 _3036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4961__A _5664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_i_clk clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 _5692_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_251_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ _4987_/A _4987_/B vssd1 vssd1 vccd1 vccd1 _5676_/D sky130_fd_sc_hd__nor2_1
X_3938_ _5081_/A _5727_/Q _5329_/A vssd1 vssd1 vccd1 vccd1 _3938_/X sky130_fd_sc_hd__mux2_1
XFILLER_258_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2955__A2 _2943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3869_ _3908_/B vssd1 vssd1 vccd1 vccd1 _3874_/B sky130_fd_sc_hd__buf_2
XFILLER_258_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4157__A1 _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5608_ _5674_/CLK _5608_/D vssd1 vssd1 vccd1 vccd1 _5608_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_11_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_142 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_164_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5539_ _5665_/CLK _5539_/D vssd1 vssd1 vccd1 vccd1 _5539_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4201__A _4372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_274_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3668__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4865__C1 _4862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4880__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5479__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4632__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4590__B _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5178__S _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3199__A2 _3133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 i_mem_data[4] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput28 i_req_data[13] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_210_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4148__A1 _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput39 i_req_data[23] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_182_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3659__B1 _3606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_284_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4871__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__C1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2882__B2 _2938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_252_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4910_ _4985_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_240_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4841_ _4646_/X _4836_/Y _4839_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _5612_/D sky130_fd_sc_hd__o211a_1
X_4772_ _4663_/X _4761_/Y _4771_/X _4769_/X vssd1 vssd1 vccd1 vccd1 _5583_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2937__A2 _3304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3723_ _5573_/Q _3607_/X _3608_/X _5589_/Q vssd1 vssd1 vccd1 vccd1 _3723_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4005__B _4130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3654_ _5630_/Q _3605_/X _3606_/X _3653_/X vssd1 vssd1 vccd1 vccd1 _3654_/X sky130_fd_sc_hd__a211o_1
XFILLER_146_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3585_ _5478_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _4006_/A sky130_fd_sc_hd__and2_1
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5324_ _5754_/Q _5295_/X _5323_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5754_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4956__A _5662_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5255_ _5255_/A vssd1 vssd1 vccd1 vccd1 _5728_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4847__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4206_ _2904_/X _4008_/X _4192_/C _2954_/X _4205_/X vssd1 vssd1 vccd1 vccd1 _4206_/Y
+ sky130_fd_sc_hd__a221oi_1
XANTENNA__4311__A1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4311__B2 _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5186_ _4599_/B _5185_/X _4599_/Y vssd1 vssd1 vccd1 vccd1 _5187_/B sky130_fd_sc_hd__o21ai_2
XFILLER_275_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4137_ _4394_/A _4127_/X _4131_/X _4133_/X _4447_/S _4469_/D vssd1 vssd1 vccd1 vccd1
+ _4138_/B sky130_fd_sc_hd__mux4_1
XFILLER_228_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4068_ _4467_/A _4232_/B _4069_/C vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__o21ai_1
X_3019_ _5391_/Q _5390_/Q vssd1 vssd1 vccd1 vccd1 _3019_/X sky130_fd_sc_hd__xor2_1
XANTENNA__3822__A0 _5478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4378__A1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2675__A_N _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3586__C1 _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4550__A1 _4499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4866__A _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4302__A1 _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4853__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3813__A0 _5474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4106__A _4130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3010__A _3063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3577__C1 _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3945__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3370_ _3419_/S vssd1 vssd1 vccd1 vccd1 _3394_/S sky130_fd_sc_hd__buf_4
XANTENNA__4541__A1 _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4829__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5700_/Q _5039_/Y _5135_/S vssd1 vssd1 vccd1 vccd1 _5041_/A sky130_fd_sc_hd__mux2_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2727__C _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4152__S0 _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3804__B1 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3280__A1 _2938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4824_ _4974_/A _4834_/B vssd1 vssd1 vccd1 vccd1 _4824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4755_ _4981_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4755_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3855__A _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4450__S _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4780__A1 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ _5576_/Q _3607_/X _3608_/X _5592_/Q vssd1 vssd1 vccd1 vccd1 _3706_/X sky130_fd_sc_hd__a22o_1
X_4686_ _4642_/Y _4684_/X _4685_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _5555_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3637_ _5619_/Q _3597_/A _3598_/X _5603_/Q vssd1 vssd1 vccd1 vccd1 _3637_/X sky130_fd_sc_hd__a22o_1
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3568_ _3599_/B _3601_/B _5644_/Q _3601_/C vssd1 vssd1 vccd1 vccd1 _3568_/X sky130_fd_sc_hd__and4b_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5307_ _5307_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__or2_1
XFILLER_255_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3499_ _5429_/Q input34/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__mux2_1
XFILLER_248_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5088__A2 _5077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5238_ _5238_/A vssd1 vssd1 vccd1 vccd1 _5722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_248_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4835__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5169_ _5179_/S _5167_/X _5168_/Y vssd1 vssd1 vccd1 vccd1 _5169_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2934__A _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5517__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3023__A1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3765__A _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5667__CLK _5667_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3326__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A i_req_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5079__A2 _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_262_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _3337_/B vssd1 vssd1 vccd1 vccd1 _5486_/D sky130_fd_sc_hd__buf_6
XFILLER_70_390 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4540_ _4532_/X _4534_/Y _4535_/X _4539_/Y _4529_/X vssd1 vssd1 vccd1 vccd1 _4540_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4471_ _4178_/X _4470_/X _4471_/S vssd1 vssd1 vccd1 vccd1 _4471_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3422_ _3422_/A vssd1 vssd1 vccd1 vccd1 _5390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3353_/A vssd1 vssd1 vccd1 vccd1 _5359_/D sky130_fd_sc_hd__clkbuf_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3304_/A _3284_/B _3775_/C vssd1 vssd1 vccd1 vccd1 _3780_/B sky130_fd_sc_hd__or3b_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5023_/A vssd1 vssd1 vccd1 vccd1 _5692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_285_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_241_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4807_ _4658_/X _4799_/Y _4806_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _5598_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2999_ input55/X _5419_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _3001_/C sky130_fd_sc_hd__mux2_1
XANTENNA__3585__A _5478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5276__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4738_ _4674_/X _4724_/Y _4737_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5569_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4669_ _5552_/Q _4687_/A vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__or2_1
XFILLER_174_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2929__A _3307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_384 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_276_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_236_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2819__B2 _5720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3244__A1 _5347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_109_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_140_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5215__A _5526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3180__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_94_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4265__S _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3971_ _5770_/A _5735_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3971_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2724__D _5603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5710_ _5716_/CLK _5710_/D vssd1 vssd1 vccd1 vccd1 _5710_/Q sky130_fd_sc_hd__dfxtp_1
X_2922_ _2922_/A _2945_/B vssd1 vssd1 vccd1 vccd1 _2923_/B sky130_fd_sc_hd__or2_1
XFILLER_250_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5641_ _5658_/CLK _5641_/D vssd1 vssd1 vccd1 vccd1 _5641_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_203_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2736__A_N _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2853_ _2830_/A _2852_/X _2829_/A _2829_/B vssd1 vssd1 vccd1 vccd1 _2853_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5572_ _5675_/CLK _5572_/D vssd1 vssd1 vccd1 vccd1 _5572_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__2740__C _5650_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2784_ _2779_/X _2780_/X _2783_/X _2791_/B _5549_/Q vssd1 vssd1 vccd1 vccd1 _3935_/A
+ sky130_fd_sc_hd__o32ai_4
X_4523_ _4600_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _4523_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5109__B _5109_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4013__B _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2886__A_N _5361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4454_ _4454_/A _4454_/B _4454_/C _4454_/D vssd1 vssd1 vccd1 vccd1 _4454_/X sky130_fd_sc_hd__or4_1
XFILLER_236_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3405_ _2845_/C _5382_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3406_/A sky130_fd_sc_hd__mux2_1
XFILLER_277_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2749__A _5553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4385_ _4385_/A vssd1 vssd1 vccd1 vccd1 _4600_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__3171__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5125__A _5125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3336_ _5352_/Q _3780_/A _3335_/X vssd1 vssd1 vccd1 vccd1 _5352_/D sky130_fd_sc_hd__o21a_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5362__CLK _5716_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_258_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _5465_/Q _3267_/B vssd1 vssd1 vccd1 vccd1 _3273_/A sky130_fd_sc_hd__nor2_1
XFILLER_252_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5006_ _5006_/A vssd1 vssd1 vccd1 vccd1 _5685_/D sky130_fd_sc_hd__clkbuf_1
X_3198_ _5670_/Q _3137_/A _3139_/A _5590_/Q vssd1 vssd1 vccd1 vccd1 _3198_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_226_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3226__A1 _5643_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4423__B1 _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2985__B1 _2840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3519__S _3523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_277_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5705__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5151__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3701__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4874__A _5685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_249_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4257__A3 _4014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4662__A0 _5707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A i_mem_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3217__A1 _5561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3429__S _3435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4768__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output81_A _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5385__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_259_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3153__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4170_ _4441_/B _4112_/X _4110_/X _4111_/Y vssd1 vssd1 vccd1 vccd1 _4171_/C sky130_fd_sc_hd__o211a_1
X_3121_ _5708_/Q _5716_/Q _4651_/S vssd1 vssd1 vccd1 vccd1 _3122_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4784__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3052_ _5539_/Q _3010_/X _3050_/Y _3051_/X _3016_/A vssd1 vssd1 vccd1 vccd1 _3052_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_255_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2735__C _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3208__A1 _5672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4008__B _4130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3208__B2 _5592_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3954_ _5517_/Q _3923_/X _3953_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5517_/D sky130_fd_sc_hd__o211a_1
X_2905_ _5359_/Q _3277_/A vssd1 vssd1 vccd1 vccd1 _2943_/C sky130_fd_sc_hd__nor2_4
X_3885_ _3885_/A vssd1 vssd1 vccd1 vccd1 _5499_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3566__C _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5624_ _5658_/CLK _5624_/D vssd1 vssd1 vccd1 vccd1 _5624_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4024__A _4024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2836_ input32/X _5427_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2840_/A sky130_fd_sc_hd__mux2_2
XFILLER_247_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4184__A2 _4045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5555_ _5747_/CLK _5555_/D vssd1 vssd1 vccd1 vccd1 _5555_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__2814__S0 _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4959__A _5663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2767_ _2762_/X _2763_/X _2766_/X _2791_/B _5551_/Q vssd1 vssd1 vccd1 vccd1 _3943_/A
+ sky130_fd_sc_hd__o32ai_4
XANTENNA__5728__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3392__A0 _2850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4506_ _4504_/Y _4494_/X _4495_/Y _4289_/C vssd1 vssd1 vccd1 vccd1 _4507_/B sky130_fd_sc_hd__a31o_1
X_5486_ _5743_/CLK _5486_/D vssd1 vssd1 vccd1 vccd1 _5486_/Q sky130_fd_sc_hd__dfxtp_1
X_2698_ _5670_/Q _2806_/A _2771_/A _2771_/B vssd1 vssd1 vccd1 vccd1 _2698_/X sky130_fd_sc_hd__and4_1
XANTENNA__5133__A1 _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4437_ _4484_/A vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__inv_2
XFILLER_104_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4368_ _4368_/A _4368_/B vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3695__A1 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input5_A i_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3319_ _3319_/A _3791_/D vssd1 vssd1 vccd1 vccd1 _3335_/B sky130_fd_sc_hd__or2_1
XFILLER_258_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4299_ _4394_/A _4127_/X _4148_/X _4149_/X _4272_/S _4146_/A vssd1 vssd1 vccd1 vccd1
+ _4299_/X sky130_fd_sc_hd__mux4_1
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3447__A1 _3082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2926__B _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3998__A2 _4289_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3301__A1_N _5365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3103__A _5707_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3922__A2 _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3948__A _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2852__A _2852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3610__A1 _5643_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3670_ _3585_/B _3935_/A _3536_/Y vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__o21a_4
XFILLER_185_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2998__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4779__A _5587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3683__A _3683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5340_ _5707_/CLK _5340_/D vssd1 vssd1 vccd1 vccd1 _5340_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4571__C1 _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 _5765_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[5] sky130_fd_sc_hd__buf_2
Xoutput116 _5563_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[15] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput127 _5508_/Q vssd1 vssd1 vccd1 vccd1 o_c_instr_page sky130_fd_sc_hd__buf_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput138 _5693_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[4] sky130_fd_sc_hd__buf_2
XANTENNA__5115__A1 _5517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput149 _3126_/X vssd1 vssd1 vccd1 vccd1 o_mem_data[14] sky130_fd_sc_hd__buf_2
XANTENNA__5115__B2 _5497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5271_ _5292_/A _5271_/B vssd1 vssd1 vccd1 vccd1 _5272_/A sky130_fd_sc_hd__and2_1
XFILLER_141_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4222_ _3710_/X _3747_/X _4231_/S vssd1 vssd1 vccd1 vccd1 _4222_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ _4300_/S _4153_/B vssd1 vssd1 vccd1 vccd1 _4347_/B sky130_fd_sc_hd__or2_1
XFILLER_255_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3104_ _3104_/A vssd1 vssd1 vccd1 vccd1 _3104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_233_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4084_ _4010_/X _4084_/B vssd1 vssd1 vccd1 vccd1 _4085_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4626__A0 _5325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3035_ _5394_/Q _3039_/C vssd1 vssd1 vccd1 vccd1 _3036_/B sky130_fd_sc_hd__xnor2_1
XFILLER_270_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4986_ _5675_/Q _4972_/B _4985_/Y _4979_/X vssd1 vssd1 vccd1 vccd1 _5675_/D sky130_fd_sc_hd__o211a_1
X_3937_ _5513_/Q _3923_/X _3936_/X _3848_/X vssd1 vssd1 vccd1 vccd1 _5513_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5550__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3868_ _3868_/A vssd1 vssd1 vccd1 vccd1 _5492_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_164_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5607_ _5623_/CLK _5607_/D vssd1 vssd1 vccd1 vccd1 _5607_/Q sky130_fd_sc_hd__dfxtp_2
X_2819_ _5757_/Q _2818_/Y _5679_/Q _5720_/Q vssd1 vssd1 vccd1 vccd1 _5331_/B sky130_fd_sc_hd__a22o_2
XFILLER_164_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3799_ _3799_/A _3799_/B vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_191_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5538_ _5665_/CLK _5538_/D vssd1 vssd1 vccd1 vccd1 _5766_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_11_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5106__A1 _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5469_ _5707_/CLK _5469_/D vssd1 vssd1 vccd1 vccd1 _5469_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__3117__A0 _5706_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3668__A1 _5629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5313__A _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_302 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput18 i_mem_data[5] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 i_req_data[14] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4148__A2 _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4599__A _5523_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3356__A0 _2829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3008__A _5760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3659__A1 _5631_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5423__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_374 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_252_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_240_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5573__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4273__S _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4840_ _4979_/A vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__clkbuf_8
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _5583_/Q _4797_/B vssd1 vssd1 vccd1 vccd1 _4771_/X sky130_fd_sc_hd__or2_1
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3722_ _5621_/Q _3597_/X _3598_/X _5605_/Q _3721_/X vssd1 vssd1 vccd1 vccd1 _3722_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4792__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3653_ _5566_/Q _3607_/X _3608_/X _5582_/Q vssd1 vssd1 vccd1 vccd1 _3653_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_228_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4544__C1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3584_ _2705_/X _2706_/X _2711_/X _2712_/X _3588_/S vssd1 vssd1 vccd1 vccd1 _3584_/X
+ sky130_fd_sc_hd__o311a_2
XFILLER_228_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5323_ _5323_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__or2_1
XFILLER_114_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4021__B _4027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5254_ _5261_/A _5254_/B vssd1 vssd1 vccd1 vccd1 _5255_/A sky130_fd_sc_hd__and2_1
XFILLER_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4956__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4205_ _2919_/X _4108_/A _4130_/B _4333_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4205_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5185_ _5771_/A _5193_/B _5184_/Y _5196_/A vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3352__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _4136_/A vssd1 vssd1 vccd1 vccd1 _4469_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4067_ _4067_/A vssd1 vssd1 vccd1 vccd1 _4467_/A sky130_fd_sc_hd__inv_2
XANTENNA__4972__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3018_ _3018_/A vssd1 vssd1 vccd1 vccd1 _3343_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_243_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5279__S _5285_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4378__A2 _4305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4969_ _4969_/A vssd1 vssd1 vccd1 vccd1 _4972_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4783__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_176 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3889__A1 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5446__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4866__B _4872_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_219_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4066__A1 _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_234_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3270__B_N _5478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3498__A _3523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4774__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3437__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4122__A _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_195_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4541__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2727__D _2775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0_0_i_clk_A clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4152__S1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3804__B2 _5469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_280_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4823_ _5605_/Q _4822_/B _4822_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5605_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3017__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4765__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4754_ _5576_/Q _4747_/B _4753_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5576_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _5624_/Q _3597_/X _3598_/X _5608_/Q _3704_/X vssd1 vssd1 vccd1 vccd1 _3705_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4780__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4685_ _5555_/Q _4687_/A vssd1 vssd1 vccd1 vccd1 _4685_/X sky130_fd_sc_hd__or2_1
X_3636_ _5667_/Q _3600_/X _3602_/X _5651_/Q vssd1 vssd1 vccd1 vccd1 _3636_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5469__CLK _5707_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3567_ _5660_/Q _5341_/Q _5343_/Q _5342_/Q vssd1 vssd1 vccd1 vccd1 _3567_/X sky130_fd_sc_hd__and4_1
XANTENNA__4967__A _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5306_ _2760_/Y _5319_/B _5305_/X _4979_/X vssd1 vssd1 vccd1 vccd1 _5745_/D sky130_fd_sc_hd__o211a_1
XFILLER_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_382 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3498_ _3523_/S vssd1 vssd1 vccd1 vccd1 _3517_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__3590__B _4363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5237_ _5331_/A _5458_/Q _5253_/S vssd1 vssd1 vccd1 vccd1 _5238_/A sky130_fd_sc_hd__and3_1
XFILLER_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5168_ _5179_/S _5315_/A vssd1 vssd1 vccd1 vccd1 _5168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4119_ _4229_/A _4231_/S vssd1 vssd1 vccd1 vccd1 _4119_/Y sky130_fd_sc_hd__nand2_1
X_5099_ _4536_/Y _5098_/Y _5087_/Y vssd1 vssd1 vccd1 vccd1 _5109_/A sky130_fd_sc_hd__a21o_1
XFILLER_216_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3111__A _5711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3271__A2 _5461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4756__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4220__A1 _4151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3765__B _4529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4877__A _5628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input43_A i_req_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4287__A1 _4347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3720__S _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5220__B _5225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3021__A _5761_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3956__A _3956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4551__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5611__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2758__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ _4469_/D _4449_/X _4469_/Y _4449_/S vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_327 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3421_ _5390_/Q _3017_/X _3435_/S vssd1 vssd1 vccd1 vccd1 _3422_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_0_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3722__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _2835_/A _5359_/Q _3368_/S vssd1 vssd1 vccd1 vccd1 _3353_/A sky130_fd_sc_hd__mux2_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3283_/A _3283_/B _3283_/C _3283_/D vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__or4_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5692_/Q _4543_/B _5030_/S vssd1 vssd1 vccd1 vccd1 _5023_/A sky130_fd_sc_hd__mux2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2754__B _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4986__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4450__A1 _4449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _5598_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__or2_1
XANTENNA__4738__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2998_ input53/X _5417_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _3001_/B sky130_fd_sc_hd__mux2_1
X_4737_ _5569_/Q _4743_/A vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__or2_1
XFILLER_119_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4668_ _4668_/A vssd1 vssd1 vccd1 vccd1 _4668_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3619_ _3619_/A _3619_/B _4379_/B _3619_/D vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__or4_2
XFILLER_266_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ _5523_/Q _4599_/B vssd1 vssd1 vccd1 vccd1 _4599_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3805__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3713__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_229_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5321__A _5321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2664__B _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4977__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3244__A2 _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5634__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3776__A _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5175__A1_N _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2755__A1 _5568_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3704__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3180__A1 _5650_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3180__B2 _5570_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3016__A _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_85_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5128__A1_N _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4968__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3970_ _5521_/Q _3923_/X _3969_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5521_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4432__A1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4432__B2 _4408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2921_ _5359_/Q _5358_/Q vssd1 vssd1 vccd1 vccd1 _2945_/B sky130_fd_sc_hd__or2_1
XFILLER_188_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3786__A3 _2943_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3686__A _4278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5640_ _5658_/CLK _5640_/D vssd1 vssd1 vccd1 vccd1 _5640_/Q sky130_fd_sc_hd__dfxtp_2
X_2852_ _2852_/A _2852_/B _2852_/C _2852_/D vssd1 vssd1 vccd1 vccd1 _2852_/X sky130_fd_sc_hd__or4_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4196__B1 _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5571_ _5747_/CLK _5571_/D vssd1 vssd1 vccd1 vccd1 _5571_/Q sky130_fd_sc_hd__dfxtp_4
X_2783_ _5613_/Q _2652_/X _2781_/X _2782_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2783_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__2740__D _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4522_ _4635_/A _4522_/B vssd1 vssd1 vccd1 vccd1 _4522_/X sky130_fd_sc_hd__or2_1
XFILLER_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4453_ _4468_/A _4320_/B _4452_/Y _4201_/Y vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__o211a_2
XFILLER_236_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3404_ _3404_/A vssd1 vssd1 vccd1 vccd1 _5381_/D sky130_fd_sc_hd__clkbuf_1
X_4384_ _4384_/A _4384_/B _4384_/C vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__or3_1
XANTENNA__2749__B _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3171__A1 _5632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3335_ _3791_/A _3335_/B _3335_/C vssd1 vssd1 vccd1 vccd1 _3335_/X sky130_fd_sc_hd__or3_1
XANTENNA__5507__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3266_ _3263_/X _3265_/X _5347_/Q vssd1 vssd1 vccd1 vccd1 _3267_/B sky130_fd_sc_hd__o21ai_4
XFILLER_285_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4120__B1 _4307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5005_ _5685_/Q _5339_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _5006_/A sky130_fd_sc_hd__mux2_1
XFILLER_273_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5214__A_N _5225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3197_ _5557_/Q _3131_/X _3194_/X _3196_/X vssd1 vssd1 vccd1 vccd1 _3197_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3360__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4671__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5657__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4423__A1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3226__A2 _3143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3596__A _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_344 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5769_ _5769_/A vssd1 vssd1 vccd1 vccd1 _5769_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3934__A0 _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3162__A1 _5550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4874__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5051__A _5528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2673__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4890__A _5634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4414__A1 _4050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3217__A2 _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_300 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output197_A _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3445__S _3451_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4130__A _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output74_A _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3153__A1 _5661_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3153__B2 _5581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3120_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_267_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4784__B _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _2852_/B _3027_/X _3343_/C vssd1 vssd1 vccd1 vccd1 _3051_/X sky130_fd_sc_hd__a21o_1
XFILLER_208_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2735__D _5634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3208__A2 _3137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _3965_/A _3953_/B vssd1 vssd1 vccd1 vccd1 _3953_/X sky130_fd_sc_hd__or2_1
XFILLER_195_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2904_ _5452_/Q vssd1 vssd1 vccd1 vccd1 _2904_/X sky130_fd_sc_hd__buf_4
XANTENNA__4305__A _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4704__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3884_ _3893_/A _3884_/B vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__and2_1
XFILLER_31_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5623_ _5623_/CLK _5623_/D vssd1 vssd1 vccd1 vccd1 _5623_/Q sky130_fd_sc_hd__dfxtp_1
X_2835_ _2835_/A _2835_/B _2966_/A _2826_/A vssd1 vssd1 vccd1 vccd1 _2852_/C sky130_fd_sc_hd__or4b_1
XANTENNA__4024__B _4024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2719__A1 _5620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5554_ _5747_/CLK _5554_/D vssd1 vssd1 vccd1 vccd1 _5554_/Q sky130_fd_sc_hd__dfxtp_4
X_2766_ _5615_/Q _2652_/A _2764_/X _2765_/X _2686_/A vssd1 vssd1 vccd1 vccd1 _2766_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4959__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2814__S1 _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4505_ _4494_/X _4495_/Y _4504_/Y vssd1 vssd1 vccd1 vccd1 _4507_/A sky130_fd_sc_hd__a21oi_1
X_5485_ _5743_/CLK _5485_/D vssd1 vssd1 vccd1 vccd1 _5485_/Q sky130_fd_sc_hd__dfxtp_4
X_2697_ _2771_/B _2771_/A _2806_/A _5638_/Q vssd1 vssd1 vccd1 vccd1 _2697_/X sky130_fd_sc_hd__and4b_1
XFILLER_144_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4436_ _4483_/A _4421_/Y _4422_/X _4435_/Y vssd1 vssd1 vccd1 vccd1 _4484_/C sky130_fd_sc_hd__a31o_1
XFILLER_144_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4341__B1 _3555_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4367_ _4386_/A _4386_/B _4386_/C vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__a21oi_1
XFILLER_258_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3695__A2 _4278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3318_ _3318_/A _5241_/B _3318_/C vssd1 vssd1 vccd1 vccd1 _3791_/D sky130_fd_sc_hd__or3_2
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4298_ _4090_/D _4296_/Y _4297_/Y vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__a21o_1
XFILLER_246_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3249_ _5508_/Q _5478_/Q _3860_/B vssd1 vssd1 vccd1 vccd1 _3250_/D sky130_fd_sc_hd__and3_1
XANTENNA__2926__C _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3103__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2645__D _5611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4885__A _5632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_249_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_201 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_264_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output112_A _5559_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4938__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2852__B _2852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4125__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3610__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5352__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput106 _5766_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[6] sky130_fd_sc_hd__buf_2
XFILLER_217_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput117 _5549_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[1] sky130_fd_sc_hd__buf_2
Xoutput128 _5741_/Q vssd1 vssd1 vccd1 vccd1 o_icache_flush sky130_fd_sc_hd__buf_2
Xoutput139 _5694_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5270_ _5733_/Q _5768_/A _5285_/S vssd1 vssd1 vccd1 vccd1 _5271_/B sky130_fd_sc_hd__mux2_1
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4221_ _4221_/A _4221_/B vssd1 vssd1 vccd1 vccd1 _4221_/X sky130_fd_sc_hd__or2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4795__A _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4152_ _4148_/X _4149_/X _4150_/X _4151_/X _4272_/S _4146_/A vssd1 vssd1 vccd1 vccd1
+ _4153_/B sky130_fd_sc_hd__mux4_1
XFILLER_233_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3103_ _5707_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3104_/A sky130_fd_sc_hd__and2_1
XFILLER_233_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4083_ _4083_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__or2_2
XFILLER_55_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4626__A1 _4457_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2746__C _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3034_ _5763_/A _3010_/X _3032_/Y _3033_/X _3016_/X vssd1 vssd1 vccd1 vccd1 _3034_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4985_ _4985_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4985_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3936_ _3948_/B _3934_/X _3935_/Y _3965_/A vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__a211o_1
XFILLER_258_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_258_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3867_ _3893_/A _3867_/B vssd1 vssd1 vccd1 vccd1 _3868_/A sky130_fd_sc_hd__and2_1
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3874__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5606_ _5654_/CLK _5606_/D vssd1 vssd1 vccd1 vccd1 _5606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2818_ input6/X vssd1 vssd1 vccd1 vccd1 _2818_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3798_ _3798_/A vssd1 vssd1 vccd1 vccd1 _5467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5537_ _5756_/CLK _5537_/D vssd1 vssd1 vccd1 vccd1 _5765_/A sky130_fd_sc_hd__dfxtp_4
X_2749_ _5553_/Q _2791_/B vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__or2_1
XFILLER_105_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_274_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5106__A2 _5125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5468_ _5707_/CLK _5468_/D vssd1 vssd1 vccd1 vccd1 _5468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_132_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4419_ _4419_/A _4419_/B vssd1 vssd1 vccd1 vccd1 _4420_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3668__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3813__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5399_ _5492_/CLK _5399_/D vssd1 vssd1 vccd1 vccd1 _5399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_246_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4078__C1 _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2656__C _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5042__A1 _4617_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5375__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 i_mem_data[6] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_314 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3356__A1 _5361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4553__B1 _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_123_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3659__A2 _3605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4721__A1_N input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_218 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4608__A1 _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5718__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2863__A _5331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3678__B _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5033__A1 _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_233_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _4658_/X _4761_/Y _4768_/X _4769_/X vssd1 vssd1 vccd1 vccd1 _5582_/D sky130_fd_sc_hd__o211a_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4241__C1 _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3721_ _5669_/Q _3600_/A _3602_/A _5653_/Q vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2635__C_N _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3652_ _5614_/Q _3597_/X _3598_/X _5598_/Q _3651_/X vssd1 vssd1 vccd1 vccd1 _3652_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3347__A1 _5357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3583_ _5482_/Q _5321_/A _3588_/S vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__mux2_4
XFILLER_228_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5322_ _5753_/Q _5295_/X _5321_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5753_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5253_ _5728_/Q _5763_/A _5253_/S vssd1 vssd1 vccd1 vccd1 _5254_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4847__A1 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4204_ _4121_/B _4203_/X _4276_/A vssd1 vssd1 vccd1 vccd1 _4271_/B sky130_fd_sc_hd__mux2_2
XANTENNA__3860__C _5472_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5184_ _5752_/Q _3840_/X _5183_/X vssd1 vssd1 vccd1 vccd1 _5184_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2757__B _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4135_ _4274_/A _4139_/B vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_228_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4066_ _4348_/A _4088_/B _4065_/X vssd1 vssd1 vccd1 vccd1 _4066_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4972__B _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3869__A _3908_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3017_ _4527_/C _3010_/X _3013_/X _3015_/Y _3016_/X vssd1 vssd1 vccd1 vccd1 _3017_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5024__A1 _4499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_196_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4968_ _4684_/X _4949_/Y _4967_/X _4957_/X vssd1 vssd1 vccd1 vccd1 _5667_/D sky130_fd_sc_hd__o211a_1
XFILLER_196_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3919_ _3919_/A vssd1 vssd1 vccd1 vccd1 _3919_/X sky130_fd_sc_hd__buf_4
X_4899_ _4974_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4899_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3338__A1 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4535__B1 _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3109__A _5710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_21 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_219_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_239 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_270_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3779__A _5460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3274__B1 _3851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3577__A1 _5558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3577__B2 _2702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3329__A1 _5347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4526__B1 _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4829__A1 _5608_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_214_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5540__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3689__A _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4462__C1 _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5690__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_240_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4822_ _4972_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_376 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4753_ _4978_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4753_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3704_ _5672_/Q _3600_/X _3602_/X _5656_/Q vssd1 vssd1 vccd1 vccd1 _3704_/X sky130_fd_sc_hd__a22o_1
X_4684_ _4684_/A vssd1 vssd1 vccd1 vccd1 _4684_/X sky130_fd_sc_hd__buf_4
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3635_ _4303_/A _3635_/B vssd1 vssd1 vccd1 vccd1 _3635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3566_ _3601_/C _3599_/B _3601_/B vssd1 vssd1 vccd1 vccd1 _3606_/A sky130_fd_sc_hd__nor3_4
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5305_ _5745_/Q _5327_/B vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__or2_1
XFILLER_255_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2768__A _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3497_ _3497_/A vssd1 vssd1 vccd1 vccd1 _5428_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5144__A _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_142_394 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5236_ _5236_/A vssd1 vssd1 vccd1 vccd1 _5721_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4150__D1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4983__A _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5167_ _4503_/A _5166_/Y _5200_/B vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__mux2_1
XFILLER_271_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4118_ _4302_/S _4118_/B vssd1 vssd1 vccd1 vccd1 _4221_/B sky130_fd_sc_hd__and2_1
XFILLER_83_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5098_ _5093_/X _5097_/X _5219_/S vssd1 vssd1 vccd1 vccd1 _5098_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_204_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3599__A _3601_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4049_ _4050_/A _4415_/A vssd1 vssd1 vccd1 vccd1 _4052_/A sky130_fd_sc_hd__or2_2
XFILLER_17_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xcore_218 vssd1 vssd1 vccd1 vccd1 core_218/HI o_mem_addr[15] sky130_fd_sc_hd__conb_1
XFILLER_271_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3111__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4205__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5319__A _5319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5413__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4508__B1 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4877__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3731__A1 _5556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5563__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4287__A2 _4199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input36_A i_req_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_181_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4995__A0 _5680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4133__A _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3970__A1 _5521_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_283 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3420_ _3420_/A vssd1 vssd1 vccd1 vccd1 _5389_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3722__A1 _5621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3351_ _3351_/A vssd1 vssd1 vccd1 vccd1 _5358_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3722__B2 _5605_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_225_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3282_ _3802_/A _3282_/B vssd1 vssd1 vccd1 vccd1 _3283_/D sky130_fd_sc_hd__or2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A vssd1 vssd1 vccd1 vccd1 _5691_/D sky130_fd_sc_hd__clkbuf_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater214 _5769_/A vssd1 vssd1 vccd1 vccd1 _4590_/B sky130_fd_sc_hd__buf_6
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2754__C _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4027__B _4027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5436__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4805_ _4653_/X _4799_/Y _4804_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _5597_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3358__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2997_ input54/X _5418_/Q _3000_/S vssd1 vssd1 vccd1 vccd1 _3001_/A sky130_fd_sc_hd__mux2_1
X_4736_ _4668_/X _4724_/Y _4735_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5568_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4667_ _5708_/Q _4666_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__mux2_2
XANTENNA__5586__CLK _5680_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4978__A _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3618_ _5480_/Q _3532_/X _3577_/X _3549_/A _3549_/B vssd1 vssd1 vccd1 vccd1 _3619_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4697__B _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4598_ _5770_/A _4511_/X _3919_/A _4597_/X vssd1 vssd1 vccd1 vccd1 _5542_/D sky130_fd_sc_hd__o211a_1
XFILLER_122_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_134_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3713__A1 _5626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3713__B2 _5610_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3549_ _3549_/A _3549_/B vssd1 vssd1 vccd1 vccd1 _3550_/A sky130_fd_sc_hd__or2_1
XFILLER_282_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5219_ _5215_/Y _5218_/X _5219_/S vssd1 vssd1 vccd1 vccd1 _5225_/A sky130_fd_sc_hd__mux2_2
XFILLER_276_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5218__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2664__C _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4652__S _4690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3401__A0 _2852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2755__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3952__A1 _5307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_87 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4888__A _5633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3704__A1 _5672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3704__B2 _5656_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_302 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3180__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4665__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4128__A _4128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5459__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3032__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_224 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_i_clk_A clkbuf_2_1_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2920_ _5242_/S vssd1 vssd1 vccd1 vccd1 _3780_/A sky130_fd_sc_hd__buf_4
XANTENNA__3640__B1 _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2994__A2 _2835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2851_ _2851_/A _2851_/B _2851_/C vssd1 vssd1 vccd1 vccd1 _2852_/D sky130_fd_sc_hd__or3_1
X_5570_ _5747_/CLK _5570_/D vssd1 vssd1 vccd1 vccd1 _5570_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2782_ _2757_/D _2782_/B _2782_/C _5597_/Q vssd1 vssd1 vccd1 vccd1 _2782_/X sky130_fd_sc_hd__and4b_1
XFILLER_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4521_ _4533_/C _4511_/X _3919_/X _4520_/X vssd1 vssd1 vccd1 vccd1 _5533_/D sky130_fd_sc_hd__o211a_1
XFILLER_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4452_ _4300_/S _4450_/X _4451_/X vssd1 vssd1 vccd1 vccd1 _4452_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3403_ _2852_/B _5381_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3404_/A sky130_fd_sc_hd__mux2_1
X_4383_ _4471_/S _4220_/X _4372_/Y _4376_/X _4382_/X vssd1 vssd1 vccd1 vccd1 _4384_/C
+ sky130_fd_sc_hd__a311o_2
XFILLER_124_180 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3171__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3334_ _5351_/Q _3293_/X _3330_/X _5365_/Q vssd1 vssd1 vccd1 vccd1 _5351_/D sky130_fd_sc_hd__a22o_1
XFILLER_252_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2782__A_N _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3265_/A _3265_/B _5348_/Q _3265_/D vssd1 vssd1 vccd1 vccd1 _3265_/X sky130_fd_sc_hd__and4_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4120__A1 _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5004_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_273_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3196_ _5637_/Q _3143_/X _3145_/X _3195_/X vssd1 vssd1 vccd1 vccd1 _3196_/X sky130_fd_sc_hd__a211o_1
XFILLER_252_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4671__A2 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4038__A _4192_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4423__A2 _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2985__A2 _2840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4187__A1 _4372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5768_ _5768_/A vssd1 vssd1 vccd1 vccd1 _5768_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4719_ _5562_/Q _4697_/A _4717_/Y _4718_/X vssd1 vssd1 vccd1 vccd1 _5562_/D sky130_fd_sc_hd__o211a_1
X_5699_ _5724_/CLK _5699_/D vssd1 vssd1 vccd1 vccd1 _5699_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3816__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3698__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3162__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5601__CLK _5680_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_257_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5051__B _5051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2673__A1 _5640_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2673__B2 _5672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_371 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4890__B _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2691__A _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5751__CLK _5756_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3622__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4178__A1 _4140_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4130__B _4130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3027__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3153__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output67_A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3461__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_255_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3050_ _3085_/A _3050_/B vssd1 vssd1 vccd1 vccd1 _3050_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5599__D _5599_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_263_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3952_ _3951_/X _5307_/A _3984_/S vssd1 vssd1 vccd1 vccd1 _3953_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2903_ _2903_/A vssd1 vssd1 vccd1 vccd1 _5453_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4305__B _4305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3883_ _5499_/Q _5311_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3884_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5622_ _5654_/CLK _5622_/D vssd1 vssd1 vccd1 vccd1 _5622_/Q sky130_fd_sc_hd__dfxtp_1
X_2834_ input42/X _5436_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2966_/A sky130_fd_sc_hd__mux2_2
XANTENNA__2719__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3916__A1 _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5553_ _5747_/CLK _5553_/D vssd1 vssd1 vccd1 vccd1 _5553_/Q sky130_fd_sc_hd__dfxtp_4
X_2765_ _5344_/Q _5346_/Q _5345_/Q _5599_/Q vssd1 vssd1 vccd1 vccd1 _2765_/X sky130_fd_sc_hd__and4b_1
XFILLER_191_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4504_ _4504_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4504_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_191_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5484_ _5722_/CLK _5484_/D vssd1 vssd1 vccd1 vccd1 _5484_/Q sky130_fd_sc_hd__dfxtp_4
X_2696_ _2782_/B vssd1 vssd1 vccd1 vccd1 _2771_/A sky130_fd_sc_hd__buf_4
X_4435_ _4372_/B _4429_/X _4434_/X vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4341__A1 _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4366_ _4377_/A _4364_/X _4365_/Y vssd1 vssd1 vccd1 vccd1 _4384_/A sky130_fd_sc_hd__o21a_1
XANTENNA__5624__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3317_ _3317_/A _3317_/B vssd1 vssd1 vccd1 vccd1 _3319_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4297_ _4090_/D _4296_/Y _5453_/Q vssd1 vssd1 vccd1 vccd1 _4297_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3371__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3248_ _5508_/Q _3248_/B vssd1 vssd1 vccd1 vccd1 _3248_/X sky130_fd_sc_hd__xor2_1
XANTENNA__2926__D _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3179_ _5602_/Q _3133_/X _3135_/X _5618_/Q _3178_/X vssd1 vssd1 vccd1 vccd1 _3179_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3852__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_213 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3604__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4580__A1 _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_200 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4885__B _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5001__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5237__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4571__A1 _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5647__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 _5767_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[7] sky130_fd_sc_hd__buf_2
Xoutput118 _5550_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[2] sky130_fd_sc_hd__buf_2
Xoutput129 _5689_/Q vssd1 vssd1 vccd1 vccd1 o_mem_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_126_275 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4220_ _4248_/C _4151_/X _4154_/X _4150_/X _4136_/A _4449_/S vssd1 vssd1 vccd1 vccd1
+ _4220_/X sky130_fd_sc_hd__mux4_2
XANTENNA__4795__B _4797_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4151_ _4132_/A _4083_/B _3613_/X _4469_/C _4469_/B vssd1 vssd1 vccd1 vccd1 _4151_/X
+ sky130_fd_sc_hd__o2111a_2
XFILLER_228_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3102_ _3102_/A vssd1 vssd1 vccd1 vccd1 _3102_/X sky130_fd_sc_hd__clkbuf_1
X_4082_ _4281_/A _4280_/B _4080_/X _4081_/Y vssd1 vssd1 vccd1 vccd1 _4240_/S sky130_fd_sc_hd__a211o_2
XFILLER_255_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2746__D _5585_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3033_ _2845_/B _3027_/X _3343_/C vssd1 vssd1 vccd1 vccd1 _3033_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3834__A0 _5484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _5674_/Q _4972_/B _4983_/Y _4979_/X vssd1 vssd1 vccd1 vccd1 _5674_/D sky130_fd_sc_hd__o211a_1
X_3935_ _3935_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _3935_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3062__A1 _2850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3866_ _5492_/Q _5067_/B _3908_/B vssd1 vssd1 vccd1 vccd1 _3867_/B sky130_fd_sc_hd__mux2_1
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5605_ _5674_/CLK _5605_/D vssd1 vssd1 vccd1 vccd1 _5605_/Q sky130_fd_sc_hd__dfxtp_4
X_2817_ _5352_/Q _2805_/X _2808_/X _2816_/X vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3366__S _3368_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3797_ _5467_/Q _3310_/B _3813_/S vssd1 vssd1 vccd1 vccd1 _3798_/A sky130_fd_sc_hd__mux2_1
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5536_ _5665_/CLK _5536_/D vssd1 vssd1 vccd1 vccd1 _5764_/A sky130_fd_sc_hd__dfxtp_4
X_2748_ _5617_/Q _2652_/A _2746_/X _2747_/X _2686_/X vssd1 vssd1 vccd1 vccd1 _2748_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_117_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5467_ _5721_/CLK _5467_/D vssd1 vssd1 vccd1 vccd1 _5467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2679_ _5575_/Q _2644_/X _2664_/X _5607_/Q vssd1 vssd1 vccd1 vccd1 _2679_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3890__A _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4314__B2 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4418_ _4418_/A vssd1 vssd1 vccd1 vccd1 _4419_/B sky130_fd_sc_hd__inv_2
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5398_ _5492_/CLK _5398_/D vssd1 vssd1 vccd1 vccd1 _5398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4865__A2 _4859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4349_ _4348_/B _4348_/C _4348_/A vssd1 vssd1 vccd1 vccd1 _4350_/C sky130_fd_sc_hd__o21ai_1
XFILLER_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4173__S0 _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_261_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__C1 _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5057__A _5460_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_359 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4553__A1 _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4608__A2 _4581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3816__A0 _5475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3720_ _3711_/X _4454_/C _4454_/B vssd1 vssd1 vccd1 vccd1 _4182_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4792__A1 _5592_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3651_ _5662_/Q _3600_/A _3602_/A _5646_/Q vssd1 vssd1 vccd1 vccd1 _3651_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_146_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4544__A1 _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3582_ _5477_/Q _3532_/X _3579_/X _4027_/A _4027_/B vssd1 vssd1 vccd1 vccd1 _3619_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5321_ _5321_/A _5325_/B vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__or2_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5252_ _5252_/A vssd1 vssd1 vccd1 vccd1 _5727_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4847__A2 _4836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4203_ _3710_/X _3740_/X _3747_/X _3726_/Y _4274_/A _4231_/S vssd1 vssd1 vccd1 vccd1
+ _4203_/X sky130_fd_sc_hd__mux4_2
XANTENNA__2858__A1 _2830_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5183_ _5523_/Q _3932_/B _3864_/C _5503_/Q vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2757__C _5648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4134_ _5454_/Q _4301_/S vssd1 vssd1 vccd1 vccd1 _4139_/B sky130_fd_sc_hd__nand2_2
XFILLER_95_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _4348_/A _4088_/B _4087_/B _4087_/A vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__o211a_1
XFILLER_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3807__A0 _5471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3016_ _3016_/A vssd1 vssd1 vccd1 vccd1 _3016_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4967_ _5667_/Q _4969_/A vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__or2_1
XFILLER_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4783__A1 _5588_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3918_ _3935_/A _3918_/B vssd1 vssd1 vccd1 vccd1 _3918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4898_ _5637_/Q _4897_/B _4897_/Y _4886_/X vssd1 vssd1 vccd1 vccd1 _5637_/D sky130_fd_sc_hd__o211a_1
XFILLER_137_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3991__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3849_ _3843_/X _3846_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _5487_/D sky130_fd_sc_hd__o21a_1
XFILLER_137_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3338__A2 _3318_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4535__A1 _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3109__B _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5519_ _5740_/CLK _5519_/D vssd1 vssd1 vccd1 vccd1 _5519_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3824__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2667__C _2747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5342__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_66 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_234_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3274__A1 _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__A _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3577__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4774__A1 _4668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3329__A2 _3780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4526__A1 _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4829__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4137__S0 _4447_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_233_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4821_ _5604_/Q _4822_/B _4820_/Y _4815_/X vssd1 vssd1 vccd1 vccd1 _5604_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3017__A1 _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4214__B1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4752_ _5575_/Q _4747_/B _4751_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5575_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4765__A1 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3703_ _3747_/A _3747_/B _3703_/C vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__or3_1
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4683_ _5711_/Q _4682_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3634_ _4232_/B _4063_/A _4302_/S vssd1 vssd1 vccd1 vccd1 _3635_/B sky130_fd_sc_hd__mux2_1
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3565_ _5341_/Q _3601_/B _5343_/Q vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__nor3b_4
XFILLER_255_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5304_ _2768_/Y _5319_/B _5303_/X _4979_/X vssd1 vssd1 vccd1 vccd1 _5744_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3496_ _5428_/Q input33/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3497_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_17_i_clk_A clkbuf_2_3_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5365__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5144__B _5311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5235_ _5463_/Q _5721_/Q _5235_/S vssd1 vssd1 vccd1 vccd1 _5236_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5166_ _5166_/A _5166_/B vssd1 vssd1 vccd1 vccd1 _5166_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4983__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4117_ _3732_/A _4418_/A _4231_/S vssd1 vssd1 vccd1 vccd1 _4221_/A sky130_fd_sc_hd__a21oi_1
XFILLER_244_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5097_ _5094_/X _5095_/X _5096_/X _5071_/B vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__o31a_1
XFILLER_216_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3599__B _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4048_ _4168_/A _4389_/A _4046_/Y _4103_/A vssd1 vssd1 vccd1 vccd1 _4055_/B sky130_fd_sc_hd__o211a_2
XFILLER_204_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcore_219 vssd1 vssd1 vccd1 vccd1 o_req_active core_219/LO sky130_fd_sc_hd__conb_1
XFILLER_71_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_231_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_221 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_271_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4205__B1 _4130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4756__A1 _5577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_149_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4220__A3 _4150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2767__B1 _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4508__A1 _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5708__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_136 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3731__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4692__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2694__A _2782_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A i_req_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_357 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_207_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4444__B1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_288 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5388__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2869__A _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3183__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5245__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4380__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3722__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3350_ _2826_/A _3277_/A _3368_/S vssd1 vssd1 vccd1 vccd1 _3351_/A sky130_fd_sc_hd__mux2_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3281_/A _3281_/B _3281_/C vssd1 vssd1 vccd1 vccd1 _3282_/B sky130_fd_sc_hd__and3_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5020_ _5691_/Q _4537_/B _5030_/S vssd1 vssd1 vccd1 vccd1 _5021_/A sky130_fd_sc_hd__mux2_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4683__A0 _5711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater215 _5539_/Q vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__buf_6
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2754__D _5632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4986__A1 _5675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4804_ _5597_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__or2_1
XFILLER_221_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4738__A1 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4324__A _5453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2996_ _2962_/Y _2850_/C _2850_/D _3084_/A _2995_/X vssd1 vssd1 vccd1 vccd1 _2996_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4735_ _5568_/Q _4743_/A vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__or2_1
XFILLER_174_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4666_ input10/X input17/X _4682_/S vssd1 vssd1 vccd1 vccd1 _4666_/X sky130_fd_sc_hd__mux2_1
XFILLER_266_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4978__B _4985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3617_ _3617_/A vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3374__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4597_ _4532_/X _4604_/B _4592_/X _4596_/Y _4529_/X vssd1 vssd1 vccd1 vccd1 _4597_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3174__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3713__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3548_ _2744_/X _2745_/X _2748_/X _2749_/X _3528_/A vssd1 vssd1 vccd1 vccd1 _3549_/B
+ sky130_fd_sc_hd__o311a_2
XFILLER_282_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_54 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3479_ _3479_/A vssd1 vssd1 vccd1 vccd1 _5419_/D sky130_fd_sc_hd__clkbuf_1
X_5218_ _5774_/A _5193_/B _5217_/Y _5196_/A vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5149_ _5520_/Q _3932_/B _3864_/C _5500_/Q vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__a22o_1
XFILLER_244_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4426__B1 _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4977__A1 _5671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_224 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4234__A _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3937__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5530__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4888__B _4894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3165__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3704__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5680__CLK _5680_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_235_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4128__B _4128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4968__A1 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3640__B2 _5555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3459__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2850_ _2850_/A _2850_/B _2850_/C _2850_/D vssd1 vssd1 vccd1 vccd1 _2851_/C sky130_fd_sc_hd__or4_1
X_2781_ _2757_/D _2782_/C _2782_/B _5565_/Q vssd1 vssd1 vccd1 vccd1 _2781_/X sky130_fd_sc_hd__and4bb_1
X_4520_ _4585_/A _4515_/Y _4519_/X vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4451_ _4471_/S _4395_/X _4372_/A vssd1 vssd1 vccd1 vccd1 _4451_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5145__A1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3156__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3402_ _3402_/A vssd1 vssd1 vccd1 vccd1 _5380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4382_ _5449_/Q _4377_/Y _4378_/Y _3678_/Y _4381_/X vssd1 vssd1 vccd1 vccd1 _4382_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3333_ _5350_/Q _3293_/X _3330_/X _5366_/Q vssd1 vssd1 vccd1 vccd1 _5350_/D sky130_fd_sc_hd__a22o_1
XFILLER_285_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3264_ _5531_/Q _5532_/Q _5351_/Q vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4656__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5684_/Q _5338_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__mux2_1
XFILLER_285_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3195_ _5653_/Q _3147_/X _3149_/X _5573_/Q vssd1 vssd1 vccd1 vccd1 _3195_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2765__C _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5403__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_121_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3631__A1 _5552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5553__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4054__A _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4187__A2 _4175_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4989__A _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5767_ _5767_/A vssd1 vssd1 vccd1 vccd1 _5767_/X sky130_fd_sc_hd__clkbuf_1
X_2979_ _5391_/Q vssd1 vssd1 vccd1 vccd1 _2979_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3893__A _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4718_ _5331_/A vssd1 vssd1 vccd1 vccd1 _4718_/X sky130_fd_sc_hd__clkbuf_4
X_5698_ _5724_/CLK _5698_/D vssd1 vssd1 vccd1 vccd1 _5698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4649_ _5548_/Q _4722_/A vssd1 vssd1 vccd1 vccd1 _4649_/X sky130_fd_sc_hd__or2_1
XANTENNA__4501__B _4501_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3698__A1 _5625_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3698__B2 _5609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2659__D _5610_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3832__S _3834_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4229__A _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3133__A _3133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2675__C _5656_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2673__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_383 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3622__A1 _5665_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3622__B2 _5649_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4899__A _4974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4178__A2 _4141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2911__S _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_220 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3308__A _3308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5426__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4638__B1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4139__A _4229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_208_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5576__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3951_ _5765_/A _5730_/Q _3988_/S vssd1 vssd1 vccd1 vccd1 _3951_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2902_ _4483_/A _2901_/X _3337_/B vssd1 vssd1 vccd1 vccd1 _2903_/A sky130_fd_sc_hd__mux2_1
X_3882_ _5498_/Q _3874_/B _3881_/Y _3848_/X vssd1 vssd1 vccd1 vccd1 _5498_/D sky130_fd_sc_hd__o211a_1
X_5621_ _5623_/CLK _5621_/D vssd1 vssd1 vccd1 vccd1 _5621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2833_ input44/X _5438_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2835_/B sky130_fd_sc_hd__mux2_2
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_251 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5552_ _5667_/CLK _5552_/D vssd1 vssd1 vccd1 vccd1 _5552_/Q sky130_fd_sc_hd__dfxtp_4
X_2764_ _5344_/Q _5345_/Q _5346_/Q _5567_/Q vssd1 vssd1 vccd1 vccd1 _2764_/X sky130_fd_sc_hd__and4bb_1
XFILLER_191_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4503_ _4503_/A _5156_/A vssd1 vssd1 vccd1 vccd1 _4504_/B sky130_fd_sc_hd__xnor2_1
XFILLER_191_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483_ _5722_/CLK _5483_/D vssd1 vssd1 vccd1 vccd1 _5483_/Q sky130_fd_sc_hd__dfxtp_4
X_2695_ _2806_/A _2727_/C _2771_/B _5606_/Q vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__and4b_1
XFILLER_247_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4434_ _4454_/D _4307_/X _4433_/Y vssd1 vssd1 vccd1 vccd1 _4434_/X sky130_fd_sc_hd__o21a_1
X_4365_ _4377_/A _4364_/X _4322_/A vssd1 vssd1 vccd1 vccd1 _4365_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3316_ _3599_/B _5486_/D _3315_/X vssd1 vssd1 vccd1 vccd1 _5343_/D sky130_fd_sc_hd__o21a_1
XFILLER_263_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4296_ _4323_/A _4070_/B _4070_/A vssd1 vssd1 vccd1 vccd1 _4296_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__4049__A _4050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3247_ _5510_/Q _3843_/B vssd1 vssd1 vccd1 vccd1 _3248_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3301__B1 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3178_ _5666_/Q _3137_/X _3139_/X _5586_/Q vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3852__A1 _3893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3604__A1 _5627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3604__B2 _5611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3368__A0 _3001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4565__C1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5449__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2967__A _2967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5599__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_252_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input11_A i_mem_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3310__B _3310_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5237__B _5458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4571__A2 _4496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput108 _5768_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[8] sky130_fd_sc_hd__buf_2
Xoutput119 _5551_/Q vssd1 vssd1 vccd1 vccd1 dbg_r0[3] sky130_fd_sc_hd__buf_2
XFILLER_126_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2877__A _3308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4150_ _4132_/A _4024_/B _3613_/X _4469_/C _4469_/B vssd1 vssd1 vccd1 vccd1 _4150_/X
+ sky130_fd_sc_hd__o2111a_2
Xoutput90 _3182_/X vssd1 vssd1 vccd1 vccd1 dbg_out[6] sky130_fd_sc_hd__buf_2
X_3101_ _5706_/Q _3113_/S vssd1 vssd1 vccd1 vccd1 _3102_/A sky130_fd_sc_hd__and2_1
XFILLER_228_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4081_ _4083_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _4081_/Y sky130_fd_sc_hd__xnor2_1
X_3032_ _3085_/A _3039_/C _3031_/X vssd1 vssd1 vccd1 vccd1 _3032_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_95_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4983_ _4983_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4983_/Y sky130_fd_sc_hd__nand2_1
XFILLER_211_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_211_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3934_ _4533_/C _5726_/Q _5329_/A vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3865_ _3905_/S vssd1 vssd1 vccd1 vccd1 _3908_/B sky130_fd_sc_hd__clkbuf_4
X_2816_ _3601_/C _2812_/X _2815_/X _5353_/Q vssd1 vssd1 vccd1 vccd1 _2816_/X sky130_fd_sc_hd__o211a_1
X_5604_ _5659_/CLK _5604_/D vssd1 vssd1 vccd1 vccd1 _5604_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_176_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3796_ _5466_/Q _3795_/A _3795_/Y _3277_/A vssd1 vssd1 vccd1 vccd1 _5466_/D sky130_fd_sc_hd__a22o_1
XFILLER_164_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5535_ _5665_/CLK _5535_/D vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__dfxtp_4
X_2747_ _2733_/A _2747_/B _5649_/Q _2747_/D vssd1 vssd1 vccd1 vccd1 _2747_/X sky130_fd_sc_hd__and4b_1
XFILLER_274_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5466_ _5692_/CLK _5466_/D vssd1 vssd1 vccd1 vccd1 _5466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2678_ _2678_/A vssd1 vssd1 vccd1 vccd1 _5321_/A sky130_fd_sc_hd__buf_4
XFILLER_172_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ _4441_/A _4441_/B _4171_/B _4060_/B _4416_/Y vssd1 vssd1 vccd1 vccd1 _4422_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_278_217 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5741__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3382__S _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5397_ _5492_/CLK _5397_/D vssd1 vssd1 vccd1 vccd1 _5397_/Q sky130_fd_sc_hd__dfxtp_1
X_4348_ _4348_/A _4348_/B _4348_/C vssd1 vssd1 vccd1 vccd1 _4350_/B sky130_fd_sc_hd__or3_1
XANTENNA_input3_A dbg_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4279_ _4014_/X _4279_/B _4350_/A vssd1 vssd1 vccd1 vccd1 _4279_/X sky130_fd_sc_hd__and3b_1
XANTENNA__4078__A1 _3572_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_246_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2645__A_N _2747_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4173__S1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3038__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4538__C1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_108_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_163_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4710__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_277_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3029__C1 _3016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4241__A1 _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5614__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4241__B2 _4024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4792__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3467__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5248__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3650_ _4454_/A _3650_/B vssd1 vssd1 vccd1 vccd1 _3650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3581_ _5554_/Q _2720_/B _2738_/X _2741_/X _3528_/A vssd1 vssd1 vccd1 vccd1 _4027_/B
+ sky130_fd_sc_hd__o221a_2
XANTENNA__4544__A2 _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _5752_/Q _5295_/X _5319_/X _4487_/X vssd1 vssd1 vccd1 vccd1 _5752_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5251_ _5261_/A _5251_/B vssd1 vssd1 vccd1 vccd1 _5252_/A sky130_fd_sc_hd__and2_1
X_4202_ _4428_/A _4200_/X _4201_/Y vssd1 vssd1 vccd1 vccd1 _4202_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2668__A_N _2733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5182_ _5182_/A _5177_/B vssd1 vssd1 vccd1 vccd1 _5192_/A sky130_fd_sc_hd__or2b_1
XFILLER_244_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2757__D _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4133_ _4373_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4133_/X sky130_fd_sc_hd__and2_1
XFILLER_228_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4064_ _4024_/B _4326_/A vssd1 vssd1 vccd1 vccd1 _4087_/B sky130_fd_sc_hd__nand2b_1
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3015_ _5390_/Q _3085_/A vssd1 vssd1 vccd1 vccd1 _3015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_243_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2773__C _2789_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4480__A1 _4482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3231__A _3419_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_13_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4966_ _4679_/X _4949_/Y _4965_/X _4957_/X vssd1 vssd1 vccd1 vccd1 _5666_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3586__A3 _2719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3917_ _3843_/B _3916_/X _4987_/A vssd1 vssd1 vccd1 vccd1 _5510_/D sky130_fd_sc_hd__a21o_1
XANTENNA__4783__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3377__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4897_ _4972_/A _4897_/B vssd1 vssd1 vccd1 vccd1 _4897_/Y sky130_fd_sc_hd__nand2_1
X_3848_ _4979_/A vssd1 vssd1 vccd1 vccd1 _3848_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3338__A3 _3310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4535__A2 _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3779_ _5460_/Q vssd1 vssd1 vccd1 vccd1 _5196_/A sky130_fd_sc_hd__buf_4
XANTENNA__3743__B1 _3608_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4940__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5518_ _5741_/CLK _5518_/D vssd1 vssd1 vccd1 vccd1 _5518_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5449_ _5692_/CLK _5449_/D vssd1 vssd1 vccd1 vccd1 _5449_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_160_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4299__A1 _4127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2667__D _5593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4774__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4526__A2 _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3734__B1 _3602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5007__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3750__S _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4137__S1 _4469_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2874__B _5363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3986__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4820_ _4970_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4214__A1 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4976_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4751_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4765__A2 _4761_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2776__A1 _2771_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3702_ _4415_/A vssd1 vssd1 vccd1 vccd1 _3703_/C sky130_fd_sc_hd__inv_2
X_4682_ input13/X input20/X _4682_/S vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3633_ _3633_/A vssd1 vssd1 vccd1 vccd1 _4302_/S sky130_fd_sc_hd__clkbuf_4
X_3564_ _5628_/Q _3605_/A _3598_/A _5596_/Q vssd1 vssd1 vccd1 vccd1 _3564_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4610__A _4626_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4922__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_255_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5303_ _5744_/Q _5327_/B vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__or2_1
XFILLER_255_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3495_ _3495_/A vssd1 vssd1 vccd1 vccd1 _5427_/D sky130_fd_sc_hd__clkbuf_1
X_5234_ _5234_/A vssd1 vssd1 vccd1 vccd1 _5719_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4150__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5165_ _5161_/Y _5164_/X _5219_/S vssd1 vssd1 vccd1 vccd1 _5166_/B sky130_fd_sc_hd__mux2_1
XFILLER_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _4116_/A _4271_/A vssd1 vssd1 vccd1 vccd1 _4454_/D sky130_fd_sc_hd__or2_4
XFILLER_256_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _5495_/Q _5082_/B _5055_/X _5491_/Q vssd1 vssd1 vccd1 vccd1 _5096_/X sky130_fd_sc_hd__a22o_1
XFILLER_216_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4047_ _4379_/B _4379_/C vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__or2_1
XANTENNA__3599__C _3601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4057__A _5453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4205__A1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4205__B2 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4756__A2 _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4949_ _5687_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4949_/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2767__B2 _5551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4508__A2 _4485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3716__B1 _3713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3192__A1 _5556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3136__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4141__B1 _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_369 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4444__A1 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3955__A0 _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3707__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3183__A1 _5667_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4380__B1 _4379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3183__B2 _5587_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3046__A _3085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _2938_/B _2923_/B _3799_/A vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__a21oi_1
XFILLER_225_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4576__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2885__A _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3480__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5261__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater216 _5764_/A vssd1 vssd1 vccd1 vccd1 _4552_/B sky130_fd_sc_hd__buf_6
XFILLER_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_238_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_306 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4435__A1 _4372_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4986__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2824__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4803_ _4646_/X _4799_/Y _4802_/X _4791_/X vssd1 vssd1 vccd1 vccd1 _5596_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_221_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4738__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2995_ _2964_/Y _2845_/A _2850_/D _3084_/A _2994_/X vssd1 vssd1 vccd1 vccd1 _2995_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_166_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4734_ _4663_/X _4724_/Y _4733_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5567_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4665_ _4642_/Y _4663_/X _4664_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5551_/D sky130_fd_sc_hd__o211a_1
XFILLER_266_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3616_ _4306_/A vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_134_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4596_ _4593_/Y _4595_/Y _4634_/A vssd1 vssd1 vccd1 vccd1 _4596_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3174__A1 _5601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3174__B2 _5617_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3547_ _5475_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _3549_/A sky130_fd_sc_hd__and2_1
XANTENNA__5482__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3478_ _5419_/Q input55/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2795__A _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5217_ _5755_/Q _3840_/X _5216_/X vssd1 vssd1 vccd1 vccd1 _5217_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5320__C1 _4487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3390__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5148_ _5520_/Q vssd1 vssd1 vccd1 vccd1 _5148_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__3882__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_244_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5079_ _3790_/X _3935_/A _5235_/S vssd1 vssd1 vccd1 vccd1 _5079_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4426__A1 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4977__A2 _4972_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_236 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_233_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4250__A _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3165__A1 _5647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3165__B2 _5567_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A i_req_data[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_279_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5081__A _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4665__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3873__C1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output128_A _5741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4968__A2 _4949_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5090__A1 _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4425__A _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_250_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5020__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5355__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2780_ _5581_/Q _2635_/Y _2657_/X _5661_/Q vssd1 vssd1 vccd1 vccd1 _2780_/X sky130_fd_sc_hd__a22o_1
XFILLER_156_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3475__S _3475_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5256__A _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4450_ _4447_/X _4449_/X _4469_/D vssd1 vssd1 vccd1 vccd1 _4450_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3156__A1 _5629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4353__B1 _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3401_ _2852_/A _5380_/Q _3415_/S vssd1 vssd1 vccd1 vccd1 _3402_/A sky130_fd_sc_hd__mux2_1
X_4381_ _5452_/Q _4103_/A _4379_/X _4380_/X vssd1 vssd1 vccd1 vccd1 _4381_/X sky130_fd_sc_hd__a211o_1
X_3332_ _5349_/Q _3293_/X _3330_/X _5367_/Q vssd1 vssd1 vccd1 vccd1 _5349_/D sky130_fd_sc_hd__a22o_1
X_3263_ _3258_/X _3262_/X _5348_/Q vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__o21ba_1
XFILLER_85_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_285_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4656__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5002_/A vssd1 vssd1 vccd1 vccd1 _5683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_273_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3194_ _5605_/Q _3133_/X _3135_/X _5621_/Q _3193_/X vssd1 vssd1 vccd1 vccd1 _3194_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2765__D _5599_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2781__C _2782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3631__A2 _3596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_i_clk clkbuf_1_1_1_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_i_clk/A
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4187__A3 _4181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5766_ _5766_/A vssd1 vssd1 vccd1 vccd1 _5766_/X sky130_fd_sc_hd__clkbuf_1
X_2978_ _5392_/Q vssd1 vssd1 vccd1 vccd1 _2978_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4592__B1 _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4717_ _4722_/A _4983_/A vssd1 vssd1 vccd1 vccd1 _4717_/Y sky130_fd_sc_hd__nand2_1
X_5697_ _5724_/CLK _5697_/D vssd1 vssd1 vccd1 vccd1 _5697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3385__S _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4648_ _4687_/A vssd1 vssd1 vccd1 vccd1 _4722_/A sky130_fd_sc_hd__buf_2
XFILLER_162_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4344__B1 _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4579_ _4585_/A _4590_/C _4579_/C vssd1 vssd1 vccd1 vccd1 _4579_/X sky130_fd_sc_hd__or3_1
XANTENNA__3698__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2658__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5378__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_232_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3622__A2 _3600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4899__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4583__A0 _5315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3950_ _5516_/Q _3923_/X _3949_/X _3945_/X vssd1 vssd1 vccd1 vccd1 _5516_/D sky130_fd_sc_hd__o211a_1
XFILLER_223_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2901_ _3281_/A _3330_/C _3775_/C _2900_/Y vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__a31o_1
X_3881_ _3956_/A _3908_/B vssd1 vssd1 vccd1 vccd1 _3881_/Y sky130_fd_sc_hd__nand2_1
X_5620_ _5623_/CLK _5620_/D vssd1 vssd1 vccd1 vccd1 _5620_/Q sky130_fd_sc_hd__dfxtp_2
X_2832_ input39/X _5433_/Q _2849_/S vssd1 vssd1 vccd1 vccd1 _2852_/B sky130_fd_sc_hd__mux2_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4574__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5551_ _5747_/CLK _5551_/D vssd1 vssd1 vccd1 vccd1 _5551_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_247_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2763_ _5583_/Q _2635_/Y _2657_/X _5663_/Q vssd1 vssd1 vccd1 vccd1 _2763_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_263 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4502_ _4502_/A _4502_/B vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__xnor2_1
XFILLER_144_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2694_ _2782_/C vssd1 vssd1 vccd1 vccd1 _2771_/B sky130_fd_sc_hd__buf_4
X_5482_ _5722_/CLK _5482_/D vssd1 vssd1 vccd1 vccd1 _5482_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_144_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4433_ _2954_/X _4430_/Y _4432_/X vssd1 vssd1 vccd1 vccd1 _4433_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4364_ _4043_/A _4009_/Y _4041_/X _4363_/Y vssd1 vssd1 vccd1 vccd1 _4364_/X sky130_fd_sc_hd__a31o_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3315_ _5371_/Q _3318_/C _3310_/X _5368_/Q _3293_/A vssd1 vssd1 vccd1 vccd1 _3315_/X
+ sky130_fd_sc_hd__a221o_1
X_4295_ _4090_/A _4090_/B _4066_/Y vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__o21ai_1
XFILLER_258_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3234__A _5300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3246_ _3854_/A _5723_/Q _5722_/Q _3856_/C vssd1 vssd1 vccd1 vccd1 _3843_/B sky130_fd_sc_hd__nor4_4
XFILLER_100_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4049__B _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5520__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3177_ _5553_/Q _3131_/X _3174_/X _3176_/X vssd1 vssd1 vccd1 vccd1 _3177_/X sky130_fd_sc_hd__o22a_2
XFILLER_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5054__A1 _5512_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4262__C1 _5452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3604__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5670__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2812__A0 _5680_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5749_ _5756_/CLK _5749_/D vssd1 vssd1 vccd1 vccd1 _5749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_210_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4317__A0 _4151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_244 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3144__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_72_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output195_A _5478_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3319__A _3319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5237__C _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput109 _5769_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[9] sky130_fd_sc_hd__buf_2
XFILLER_126_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output72_A _5766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5543__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 _3162_/X vssd1 vssd1 vccd1 vccd1 dbg_out[2] sky130_fd_sc_hd__buf_2
XFILLER_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput91 _3187_/X vssd1 vssd1 vccd1 vccd1 dbg_out[7] sky130_fd_sc_hd__buf_2
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3100_ _3100_/A vssd1 vssd1 vccd1 vccd1 _3100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_233_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4080_ _4079_/B _4079_/C _4274_/A vssd1 vssd1 vccd1 vccd1 _4080_/X sky130_fd_sc_hd__o21a_1
XFILLER_163_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3031_ _5393_/Q _3031_/B vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__or2_1
XANTENNA__2893__A _5453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4584__S _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5693__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_263_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3047__B1 _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4982_ _5673_/Q _4972_/B _4981_/Y _4979_/X vssd1 vssd1 vccd1 vccd1 _5673_/D sky130_fd_sc_hd__o211a_1
XFILLER_211_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3933_ _3993_/B vssd1 vssd1 vccd1 vccd1 _3948_/B sky130_fd_sc_hd__buf_2
XANTENNA__2832__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4613__A _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3864_ _4635_/A _4988_/B _3864_/C vssd1 vssd1 vccd1 vccd1 _3905_/S sky130_fd_sc_hd__and3_2
X_5603_ _5653_/CLK _5603_/D vssd1 vssd1 vccd1 vccd1 _5603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2815_ _2815_/A _2815_/B vssd1 vssd1 vccd1 vccd1 _2815_/X sky130_fd_sc_hd__or2_1
X_3795_ _3795_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3795_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5534_ _5685_/CLK _5534_/D vssd1 vssd1 vccd1 vccd1 _5762_/A sky130_fd_sc_hd__dfxtp_2
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2746_ _2747_/D _2733_/A _2747_/B _5585_/Q vssd1 vssd1 vccd1 vccd1 _2746_/X sky130_fd_sc_hd__and4bb_1
XFILLER_127_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5465_ _5743_/CLK _5465_/D vssd1 vssd1 vccd1 vccd1 _5465_/Q sky130_fd_sc_hd__dfxtp_1
X_2677_ _2672_/X _2673_/X _2676_/X _2791_/B _5560_/Q vssd1 vssd1 vccd1 vccd1 _2678_/A
+ sky130_fd_sc_hd__o32a_1
X_4416_ _4050_/A _4415_/Y _4422_/A vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_278_229 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5396_ _5492_/CLK _5396_/D vssd1 vssd1 vccd1 vccd1 _5396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4347_ _4347_/A _4347_/B _4347_/C vssd1 vssd1 vccd1 vccd1 _4347_/X sky130_fd_sc_hd__and3_1
XFILLER_207_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4278_ _4278_/A _4278_/B _4278_/C vssd1 vssd1 vccd1 vccd1 _4279_/B sky130_fd_sc_hd__or3_1
XFILLER_86_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3229_ _5356_/Q _5678_/Q vssd1 vssd1 vccd1 vccd1 _3345_/A sky130_fd_sc_hd__nor2_2
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4235__C1 _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__A1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4523__A _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5416__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3139__A _3139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3210__B1 _3149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5566__CLK _5674_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3573__S _3588_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2697__B _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3513__A1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3602__A _3602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5018__A1 _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output110_A _5548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output208_A _5307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4241__A2 _4326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3748__S _4272_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3201__B1 _3145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3580_ _5476_/Q _3585_/B vssd1 vssd1 vccd1 vccd1 _4027_/A sky130_fd_sc_hd__and2_1
XFILLER_158_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2888__A _3281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2960__C1 _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5250_ _5727_/Q _5081_/A _5253_/S vssd1 vssd1 vccd1 vccd1 _5251_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4201_ _4372_/B vssd1 vssd1 vccd1 vccd1 _4201_/Y sky130_fd_sc_hd__inv_2
X_5181_ _5181_/A vssd1 vssd1 vccd1 vccd1 _5714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_244_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4132_ _4132_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _4373_/B sky130_fd_sc_hd__or2_1
XFILLER_68_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5257__A1 _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2827__S _3000_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4063_ _4063_/A _4030_/A vssd1 vssd1 vccd1 vccd1 _4088_/B sky130_fd_sc_hd__or2b_1
XFILLER_83_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_271_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ _3089_/A vssd1 vssd1 vccd1 vccd1 _3085_/A sky130_fd_sc_hd__buf_2
XFILLER_209_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2773__D _5582_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4480__A2 _4485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5439__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4965_ _5666_/Q _4969_/A vssd1 vssd1 vccd1 vccd1 _4965_/X sky130_fd_sc_hd__or2_1
XFILLER_224_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3916_ _5510_/Q _5067_/B _3918_/B vssd1 vssd1 vccd1 vccd1 _3916_/X sky130_fd_sc_hd__mux2_1
X_4896_ _5636_/Q _4897_/B _4895_/Y _4886_/X vssd1 vssd1 vccd1 vccd1 _5636_/D sky130_fd_sc_hd__o211a_1
XFILLER_149_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3991__A1 _5526_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5589__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3847_ _5263_/A vssd1 vssd1 vccd1 vccd1 _4979_/A sky130_fd_sc_hd__buf_4
XFILLER_164_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3778_ _3778_/A vssd1 vssd1 vccd1 vccd1 _5459_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4535__A3 _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3743__A1 _5575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5517_ _5740_/CLK _5517_/D vssd1 vssd1 vccd1 vccd1 _5517_/Q sky130_fd_sc_hd__dfxtp_2
X_2729_ _5587_/Q _2635_/Y _2686_/X _2727_/X _2728_/X vssd1 vssd1 vccd1 vccd1 _2729_/X
+ sky130_fd_sc_hd__a2111o_1
X_5448_ _5692_/CLK _5448_/D vssd1 vssd1 vccd1 vccd1 _5448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4299__A2 _4148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5379_ _5722_/CLK _5379_/D vssd1 vssd1 vccd1 vccd1 _5379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3259__B1 _5530_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4518__A _4533_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3734__A1 _5670_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4144__D1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3689__D _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4214__A2 _4132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3478__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5731__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _5574_/Q _4747_/B _4749_/Y _4745_/X vssd1 vssd1 vccd1 vccd1 _5574_/D sky130_fd_sc_hd__o211a_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3701_ _5561_/Q _3596_/X _3698_/X _3700_/X vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__o22a_4
XFILLER_174_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4681_ _4642_/Y _4679_/X _4680_/X _4670_/X vssd1 vssd1 vccd1 vccd1 _5554_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3632_ _3673_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _3633_/A sky130_fd_sc_hd__and2_1
XANTENNA__3725__A1 _5557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3563_ _5341_/Q _5343_/Q _5342_/Q vssd1 vssd1 vccd1 vccd1 _3598_/A sky130_fd_sc_hd__and3b_4
XANTENNA__4610__B _5321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5302_ _5325_/B vssd1 vssd1 vccd1 vccd1 _5319_/B sky130_fd_sc_hd__buf_2
XFILLER_154_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3494_ _5427_/Q input32/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3495_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5233_ _5719_/Q _5232_/X _5233_/S vssd1 vssd1 vccd1 vccd1 _5234_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4686__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4150__A1 _4132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5164_ _4590_/B _5193_/B _5163_/Y _5196_/A vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_271_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4115_ _4441_/B _4171_/B _4114_/A vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5095_ _5744_/Q _3840_/A _5051_/B _5531_/Q vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3242__A _5461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_256_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4046_ _4403_/A _4183_/A vssd1 vssd1 vccd1 vccd1 _4046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_392 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4205__A2 _4108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3388__S _3394_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3413__A0 _2835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4948_ _5659_/Q _4935_/B _4947_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5659_/D sky130_fd_sc_hd__o211a_1
XFILLER_212_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3964__A1 _5313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4879_ _5629_/Q _4910_/B vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__or2_1
XFILLER_149_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4801__A _4819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3716__A1 _5562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3192__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3136__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4126__D1 _4128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4141__A1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5604__CLK _5659_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4248__A _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4444__A2 _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_262_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3652__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_346 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4601__C1 _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2758__A2 _2652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3707__A1 _5640_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5018__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3183__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_320 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4380__A1 _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater217 _5762_/A vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__buf_6
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_348 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_241_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4435__A2 _4429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_318 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3997__A _5461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3643__B1 _3607_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_351 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_221_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4802_ _5596_/Q _4834_/B vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__or2_1
XFILLER_61_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2994_ _2965_/Y _2835_/B _2845_/A _2964_/Y _2993_/X vssd1 vssd1 vccd1 vccd1 _2994_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3946__A1 _5515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4733_ _5567_/Q _4759_/B vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__or2_1
XFILLER_159_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4621__A _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4664_ _5551_/Q _4722_/A vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__or2_1
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3615_ _4276_/A _4124_/B _4248_/C vssd1 vssd1 vccd1 vccd1 _3615_/X sky130_fd_sc_hd__and3_2
XFILLER_266_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4595_ _4600_/A _4490_/B _4594_/X vssd1 vssd1 vccd1 vccd1 _4595_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_174_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3237__A _5482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3174__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3546_ _5454_/Q vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__5627__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3477_ _3523_/S vssd1 vssd1 vccd1 vccd1 _3496_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5216_ _5526_/Q _3932_/B _3864_/C _5506_/Q _5053_/X vssd1 vssd1 vccd1 vccd1 _5216_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_215_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_215_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5147_ _5147_/A vssd1 vssd1 vccd1 vccd1 _5711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5078_ _5015_/Y _5156_/B _5077_/X _3790_/X vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__a211o_1
XFILLER_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4029_ _4067_/A _4232_/B vssd1 vssd1 vccd1 vccd1 _4029_/X sky130_fd_sc_hd__or2_1
XANTENNA__3634__A0 _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4831__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3937__A1 _5513_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3147__A _3147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4898__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3165__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5081__B _5125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4665__A2 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input34_A i_req_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2676__A1 _5624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_282_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3625__B1 _3606_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5090__A2 _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4425__B _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4889__C1 _4886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3057__A _5768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4353__A1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3156__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3400_ _3400_/A vssd1 vssd1 vccd1 vccd1 _5379_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4380_ _5450_/Q _4379_/B _4379_/C _4160_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4380_/X
+ sky130_fd_sc_hd__a221o_1
X_3331_ _5348_/Q _3293_/X _3330_/X _5368_/Q vssd1 vssd1 vccd1 vccd1 _5348_/D sky130_fd_sc_hd__a22o_1
XFILLER_258_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3262_ _5351_/Q _3259_/Y _3260_/X _3261_/X _5349_/Q vssd1 vssd1 vccd1 vccd1 _3262_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3313__C1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5001_ _5683_/Q _5337_/Q _5720_/D vssd1 vssd1 vccd1 vccd1 _5002_/A sky130_fd_sc_hd__mux2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3193_ _5669_/Q _3137_/X _3139_/X _5589_/Q vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__a22o_1
XFILLER_273_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4813__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4716__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2781__D _5565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5765_ _5765_/A vssd1 vssd1 vccd1 vccd1 _5765_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_194_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2977_ _5393_/Q vssd1 vssd1 vccd1 vccd1 _2977_/Y sky130_fd_sc_hd__inv_2
X_4716_ input12/X _4689_/X _4690_/X _4715_/Y vssd1 vssd1 vccd1 vccd1 _4983_/A sky130_fd_sc_hd__o2bb2a_4
XANTENNA__4592__A1 _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5696_ _5724_/CLK _5696_/D vssd1 vssd1 vccd1 vccd1 _5696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4647_ _5680_/Q _4950_/B vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__and2_1
XANTENNA__4344__A1 _2936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4344__B2 _2954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4578_ _5539_/Q _4577_/C _5768_/A vssd1 vssd1 vccd1 vccd1 _4579_/C sky130_fd_sc_hd__a21oi_1
X_3529_ _5473_/Q _2768_/Y _3588_/S vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__mux2_8
XFILLER_115_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2658__A1 _5642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2658__B2 _5674_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4583__A1 _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3605__A _3605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4200__S _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2649__A1 _5563_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_267_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2900_ _3281_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _2900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _3880_/A vssd1 vssd1 vccd1 vccd1 _5497_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5472__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2831_ input38/X _5432_/Q _5409_/Q vssd1 vssd1 vccd1 vccd1 _2852_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3486__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4171__A _4171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__A1 _5539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5550_ _5674_/CLK _5550_/D vssd1 vssd1 vccd1 vccd1 _5550_/Q sky130_fd_sc_hd__dfxtp_4
X_2762_ _5631_/Q _2655_/X _2761_/X _5647_/Q vssd1 vssd1 vccd1 vccd1 _2762_/X sky130_fd_sc_hd__a22o_1
XFILLER_191_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4501_ _4501_/A _4501_/B vssd1 vssd1 vccd1 vccd1 _4502_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5481_ _5722_/CLK _5481_/D vssd1 vssd1 vccd1 vccd1 _5481_/Q sky130_fd_sc_hd__dfxtp_4
X_2693_ _2782_/B vssd1 vssd1 vccd1 vccd1 _2727_/C sky130_fd_sc_hd__buf_4
XFILLER_184_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4432_ _2904_/X _4410_/B _4431_/X _4408_/A _4161_/X vssd1 vssd1 vccd1 vccd1 _4432_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_144_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4363_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4363_/Y sky130_fd_sc_hd__nor2_1
XFILLER_263_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3314_ _3601_/B _5486_/D _3313_/X vssd1 vssd1 vccd1 vccd1 _5342_/D sky130_fd_sc_hd__o21a_1
X_4294_ _4294_/A _4294_/B vssd1 vssd1 vccd1 vccd1 _4294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3245_ _3851_/B _3245_/B vssd1 vssd1 vccd1 vccd1 _3245_/Y sky130_fd_sc_hd__nor2_1
XFILLER_273_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3176_ _5633_/Q _3143_/X _3145_/X _3175_/X vssd1 vssd1 vccd1 vccd1 _3176_/X sky130_fd_sc_hd__a211o_1
XFILLER_273_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3250__A _3250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2812__A1 _5681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_167_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4081__A _4083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4565__A1 _4532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5748_ _5756_/CLK _5748_/D vssd1 vssd1 vccd1 vccd1 _5748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5679_ _5721_/CLK _5679_/D vssd1 vssd1 vccd1 vccd1 _5679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3144__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5345__CLK _5738_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3828__A0 _5481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5495__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3056__A1 _2845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4253__B1 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_260_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_198_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3319__B _3791_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output188_A _5471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4308__A1 _4271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5026__S _5030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3335__A _3791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 _5764_/A vssd1 vssd1 vccd1 vccd1 dbg_out[20] sky130_fd_sc_hd__buf_2
Xoutput81 _5774_/A vssd1 vssd1 vccd1 vccd1 dbg_out[30] sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0_i_clk clkbuf_0_i_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_i_clk/A
+ sky130_fd_sc_hd__clkbuf_8
Xoutput92 _3192_/X vssd1 vssd1 vccd1 vccd1 dbg_out[8] sky130_fd_sc_hd__buf_2
XANTENNA_output65_A _5760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_324 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_283_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3030_ _5393_/Q _3031_/B vssd1 vssd1 vccd1 vccd1 _3039_/C sky130_fd_sc_hd__and2_1
XFILLER_95_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_236_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_251_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3047__A1 _2852_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4981_ _4981_/A _4985_/B vssd1 vssd1 vccd1 vccd1 _4981_/Y sky130_fd_sc_hd__nand2_1
X_3932_ _4635_/A _3932_/B vssd1 vssd1 vccd1 vccd1 _3993_/B sky130_fd_sc_hd__nand2_1
XFILLER_251_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3863_ _5082_/B vssd1 vssd1 vccd1 vccd1 _3864_/C sky130_fd_sc_hd__buf_2
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4613__B _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5602_ _5653_/CLK _5602_/D vssd1 vssd1 vccd1 vccd1 _5602_/Q sky130_fd_sc_hd__dfxtp_2
X_2814_ _5684_/Q _5685_/Q _5686_/Q _5687_/Q _3599_/B _3601_/B vssd1 vssd1 vccd1 vccd1
+ _2815_/B sky130_fd_sc_hd__mux4_1
XFILLER_258_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3794_ _3794_/A vssd1 vssd1 vccd1 vccd1 _5465_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4332__C _4332_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5533_ _5685_/CLK _5533_/D vssd1 vssd1 vccd1 vccd1 _5761_/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__3229__B _5678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2745_ _5633_/Q _2655_/X _2657_/X _5665_/Q vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5464_ _5707_/CLK _5464_/D vssd1 vssd1 vccd1 vccd1 _5464_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_172_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2676_ _5624_/Q _2652_/A _2674_/X _2675_/X _2686_/A vssd1 vssd1 vccd1 vccd1 _2676_/X
+ sky130_fd_sc_hd__a2111o_1
X_4415_ _4415_/A _4440_/A vssd1 vssd1 vccd1 vccd1 _4415_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5368__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5395_ _5404_/CLK _5395_/D vssd1 vssd1 vccd1 vccd1 _5395_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3245__A _3851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4346_ _4347_/A _4175_/B _4337_/Y _4345_/Y vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__a211o_4
XANTENNA__2730__B1 _2726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4277_ _4276_/A _4303_/A _4273_/X _4276_/Y _4271_/A vssd1 vssd1 vccd1 vccd1 _4277_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3228_ _3228_/A vssd1 vssd1 vccd1 vccd1 _4987_/B sky130_fd_sc_hd__inv_2
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4076__A _4076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3159_ _5598_/Q _3133_/X _3135_/X _5614_/Q _3158_/X vssd1 vssd1 vccd1 vccd1 _3159_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3038__A1 _4552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4235__B1 _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3589__A2 _4045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4804__A _5597_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4523__B _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4538__A1 _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_335 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_182_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3210__A1 _5656_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3210__B2 _5576_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2697__C _2806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4710__A1 _5560_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_265_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3029__A1 _5081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3201__A1 _5638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_126 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3764__S _4585_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5510__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2888__B _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_114_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _4153_/B _4138_/B _4471_/S vssd1 vssd1 vccd1 vccd1 _4200_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4162__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5180_ _5714_/Q _5179_/X _5233_/S vssd1 vssd1 vccd1 vccd1 _5181_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5660__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4131_ _4373_/A _4177_/B vssd1 vssd1 vccd1 vccd1 _4131_/X sky130_fd_sc_hd__and2_1
XFILLER_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5280__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4062_ _4379_/B _4112_/B _4112_/C vssd1 vssd1 vccd1 vccd1 _4441_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__4465__B1 _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3013_ _2840_/C _3089_/A _3018_/A vssd1 vssd1 vccd1 vccd1 _3013_/X sky130_fd_sc_hd__a21o_1
XFILLER_283_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_202 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_91_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2843__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4964_ _4674_/X _4949_/Y _4963_/X _4957_/X vssd1 vssd1 vccd1 vccd1 _5665_/D sky130_fd_sc_hd__o211a_1
XFILLER_251_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3915_ _5743_/Q _4600_/A _5094_/C _3996_/B vssd1 vssd1 vccd1 vccd1 _3918_/B sky130_fd_sc_hd__and4_1
X_4895_ _4970_/A _4897_/B vssd1 vssd1 vccd1 vccd1 _4895_/Y sky130_fd_sc_hd__nand2_1
X_3846_ _5229_/S _4523_/B _5294_/B vssd1 vssd1 vccd1 vccd1 _3846_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_164_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3777_ _5294_/A _3775_/X _3813_/S vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__mux2_1
XFILLER_285_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3743__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2728_ _2727_/C _2775_/B _5651_/Q _2775_/D vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__and4b_1
X_5516_ _5741_/CLK _5516_/D vssd1 vssd1 vccd1 vccd1 _5516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_285_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2798__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5447_ _5692_/CLK _5447_/D vssd1 vssd1 vccd1 vccd1 _5447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2659_ _2747_/D _2682_/A _2761_/B _5610_/Q vssd1 vssd1 vccd1 vccd1 _2659_/X sky130_fd_sc_hd__and4b_1
XFILLER_218_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4299__A3 _4149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5378_ _5441_/CLK _5378_/D vssd1 vssd1 vccd1 vccd1 _5378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4329_ _5450_/Q _4033_/A _4071_/B _5446_/Q _4160_/A vssd1 vssd1 vccd1 vccd1 _4329_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3259__A1 _5528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4518__B _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_215_311 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3195__B1 _3149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3734__A2 _3600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5683__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_92_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _5641_/Q _3605_/X _3606_/X _3699_/X vssd1 vssd1 vccd1 vccd1 _3700_/X sky130_fd_sc_hd__a211o_1
XFILLER_186_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680_ _5554_/Q _4687_/A vssd1 vssd1 vccd1 vccd1 _4680_/X sky130_fd_sc_hd__or2_1
XFILLER_169_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3631_ _5552_/Q _3596_/A _3628_/X _3630_/X vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__o22a_4
XFILLER_186_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5175__B2 _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3494__S _3496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3186__B1 _3145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4383__C1 _4382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3725__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3562_ _5342_/Q _3599_/B _3601_/C vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__and3b_4
XANTENNA__4922__A1 _4663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5301_ _5301_/A vssd1 vssd1 vccd1 vccd1 _5743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3493_ _3493_/A vssd1 vssd1 vccd1 vccd1 _5426_/D sky130_fd_sc_hd__clkbuf_1
X_5232_ _5231_/X _2650_/Y _5464_/Q vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4150__A2 _4024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2838__S _5409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5163_ _5750_/Q _3840_/X _5162_/X vssd1 vssd1 vccd1 vccd1 _5163_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4114_ _4114_/A _4441_/B _4171_/B vssd1 vssd1 vccd1 vccd1 _4114_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__5406__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5094_ _5515_/Q _5094_/B _5094_/C vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__and3_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4045_ _4045_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__nor2_1
XFILLER_204_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_271_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5556__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4947_ _4985_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4947_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4878_ _4646_/X _4874_/Y _4877_/X _4862_/X vssd1 vssd1 vccd1 vccd1 _5628_/D sky130_fd_sc_hd__o211a_1
X_3829_ _3829_/A vssd1 vssd1 vccd1 vccd1 _5481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_229_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3716__A2 _3596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4126__C1 _4128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3136__C input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4677__A0 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4141__A2 _4363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4529__A _4529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4248__B _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3652__A1 _5614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3652__B2 _5598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2860__C1 _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_i_clk clkbuf_2_1_0_i_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_i_clk/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_130_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_358 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5157__A1 _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3608__A _3608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3168__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__A1 _5640_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3707__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output170_A _3091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4380__A2 _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5429__CLK _5441_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater216_A _5764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3343__A _5331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_238_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5579__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3997__B _5051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3643__A1 _5634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3643__B2 _5570_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_363 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_261_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4801_ _4819_/A vssd1 vssd1 vccd1 vccd1 _4834_/B sky130_fd_sc_hd__buf_6
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2993_ _2965_/Y _2835_/B _2992_/X vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__o21a_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4732_ _4658_/X _4724_/Y _4731_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5566_/D sky130_fd_sc_hd__o211a_1
XFILLER_119_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4663_ _4663_/A vssd1 vssd1 vccd1 vccd1 _4663_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2752__A_N _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3159__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3614_ _4132_/A _3572_/X _4469_/B _4469_/C _3613_/X vssd1 vssd1 vccd1 vccd1 _4248_/C
+ sky130_fd_sc_hd__o2111a_1
X_4594_ _4626_/S _5317_/A _5229_/S vssd1 vssd1 vccd1 vccd1 _4594_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3237__B _5485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3545_ _5455_/Q vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__inv_2
XFILLER_127_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3952__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3476_ _3476_/A vssd1 vssd1 vccd1 vccd1 _5418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_282_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5215_ _5526_/Q vssd1 vssd1 vccd1 vccd1 _5215_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_282_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3253__A _5291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5146_ _5711_/Q _5145_/Y _5233_/S vssd1 vssd1 vccd1 vccd1 _5147_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_350 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5077_ _5060_/B _5060_/Y _5077_/S vssd1 vssd1 vccd1 vccd1 _5077_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4028_ _4033_/A _4071_/B vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__or2_1
XFILLER_244_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3634__A1 _4063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3399__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4812__A _5601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5139__A1 _5539_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4259__A _5453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5721__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_208 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2676__A2 _2652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input27_A i_req_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3625__A1 _5633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4425__C _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2775__A_N _2727_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3057__B _3063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4353__A2 _4121_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3561__B1 _3608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _5242_/S _3775_/B _3330_/C _3775_/C vssd1 vssd1 vccd1 vccd1 _3330_/X sky130_fd_sc_hd__and4_1
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3261_ _5528_/Q _3265_/A _5351_/Q vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__a21bo_1
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3313__B1 _3310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5000_ _5000_/A vssd1 vssd1 vccd1 vccd1 _5682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3192_ _5556_/Q _3131_/X _3189_/X _3191_/X vssd1 vssd1 vccd1 vccd1 _3192_/X sky130_fd_sc_hd__o22a_1
XFILLER_285_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_81_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_179 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3077__C1 _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3947__S _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5764_ _5764_/A vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__clkbuf_1
X_2976_ _5394_/Q vssd1 vssd1 vccd1 vccd1 _2976_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4715_ _5718_/Q vssd1 vssd1 vccd1 vccd1 _4715_/Y sky130_fd_sc_hd__inv_2
X_5695_ _5724_/CLK _5695_/D vssd1 vssd1 vccd1 vccd1 _5695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3248__A _5508_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4646_ _4646_/A vssd1 vssd1 vccd1 vccd1 _4646_/X sky130_fd_sc_hd__buf_4
XFILLER_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4577_ _5768_/A _5767_/A _4577_/C vssd1 vssd1 vccd1 vccd1 _4590_/C sky130_fd_sc_hd__and3_1
XANTENNA__5744__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3528_ _3528_/A vssd1 vssd1 vccd1 vccd1 _3588_/S sky130_fd_sc_hd__buf_6
XFILLER_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4079__A _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3459_ _5410_/Q input24/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3460_/A sky130_fd_sc_hd__mux2_1
XFILLER_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2658__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_257_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129_ _4599_/B _5128_/X _4561_/Y vssd1 vssd1 vccd1 vccd1 _5131_/C sky130_fd_sc_hd__o21a_1
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3068__C1 _3016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4542__A _5516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_200_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_267_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4740__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_267_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3846__A1 _5229_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2649__A2 _2791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2830_ _2830_/A _3003_/C vssd1 vssd1 vccd1 vccd1 _2830_/Y sky130_fd_sc_hd__nor2_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4574__A2 _4511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2761_ _2682_/A _2761_/B _5344_/Q vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__and3b_1
XFILLER_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4500_ _4500_/A _5015_/A vssd1 vssd1 vccd1 vccd1 _4501_/B sky130_fd_sc_hd__xor2_2
XFILLER_191_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5480_ _5722_/CLK _5480_/D vssd1 vssd1 vccd1 vccd1 _5480_/Q sky130_fd_sc_hd__dfxtp_4
X_2692_ _2757_/D vssd1 vssd1 vccd1 vccd1 _2806_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_129_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4431_ _5445_/Q _4484_/A _2919_/X vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5283__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4362_ _4362_/A _5156_/A _4362_/C _4362_/D vssd1 vssd1 vccd1 vccd1 _4401_/B sky130_fd_sc_hd__or4_1
X_3313_ _5372_/Q _3318_/C _3310_/X _5369_/Q _3293_/A vssd1 vssd1 vccd1 vccd1 _3313_/X
+ sky130_fd_sc_hd__a221o_1
X_4293_ _4071_/C _4033_/X _4322_/B _4350_/A vssd1 vssd1 vccd1 vccd1 _4294_/B sky130_fd_sc_hd__o31a_1
XFILLER_258_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3244_ _5347_/Q _4619_/B _3989_/S _5291_/S vssd1 vssd1 vccd1 vccd1 _3245_/B sky130_fd_sc_hd__o31a_1
XFILLER_273_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2846__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3175_ _5649_/Q _3147_/X _3149_/X _5569_/Q vssd1 vssd1 vccd1 vccd1 _3175_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3531__A _5468_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4798__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4262__A1 _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4262__B2 _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4362__A _4362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4014__A1 _4278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5177__B _5177_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4081__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5747_ _5747_/CLK _5747_/D vssd1 vssd1 vccd1 vccd1 _5747_/Q sky130_fd_sc_hd__dfxtp_1
X_2959_ _2959_/A vssd1 vssd1 vccd1 vccd1 _5446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3773__B1 _3775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5678_ _5743_/CLK _5678_/D vssd1 vssd1 vccd1 vccd1 _5678_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4629_ _4629_/A _4629_/B vssd1 vssd1 vccd1 vccd1 _4633_/B sky130_fd_sc_hd__nor2_1
XFILLER_237_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5193__A _5772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4301__S _4301_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3144__C input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4537__A _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_272_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4789__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4253__A1 _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3764__A0 _4527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4700__A2_N _4689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3616__A _4306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4211__S _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput60 _3207_/X vssd1 vssd1 vccd1 vccd1 dbg_out[11] sky130_fd_sc_hd__buf_2
Xoutput71 _5765_/A vssd1 vssd1 vccd1 vccd1 dbg_out[21] sky130_fd_sc_hd__buf_2
Xoutput82 _5775_/A vssd1 vssd1 vccd1 vccd1 dbg_out[31] sky130_fd_sc_hd__buf_2
Xoutput93 _3197_/X vssd1 vssd1 vccd1 vccd1 dbg_out[9] sky130_fd_sc_hd__buf_2
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output58_A _3152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5042__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_323 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4244__A1 _4171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4980_ _5672_/Q _4972_/B _4978_/Y _4979_/X vssd1 vssd1 vccd1 vccd1 _5672_/D sky130_fd_sc_hd__o211a_1
XFILLER_63_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3931_ _3931_/A vssd1 vssd1 vccd1 vccd1 _3932_/B sky130_fd_sc_hd__buf_2
XANTENNA__4182__A _4454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3862_ _3862_/A vssd1 vssd1 vccd1 vccd1 _5082_/B sky130_fd_sc_hd__clkbuf_2
X_5601_ _5680_/CLK _5601_/D vssd1 vssd1 vccd1 vccd1 _5601_/Q sky130_fd_sc_hd__dfxtp_2
X_2813_ _3601_/C vssd1 vssd1 vccd1 vccd1 _2815_/A sky130_fd_sc_hd__clkinv_2
X_3793_ _5465_/Q _5456_/Q _3813_/S vssd1 vssd1 vccd1 vccd1 _3794_/A sky130_fd_sc_hd__mux2_1
X_5532_ _5707_/CLK _5532_/D vssd1 vssd1 vccd1 vccd1 _5532_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4910__A _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2744_ _5569_/Q _2644_/X _2664_/X _5601_/Q vssd1 vssd1 vccd1 vccd1 _2744_/X sky130_fd_sc_hd__a22o_1
XFILLER_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5463_ _5757_/CLK _5463_/D vssd1 vssd1 vccd1 vccd1 _5463_/Q sky130_fd_sc_hd__dfxtp_1
X_2675_ _2733_/A _2761_/B _5656_/Q _2681_/A vssd1 vssd1 vccd1 vccd1 _2675_/X sky130_fd_sc_hd__and4b_1
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4414_ _4050_/A _3703_/C _4440_/A vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__a21boi_2
XFILLER_132_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5394_ _5404_/CLK _5394_/D vssd1 vssd1 vccd1 vccd1 _5394_/Q sky130_fd_sc_hd__dfxtp_1
X_4345_ _4171_/A _4339_/X _4340_/X _4341_/X _4344_/Y vssd1 vssd1 vccd1 vccd1 _4345_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_98_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3960__S _3984_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2730__A1 _5555_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4276_ _4276_/A _4276_/B vssd1 vssd1 vccd1 vccd1 _4276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3227_ _5563_/Q _3131_/A _3224_/X _3226_/X vssd1 vssd1 vccd1 vccd1 _3227_/X sky130_fd_sc_hd__o22a_2
XFILLER_223_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_252 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3158_ _5662_/Q _3137_/X _3139_/X _5582_/Q vssd1 vssd1 vccd1 vccd1 _3158_/X sky130_fd_sc_hd__a22o_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4235__A1 _4454_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3089_ _3089_/A _3089_/B vssd1 vssd1 vccd1 vccd1 _3089_/Y sky130_fd_sc_hd__nor2_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4804__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4092__A _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4538__A2 _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_347 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4820__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3210__A2 _3147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2697__D _5638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5462__CLK _5692_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3737__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4934__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3201__A2 _3143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5037__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__A _4987_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2960__B2 _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_385 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4162__B1 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4130_ _5454_/Q _4130_/B vssd1 vssd1 vccd1 vccd1 _4177_/B sky130_fd_sc_hd__or2_1
XFILLER_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2709__A_N _2775_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_283_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4061_ _4403_/A _4183_/A vssd1 vssd1 vccd1 vccd1 _4112_/C sky130_fd_sc_hd__or2_1
XANTENNA__4177__A _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3012_ _5355_/Q _5678_/Q vssd1 vssd1 vccd1 vccd1 _3018_/A sky130_fd_sc_hd__or2_2
XFILLER_260_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_76_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4905__A _4981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4217__A1 _4483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ _5665_/Q _4969_/A vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__or2_1
XFILLER_269_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2779__A1 _5629_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2779__B2 _5645_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3914_ _3914_/A vssd1 vssd1 vccd1 vccd1 _5509_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3020__S _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4894_ _4894_/A vssd1 vssd1 vccd1 vccd1 _4897_/B sky130_fd_sc_hd__buf_4
XFILLER_149_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5335__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3845_ _5219_/S vssd1 vssd1 vccd1 vccd1 _5229_/S sky130_fd_sc_hd__buf_4
XANTENNA__3955__S _5329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_192_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3728__B1 _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3776_ _5242_/S vssd1 vssd1 vccd1 vccd1 _3813_/S sky130_fd_sc_hd__buf_4
XFILLER_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5515_ _5741_/CLK _5515_/D vssd1 vssd1 vccd1 vccd1 _5515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2727_ _5667_/Q _2775_/D _2727_/C _2775_/B vssd1 vssd1 vccd1 vccd1 _2727_/X sky130_fd_sc_hd__and4_1
XANTENNA__4940__A2 _4935_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3256__A _5529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5446_ _5692_/CLK _5446_/D vssd1 vssd1 vccd1 vccd1 _5446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5485__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2658_ _5642_/Q _2655_/X _2657_/X _5674_/Q vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__a22o_1
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5377_ _5441_/CLK _5377_/D vssd1 vssd1 vccd1 vccd1 _5377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2703__A1 _5558_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2703__B2 _2702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4328_ _3555_/C _4265_/X _4327_/X _4116_/A vssd1 vssd1 vccd1 vccd1 _4332_/C sky130_fd_sc_hd__a211o_1
XFILLER_259_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input1_A dbg_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4087__A _4087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4259_ _5453_/Q _4259_/B vssd1 vssd1 vccd1 vccd1 _4259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_234_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4456__A1 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4815__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3967__A0 _4590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3719__A0 _3717_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4916__C1 _4908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4392__B1 _2904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3195__B2 _5573_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_341 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4144__B1 _4469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input57_A i_rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4709__B _4978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__A1 _4140_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output213_A _3250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4725__A _5681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3670__A2 _3935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5358__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ _5632_/Q _3605_/X _3606_/A _3629_/X vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__a211o_1
XFILLER_186_296 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3186__A1 _5635_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3561_ _5612_/Q _3597_/A _3608_/A _5580_/Q vssd1 vssd1 vccd1 vccd1 _3561_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4922__A2 _4912_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3076__A _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5300_ _5300_/A _5300_/B vssd1 vssd1 vccd1 vccd1 _5301_/A sky130_fd_sc_hd__or2_1
X_3492_ _5426_/Q input31/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3493_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5231_ _4482_/B _5230_/Y _5231_/S vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4686__A1 _4642_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5162_ _5521_/Q _3932_/B _3864_/C _5501_/Q vssd1 vssd1 vccd1 vccd1 _5162_/X sky130_fd_sc_hd__a22o_1
XFILLER_271_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4619__B _4619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4113_ _4110_/X _4111_/Y _4441_/B _4112_/X vssd1 vssd1 vccd1 vccd1 _4171_/B sky130_fd_sc_hd__a211oi_4
XFILLER_256_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_271_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5093_ _5763_/A _5125_/A vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__and2_1
XFILLER_271_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _4009_/Y _4041_/X _4108_/C vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__a21oi_2
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2854__S _3768_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4635__A _4635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _5658_/Q _4935_/B _4945_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5658_/D sky130_fd_sc_hd__o211a_1
XFILLER_220_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _5628_/Q _4910_/B vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__or2_1
XFILLER_165_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3828_ _5481_/Q _5385_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3829_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4374__A0 _4140_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3177__A1 _5553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3759_ _5512_/Q _3844_/A vssd1 vssd1 vccd1 vccd1 _3759_/X sky130_fd_sc_hd__or2_1
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3582__D1 _4027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4126__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5429_ _5441_/CLK _5429_/D vssd1 vssd1 vccd1 vccd1 _5429_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4677__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5500__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3652__A2 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4601__A1 _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3168__A1 _5664_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4365__B1 _4322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3168__B2 _5584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4904__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4117__B1 _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5314__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2679__B1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3343__B _3343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_238_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3643__A2 _3605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _5683_/Q _4950_/B vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__and2_4
XFILLER_206_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_375 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2992_ _2968_/X _2969_/X _2972_/X _2991_/X vssd1 vssd1 vccd1 vccd1 _2992_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4731_ _5566_/Q _4759_/B vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__or2_1
XFILLER_221_189 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5286__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4662_ _5707_/Q _4661_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3159__A1 _5598_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3613_ _4128_/C vssd1 vssd1 vccd1 vccd1 _3613_/X sky130_fd_sc_hd__buf_2
XANTENNA__4356__B1 _4232_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3159__B2 _5614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4593_ _5522_/Q _4599_/B vssd1 vssd1 vccd1 vccd1 _4593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3237__C _5484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3544_ _4326_/A _4122_/B vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__2849__S _2849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3475_ _5418_/Q input54/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3476_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4203__S0 _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _5225_/B _5214_/B vssd1 vssd1 vccd1 vccd1 _5220_/A sky130_fd_sc_hd__and2b_1
XFILLER_276_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5145_ _5179_/S _5143_/X _5144_/Y vssd1 vssd1 vccd1 vccd1 _5145_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__5523__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_229_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5076_ _5219_/S _5071_/X _5075_/X _4514_/X vssd1 vssd1 vccd1 vccd1 _5077_/S sky130_fd_sc_hd__a31o_2
XANTENNA__5084__A1 _5514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4027_ _4027_/A _4027_/B vssd1 vssd1 vccd1 vccd1 _4033_/A sky130_fd_sc_hd__or2_2
XFILLER_37_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4831__A1 _5609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5673__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _5651_/Q _4931_/A vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__or2_1
XANTENNA__4812__B _4819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5196__A _5196_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3709__A _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4304__S _4304_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5346__D _5346_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4898__A1 _5637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5135__S _5135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5075__A1 _5742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3086__B1 _3018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3625__A2 _3605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4722__B _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4889__A1 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3561__A1 _5612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output88_A _3172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3561__B2 _5580_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5546__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_325 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3260_ _5530_/Q _5350_/Q _5528_/Q vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4510__B1 _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3191_ _5636_/Q _3143_/X _3145_/X _3190_/X vssd1 vssd1 vccd1 vccd1 _3191_/X sky130_fd_sc_hd__a211o_1
XFILLER_285_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5696__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_294 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_226_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_361 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4813__A1 _4674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4913__A _5686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5763_ _5763_/A vssd1 vssd1 vccd1 vccd1 _5763_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_277_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ _5395_/Q vssd1 vssd1 vccd1 vccd1 _2975_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_380 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4714_ _5561_/Q _4697_/A _4713_/Y _4670_/X vssd1 vssd1 vccd1 vccd1 _5561_/D sky130_fd_sc_hd__o211a_1
X_5694_ _5724_/CLK _5694_/D vssd1 vssd1 vccd1 vccd1 _5694_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4329__B1 _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4645_ _5704_/Q _4643_/X _4690_/A vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3963__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4576_ _5520_/Q _4575_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _4576_/X sky130_fd_sc_hd__mux2_1
X_3527_ _5468_/Q vssd1 vssd1 vccd1 vccd1 _3528_/A sky130_fd_sc_hd__clkinv_4
XFILLER_115_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4079__B _4079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_170_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3458_ _5678_/Q _4987_/A _3458_/C _3458_/D vssd1 vssd1 vccd1 vccd1 _5409_/D sky130_fd_sc_hd__nor4_1
XFILLER_226_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3389_ _3389_/A vssd1 vssd1 vccd1 vccd1 _5374_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5128_ _5766_/A _5193_/B _5127_/Y _5460_/Q vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_217_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5059_ _5050_/X _5058_/X _5460_/Q _3759_/X vssd1 vssd1 vccd1 vccd1 _5060_/B sky130_fd_sc_hd__o211a_2
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5419__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5569__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_193_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5296__A1 _5742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3846__A2 _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4717__B _4983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_263_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output126_A _5742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3113__S _3113_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2952__S _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4733__A _5567_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3349__A _3419_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_129_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2760_ _3948_/A vssd1 vssd1 vccd1 vccd1 _2760_/Y sky130_fd_sc_hd__inv_2
X_2691_ _2791_/B vssd1 vssd1 vccd1 vccd1 _2720_/B sky130_fd_sc_hd__buf_6
XFILLER_247_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4430_ _4483_/B vssd1 vssd1 vccd1 vccd1 _4430_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3534__A1 _3532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4361_ _4361_/A _5132_/A _4543_/B _4499_/B vssd1 vssd1 vccd1 vccd1 _4362_/D sky130_fd_sc_hd__or4_1
XFILLER_6_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_152_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3312_ _3601_/C _5486_/D _3311_/X vssd1 vssd1 vccd1 vccd1 _5341_/D sky130_fd_sc_hd__o21a_1
XFILLER_112_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4292_ _4033_/X _4322_/B _4071_/C vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__o21ai_1
XFILLER_193_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3243_ _4988_/B vssd1 vssd1 vccd1 vccd1 _5291_/S sky130_fd_sc_hd__buf_6
XANTENNA__3298__B1 _3795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4908__A _4979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3174_ _5601_/Q _3133_/X _3135_/X _5617_/Q _3173_/X vssd1 vssd1 vccd1 vccd1 _3174_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_273_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_395 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_275 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4262__A2 _3617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2812__A3 _5683_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4362__B _5156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4014__A2 _4278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5211__A1 _5323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5711__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_194_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5746_ _5747_/CLK _5746_/D vssd1 vssd1 vccd1 vccd1 _5746_/Q sky130_fd_sc_hd__dfxtp_1
X_2958_ _5446_/Q _3283_/C _3337_/B vssd1 vssd1 vccd1 vccd1 _2959_/A sky130_fd_sc_hd__mux2_1
XFILLER_194_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3773__A1 _5458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5677_ _5716_/CLK _5677_/D vssd1 vssd1 vccd1 vccd1 _5677_/Q sky130_fd_sc_hd__dfxtp_1
X_2889_ _2922_/A _2889_/B vssd1 vssd1 vccd1 vccd1 _3799_/B sky130_fd_sc_hd__or2_4
XFILLER_135_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4628_ _5774_/A vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__inv_2
X_4559_ _4577_/C vssd1 vssd1 vccd1 vccd1 _4559_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_312 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_150_228 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_249_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4537__B _4537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_301 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3134__C_N input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5202__A1 _5321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5391__CLK _5404_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3213__B1 _3139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3284__C_N _3775_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_214 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_147_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_353 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_126_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3335__C _3335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput61 _3212_/X vssd1 vssd1 vccd1 vccd1 dbg_out[12] sky130_fd_sc_hd__buf_2
Xoutput72 _5766_/A vssd1 vssd1 vccd1 vccd1 dbg_out[22] sky130_fd_sc_hd__buf_2
Xoutput83 _4987_/B vssd1 vssd1 vccd1 vccd1 dbg_out[32] sky130_fd_sc_hd__buf_2
Xoutput94 _5760_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[0] sky130_fd_sc_hd__buf_2
XANTENNA__4477__C1 _3986_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_255_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_245 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_251_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5734__CLK _5740_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _5094_/B _5094_/C vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__and2_2
XFILLER_251_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3861_ _5471_/Q _3996_/B _5055_/C vssd1 vssd1 vccd1 vccd1 _3862_/A sky130_fd_sc_hd__and3_1
X_5600_ _5680_/CLK _5600_/D vssd1 vssd1 vccd1 vccd1 _5600_/Q sky130_fd_sc_hd__dfxtp_1
X_2812_ _5680_/Q _5681_/Q _5682_/Q _5683_/Q _3599_/B _3601_/B vssd1 vssd1 vccd1 vccd1
+ _2812_/X sky130_fd_sc_hd__mux4_1
XFILLER_258_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3204__B1 _3135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5185__A1_N _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3792_ _3790_/X _3780_/A _3791_/X vssd1 vssd1 vccd1 vccd1 _5464_/D sky130_fd_sc_hd__o21a_1
X_5531_ _5707_/CLK _5531_/D vssd1 vssd1 vccd1 vccd1 _5531_/Q sky130_fd_sc_hd__dfxtp_2
X_2743_ _3956_/A vssd1 vssd1 vccd1 vccd1 _2743_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4910__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5294__A _5294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5462_ _5692_/CLK _5462_/D vssd1 vssd1 vccd1 vccd1 _5462_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_172_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2674_ _2681_/A _2682_/A _2761_/B _5592_/Q vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__and4bb_1
XFILLER_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4704__B1 _4690_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4413_ _4413_/A _4413_/B vssd1 vssd1 vccd1 vccd1 _4484_/B sky130_fd_sc_hd__nor2_2
XANTENNA__2788__A_N _2774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_274_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5393_ _5404_/CLK _5393_/D vssd1 vssd1 vccd1 vccd1 _5393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4344_ _2936_/X _4348_/B _4087_/A _2954_/X _4343_/X vssd1 vssd1 vccd1 vccd1 _4344_/Y
+ sky130_fd_sc_hd__a221oi_1
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2730__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4275_ _4304_/S _4229_/B _4234_/B _4274_/Y vssd1 vssd1 vccd1 vccd1 _4276_/B sky130_fd_sc_hd__o22a_1
XANTENNA__3542__A _4276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3226_ _5643_/Q _3143_/A _3145_/A _3225_/X vssd1 vssd1 vccd1 vccd1 _3226_/X sky130_fd_sc_hd__a211o_1
XFILLER_39_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3157_ _5549_/Q _3131_/X _3154_/X _3156_/X vssd1 vssd1 vccd1 vccd1 _3157_/X sky130_fd_sc_hd__o22a_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3088_ _5405_/Q _3088_/B vssd1 vssd1 vccd1 vccd1 _3089_/B sky130_fd_sc_hd__xnor2_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4373__A _4373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4092__B _4092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5729_ _5740_/CLK _5729_/D vssd1 vssd1 vccd1 vccd1 _5729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4820__B _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_117_86 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5143__S _5200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5120__B1 _5156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5757__CLK _5757_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_370 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_280_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_133_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_195 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4631__C1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3737__A1 _5638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output193_A _5476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4222__S _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3346__B _3346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4698__C1 _4670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4162__A1 _2919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4162__B2 _4333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output70_A _5764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4458__A _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4060_ _4441_/A _4060_/B vssd1 vssd1 vccd1 vccd1 _4114_/A sky130_fd_sc_hd__and2b_1
XFILLER_209_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3011_ _3011_/A vssd1 vssd1 vccd1 vccd1 _3089_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_283_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_190_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_223 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4905__B _4910_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4217__A2 _4213_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5289__A _5292_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_224_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4962_ _4668_/X _4949_/Y _4961_/X _4957_/X vssd1 vssd1 vccd1 vccd1 _5664_/D sky130_fd_sc_hd__o211a_1
XFILLER_196_209 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2779__A2 _2655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3913_ _5261_/A _3913_/B vssd1 vssd1 vccd1 vccd1 _3914_/A sky130_fd_sc_hd__and2_1
XANTENNA__3976__A1 _5319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4893_ _4684_/X _4874_/Y _4892_/X _4886_/X vssd1 vssd1 vccd1 vccd1 _5635_/D sky130_fd_sc_hd__o211a_1
XFILLER_269_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5178__A0 _4490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4921__A _5647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3844_ _3844_/A vssd1 vssd1 vccd1 vccd1 _5219_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_149_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3728__A1 _5572_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3728__B2 _5604_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3775_ _3775_/A _3775_/B _3775_/C vssd1 vssd1 vccd1 vccd1 _3775_/X sky130_fd_sc_hd__and3_1
XFILLER_164_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_157_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5514_ _5741_/CLK _5514_/D vssd1 vssd1 vccd1 vccd1 _5514_/Q sky130_fd_sc_hd__dfxtp_2
X_2726_ _5619_/Q _2652_/X _2723_/X _2724_/X _2725_/X vssd1 vssd1 vccd1 vccd1 _2726_/X
+ sky130_fd_sc_hd__a2111o_4
X_5445_ _5528_/CLK _5445_/D vssd1 vssd1 vccd1 vccd1 _5445_/Q sky130_fd_sc_hd__dfxtp_4
X_2657_ _2657_/A vssd1 vssd1 vccd1 vccd1 _2657_/X sky130_fd_sc_hd__buf_4
XANTENNA__3971__S _3988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5376_ _5743_/CLK _5376_/D vssd1 vssd1 vccd1 vccd1 _5376_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2703__A2 _2720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4327_ _3617_/A _4454_/B _4454_/C _4306_/X _4326_/X vssd1 vssd1 vccd1 vccd1 _4327_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_247_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_259_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5102__B1 _5235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4258_ _5449_/Q _4257_/X vssd1 vssd1 vccd1 vccd1 _4258_/X sky130_fd_sc_hd__or2b_1
X_3209_ _5608_/Q _3133_/A _3135_/A _5624_/Q _3208_/X vssd1 vssd1 vccd1 vccd1 _3209_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4189_ _4617_/A _4617_/B _5200_/A vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__nand3_1
XFILLER_227_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3719__A1 _4307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4392__A1 _5449_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3195__A2 _3147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_128_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4144__A1 _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_151_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4278__A _4278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_307 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4725__B _4949_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_93 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3407__A0 _2850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output206_A _2768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3121__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A1 _5518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__B1 _4274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4741__A _5571_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3186__A2 _3143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4383__A1 _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ _3601_/C _3599_/B _5342_/Q vssd1 vssd1 vccd1 vccd1 _3608_/A sky130_fd_sc_hd__nor3b_4
X_3491_ _3491_/A vssd1 vssd1 vccd1 vccd1 _5425_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5230_ _5230_/A _5230_/B vssd1 vssd1 vccd1 vccd1 _5230_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4686__A2 _4684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5161_ _5521_/Q vssd1 vssd1 vccd1 vccd1 _5161_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4112_ _4379_/B _4112_/B _4112_/C vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__and3_1
X_5092_ _5090_/Y _5091_/X _5706_/Q _5235_/S vssd1 vssd1 vccd1 vccd1 _5706_/D sky130_fd_sc_hd__a2bb2o_1
XFILLER_256_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4043_ _4043_/A _4043_/B vssd1 vssd1 vccd1 vccd1 _4108_/C sky130_fd_sc_hd__nand2_2
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3646__A0 _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4843__C1 _4840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_209_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4635__B _4635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_271_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_212_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4945_ _4983_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4876_ _4894_/A vssd1 vssd1 vccd1 vccd1 _4910_/B sky130_fd_sc_hd__buf_4
XANTENNA__5452__CLK _5528_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3827_ _3827_/A vssd1 vssd1 vccd1 vccd1 _5480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_220_382 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4374__A1 _4141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3177__A2 _3131_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3758_ _5459_/Q vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__inv_2
XFILLER_229_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2709_ _2775_/D _2727_/C _2775_/B _5589_/Q vssd1 vssd1 vccd1 vccd1 _2709_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__3601__A_N _3599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3689_ _5452_/Q _5451_/Q _5448_/Q _5450_/Q vssd1 vssd1 vccd1 vccd1 _3690_/D sky130_fd_sc_hd__or4_1
XFILLER_133_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4126__A1 _5454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5428_ _5441_/CLK _5428_/D vssd1 vssd1 vccd1 vccd1 _5428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5359_ _5724_/CLK _5359_/D vssd1 vssd1 vccd1 vccd1 _5359_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_245_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4429__A2 _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5087__C1 _5060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4826__A _4976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3637__B1 _3598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2860__A1 _5357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4561__A _5518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_156_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3168__A2 _3137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2915__A2 _5486_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3325__C1 _3293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2679__A1 _5575_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2679__B2 _5607_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3343__C _3343_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3628__B1 _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_340 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4455__B _4455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_249 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5475__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2991_ _2987_/X _2989_/X _2990_/X vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _4653_/X _4724_/Y _4729_/X _4718_/X vssd1 vssd1 vccd1 vccd1 _5565_/D sky130_fd_sc_hd__o211a_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4661_ input9/X input16/X _4682_/S vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2717__B_N _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3612_ _4124_/A _4484_/A vssd1 vssd1 vccd1 vccd1 _4128_/C sky130_fd_sc_hd__or2_1
XANTENNA__4356__A1 _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3159__A2 _3133_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4592_ _4590_/B _4590_/C _5770_/A vssd1 vssd1 vccd1 vccd1 _4592_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3543_ _4132_/A _4307_/B vssd1 vssd1 vccd1 vccd1 _4122_/B sky130_fd_sc_hd__nand2_4
XFILLER_115_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3815__A _5242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3474_ _3474_/A vssd1 vssd1 vccd1 vccd1 _5417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5213_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5717_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4203__S1 _4231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_360 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3331__A2 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5144_ _5179_/S _5311_/A vssd1 vssd1 vccd1 vccd1 _5144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_215_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_96_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5075_ _5742_/Q _3840_/A _5072_/X _5073_/X _5074_/X vssd1 vssd1 vccd1 vccd1 _5075_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4816__C1 _4815_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4026_ _4034_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__or2_1
XFILLER_37_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4831__A2 _4822_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4595__A1 _4600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _4679_/X _4912_/Y _4927_/X _4908_/X vssd1 vssd1 vccd1 vccd1 _5650_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4972_/A _4859_/B vssd1 vssd1 vccd1 vccd1 _4859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4898__A2 _4897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_180_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5348__CLK _5721_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3858__B1 _3919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_279_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4556__A _5765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4807__C1 _4791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5498__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3086__A1 _2850_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_310 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_243_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4338__A1 _4240_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4889__A2 _4874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3635__A _4303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3561__A2 _3597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3849__B1 _3848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3313__A2 _3318_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4510__A1 _5347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3190_ _5652_/Q _3147_/X _3149_/X _5572_/Q vssd1 vssd1 vccd1 vccd1 _3190_/X sky130_fd_sc_hd__a22o_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_210 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4466__A _4466_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_266_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3370__A _3419_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_205 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_281_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3077__A1 _2835_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_373 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4813__A2 _4799_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4913__B _4950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5762_ _5762_/A vssd1 vssd1 vccd1 vccd1 _5762_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_201_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2974_ _5397_/Q vssd1 vssd1 vccd1 vccd1 _2974_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4713_ _4722_/A _4981_/A vssd1 vssd1 vccd1 vccd1 _4713_/Y sky130_fd_sc_hd__nand2_1
XFILLER_277_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5693_ _5724_/CLK _5693_/D vssd1 vssd1 vccd1 vccd1 _5693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_212 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_277_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4329__A1 _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4644_ _5679_/Q vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__clkbuf_4
X_4575_ _5313_/A _5156_/A _4626_/S vssd1 vssd1 vccd1 vccd1 _4575_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3552__A2 _3948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3526_ _5347_/Q _5469_/Q _3761_/A _5291_/S vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__o31ai_4
XFILLER_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3457_ _3346_/B _3345_/A _3768_/S vssd1 vssd1 vccd1 vccd1 _3458_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__4079__C _4079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5760__A _5760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_130_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5640__CLK _5658_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3388_ _2840_/C _5374_/Q _3394_/S vssd1 vssd1 vccd1 vccd1 _3389_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5127_ _5747_/Q _3840_/A _5126_/X vssd1 vssd1 vccd1 vccd1 _5127_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_284_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5058_ _5051_/X _5052_/X _5054_/X _5056_/X _5071_/B vssd1 vssd1 vccd1 vccd1 _5058_/X
+ sky130_fd_sc_hd__o41a_1
XANTENNA__3068__A1 _5770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4009_ _4037_/A _4192_/A _4008_/X vssd1 vssd1 vccd1 vccd1 _4009_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_111_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_145 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_71_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_289 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4740__A1 _4679_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4179__S0 _4146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5296__A2 _3843_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input32_A i_req_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output119_A _5551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4733__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_188_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_178 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5513__CLK _5741_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2690_ _2690_/A vssd1 vssd1 vccd1 vccd1 _5319_/A sky130_fd_sc_hd__buf_6
XFILLER_184_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2990__B1 _2845_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4360_ _4347_/X _4350_/X _4359_/X _4232_/B _4438_/B vssd1 vssd1 vccd1 vccd1 _4499_/B
+ sky130_fd_sc_hd__o32a_4
XANTENNA__3534__A2 _4523_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5663__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2700__C _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3311_ _5373_/Q _3318_/C _3310_/X _5370_/Q _3293_/A vssd1 vssd1 vccd1 vccd1 _3311_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2742__B1 _2738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4291_ _4031_/X _4348_/B _4348_/C _4069_/C _4029_/X vssd1 vssd1 vccd1 vccd1 _4322_/B
+ sky130_fd_sc_hd__o311a_1
X_3242_ _5461_/Q _5094_/B _5094_/C vssd1 vssd1 vccd1 vccd1 _3989_/S sky130_fd_sc_hd__and3_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3173_ _5665_/Q _3137_/X _3139_/X _5585_/Q vssd1 vssd1 vccd1 vccd1 _3173_/X sky130_fd_sc_hd__a22o_1
XFILLER_239_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4247__A0 _4151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_287 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4798__A1 _5595_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2957_ _3799_/A _2957_/B vssd1 vssd1 vccd1 vccd1 _3283_/C sky130_fd_sc_hd__and2b_1
XANTENNA__3222__A1 _5562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5745_ _5747_/CLK _5745_/D vssd1 vssd1 vccd1 vccd1 _5745_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3773__A2 _3293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2888_ _3281_/A _3277_/A vssd1 vssd1 vccd1 vccd1 _2889_/B sky130_fd_sc_hd__or2_1
X_5676_ _5743_/CLK _5676_/D vssd1 vssd1 vccd1 vccd1 _5676_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2981__B1 _2840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4627_ _5526_/Q _4626_/X _5229_/S vssd1 vssd1 vccd1 vccd1 _4627_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_321 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4558_ _5766_/A _4560_/B vssd1 vssd1 vccd1 vccd1 _4577_/C sky130_fd_sc_hd__and2_1
XFILLER_237_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3509_ _5434_/Q input40/X _3517_/S vssd1 vssd1 vccd1 vccd1 _3510_/A sky130_fd_sc_hd__mux2_1
XFILLER_277_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4489_ _4617_/A _4617_/B _5200_/A vssd1 vssd1 vccd1 vccd1 _4491_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4486__B1 _4458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4834__A _4985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_313 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5536__CLK _5665_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_201_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_317 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_185_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3213__A1 _5673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3213__B2 _5593_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_278_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5686__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput62 _3217_/X vssd1 vssd1 vccd1 vccd1 dbg_out[13] sky130_fd_sc_hd__buf_2
XANTENNA__3913__A _5261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 _5767_/A vssd1 vssd1 vccd1 vccd1 dbg_out[23] sky130_fd_sc_hd__buf_2
Xoutput84 _5357_/Q vssd1 vssd1 vccd1 vccd1 dbg_out[33] sky130_fd_sc_hd__buf_2
Xoutput95 _5770_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[10] sky130_fd_sc_hd__buf_2
XANTENNA__3632__B _3673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4744__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_257 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3860_ _5473_/Q _3860_/B _5472_/Q vssd1 vssd1 vccd1 vccd1 _5055_/C sky130_fd_sc_hd__and3b_1
XANTENNA_clkbuf_leaf_7_i_clk_A clkbuf_2_2_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4182__C _4454_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2811_ _5342_/Q vssd1 vssd1 vccd1 vccd1 _3601_/B sky130_fd_sc_hd__buf_4
XANTENNA__3204__A1 _5607_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3791_ _3791_/A _3791_/B _3791_/C _3791_/D vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__or4_2
XFILLER_188_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _5692_/CLK _5530_/D vssd1 vssd1 vccd1 vccd1 _5530_/Q sky130_fd_sc_hd__dfxtp_4
X_2742_ _5554_/Q _2720_/B _2738_/X _2741_/X vssd1 vssd1 vccd1 vccd1 _3956_/A sky130_fd_sc_hd__o22ai_4
XFILLER_75_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5461_ _5721_/CLK _5461_/D vssd1 vssd1 vccd1 vccd1 _5461_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_157_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2673_ _5640_/Q _2655_/X _2657_/X _5672_/Q vssd1 vssd1 vccd1 vccd1 _2673_/X sky130_fd_sc_hd__a22o_1
XFILLER_184_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4412_ _4483_/B _4405_/A _4406_/Y _4322_/A vssd1 vssd1 vccd1 vccd1 _4413_/B sky130_fd_sc_hd__a31o_1
XFILLER_172_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5392_ _5404_/CLK _5392_/D vssd1 vssd1 vccd1 vccd1 _5392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2715__B1 _2664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4343_ _2919_/X _4030_/A _3692_/X _4063_/A _4342_/X vssd1 vssd1 vccd1 vccd1 _4343_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4919__A _5646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5409__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4274_ _4274_/A _4303_/A vssd1 vssd1 vccd1 vccd1 _4274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_207_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3225_ _5659_/Q _3147_/A _3149_/A _5579_/Q vssd1 vssd1 vccd1 vccd1 _3225_/X sky130_fd_sc_hd__a22o_1
XFILLER_223_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3140__B1 _3139_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3156_ _5629_/Q _3143_/X _3145_/X _3155_/X vssd1 vssd1 vccd1 vccd1 _3156_/X sky130_fd_sc_hd__a211o_1
XFILLER_254_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_223_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5559__CLK _5675_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_254_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4654__A _5549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3087_ _5774_/A _3063_/B _3085_/Y _3086_/X _3016_/A vssd1 vssd1 vccd1 vccd1 _3087_/X
+ sky130_fd_sc_hd__o221a_2
XFILLER_199_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4640__A0 _5720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _3988_/X _5325_/A _3989_/S vssd1 vssd1 vccd1 vccd1 _3990_/B sky130_fd_sc_hd__mux2_1
X_5728_ _5741_/CLK _5728_/D vssd1 vssd1 vccd1 vccd1 _5728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3717__B _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5659_ _5659_/CLK _5659_/D vssd1 vssd1 vccd1 vccd1 _5659_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2706__B1 _2657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_240 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_77_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2721__A3 _2719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_264_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_245_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3198__B1 _3139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3908__A _4635_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4934__A1 _5652_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3737__A2 _3605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output186_A _5484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3119__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4147__C1 _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2958__S _3337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4162__A2 _4050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4739__A _5570_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_11 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output63_A _3222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_273 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_268_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_203 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5111__A1 _4543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5701__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3010_ _3063_/B vssd1 vssd1 vccd1 vccd1 _3010_/X sky130_fd_sc_hd__buf_2
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4961_ _5664_/Q _4969_/A vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__or2_1
X_3912_ _5511_/Q _3245_/B _3245_/Y _5509_/Q vssd1 vssd1 vccd1 vccd1 _3913_/B sky130_fd_sc_hd__a22o_1
X_4892_ _5635_/Q _4894_/A vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__or2_1
XFILLER_232_391 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_189_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3843_ _5487_/Q _3843_/B _5294_/B vssd1 vssd1 vccd1 vccd1 _3843_/X sky130_fd_sc_hd__and3_1
XANTENNA__4921__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3189__B1 _3135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3728__A2 _3607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3774_ _4619_/B vssd1 vssd1 vccd1 vccd1 _5294_/A sky130_fd_sc_hd__clkbuf_4
X_5513_ _5741_/CLK _5513_/D vssd1 vssd1 vccd1 vccd1 _5513_/Q sky130_fd_sc_hd__dfxtp_1
X_2725_ _2775_/D _2775_/B _2727_/C _5571_/Q vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__and4bb_1
XFILLER_145_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5444_ _5692_/CLK _5444_/D vssd1 vssd1 vccd1 vccd1 _5444_/Q sky130_fd_sc_hd__dfxtp_1
X_2656_ _5344_/Q _5346_/Q _5345_/Q vssd1 vssd1 vccd1 vccd1 _2657_/A sky130_fd_sc_hd__and3_1
XFILLER_172_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5375_ _5441_/CLK _5375_/D vssd1 vssd1 vccd1 vccd1 _5375_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4649__A _5548_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5244__S _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4326_ _4326_/A _4326_/B vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__or2_1
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5381__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4257_ _4322_/A _4012_/X _4014_/X _4259_/B _4171_/A vssd1 vssd1 vccd1 vccd1 _4257_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_59_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_113_295 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_234_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4310__C1 _4161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3208_ _5672_/Q _3137_/A _3139_/A _5592_/Q vssd1 vssd1 vccd1 vccd1 _3208_/X sky130_fd_sc_hd__a22o_1
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4188_ _4322_/A _4055_/B _4169_/X _4171_/X _4187_/X vssd1 vssd1 vccd1 vccd1 _5200_/A
+ sky130_fd_sc_hd__o311a_4
XFILLER_67_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3139_ _3139_/A vssd1 vssd1 vccd1 vccd1 _3139_/X sky130_fd_sc_hd__buf_4
XFILLER_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5169__A1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2773__B_N _2789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4916__A1 _4646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2632__A _5345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_136_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4144__A2 _4059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5724__CLK _5724_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_345 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3352__A0 _2835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_389 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4278__B _4278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4993__S _5720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_265_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_319 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3655__A1 _5550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__A1 _4079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4383__A2 _4220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3490_ _5425_/Q input30/X _3496_/S vssd1 vssd1 vccd1 vccd1 _3491_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4469__A _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _5160_/A vssd1 vssd1 vccd1 vccd1 _5712_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4540__C1 _4529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4111_ _4368_/A _4370_/B _4368_/B vssd1 vssd1 vccd1 vccd1 _4111_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5091_ _3790_/X _4523_/B _5235_/S vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__a21o_1
XFILLER_271_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4042_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4043_/B sky130_fd_sc_hd__or2_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3646__A1 _4071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4932__A _4970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4944_ _5657_/Q _4935_/B _4943_/Y _4933_/X vssd1 vssd1 vccd1 vccd1 _5657_/D sky130_fd_sc_hd__o211a_1
XFILLER_33_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4875_ _5685_/Q _4950_/B vssd1 vssd1 vccd1 vccd1 _4894_/A sky130_fd_sc_hd__and2_4
XFILLER_32_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_177_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3826_ _5480_/Q _5384_/Q _3834_/S vssd1 vssd1 vccd1 vccd1 _3827_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3267__B _3267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3757_ _5067_/B _3755_/Y _4550_/S vssd1 vssd1 vccd1 vccd1 _3757_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5747__CLK _5747_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5763__A _5763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2708_ _2782_/C vssd1 vssd1 vccd1 vccd1 _2775_/B sky130_fd_sc_hd__buf_4
X_3688_ _5445_/Q _5449_/Q _5446_/Q _5444_/Q vssd1 vssd1 vccd1 vccd1 _3691_/A sky130_fd_sc_hd__or4_1
XFILLER_118_387 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_279_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2790__D1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4379__A _5445_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4126__A2 _4161_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5427_ _5441_/CLK _5427_/D vssd1 vssd1 vccd1 vccd1 _5427_/Q sky130_fd_sc_hd__dfxtp_1
X_2639_ _5344_/Q vssd1 vssd1 vccd1 vccd1 _2747_/D sky130_fd_sc_hd__buf_2
XFILLER_279_339 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_160_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5358_ _5724_/CLK _5358_/D vssd1 vssd1 vccd1 vccd1 _5358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_293 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4309_ _4306_/X _4230_/Y _4308_/Y vssd1 vssd1 vccd1 vccd1 _4309_/X sky130_fd_sc_hd__o21a_2
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5087__B1 _5077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5289_ _5292_/A _5289_/B vssd1 vssd1 vccd1 vccd1 _5290_/A sky130_fd_sc_hd__and2_1
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3637__A1 _5619_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4826__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3637__B2 _5603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4842__A _5613_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4062__A1 _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3458__A _5678_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5011__A0 _5687_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3892__S _3905_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3573__A0 _5484_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_365 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4770__C1 _4769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4117__A2 _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4289__A _4537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3325__B1 _3335_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_379 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2679__A2 _2644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3628__B2 _5600_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_253_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_352 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_206_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4589__C1 _3919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2990_ _2970_/Y _2850_/A _2845_/C _2988_/Y vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__a22o_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_282 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_202_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4660_ _4642_/Y _4658_/X _4659_/X _3986_/X vssd1 vssd1 vccd1 vccd1 _5550_/D sky130_fd_sc_hd__o211a_1
X_3611_ _5563_/Q _3596_/X _3604_/X _3610_/X vssd1 vssd1 vccd1 vccd1 _4484_/A sky130_fd_sc_hd__o22a_4
XANTENNA__4356__A2 _4067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4591_ _4613_/C vssd1 vssd1 vccd1 vccd1 _4604_/B sky130_fd_sc_hd__inv_2
XANTENNA__3564__B1 _3598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3542_ _4276_/A _4124_/B vssd1 vssd1 vccd1 vccd1 _4307_/B sky130_fd_sc_hd__nand2_2
XFILLER_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3473_ _5417_/Q input53/X _3475_/S vssd1 vssd1 vccd1 vccd1 _3474_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3316__B1 _3315_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5212_ _5717_/Q _5211_/X _5233_/S vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__mux2_1
XFILLER_276_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_215_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_372 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2943__A_N _3799_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5143_ _4496_/A _5142_/Y _5200_/B vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4927__A _5650_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5074_ _5513_/Q _3931_/A _5125_/A _5761_/A vssd1 vssd1 vccd1 vccd1 _5074_/X sky130_fd_sc_hd__a22o_1
XFILLER_284_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4025_ _4010_/X _4016_/X _4023_/X _4084_/B vssd1 vssd1 vccd1 vccd1 _4025_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4927_ _5650_/Q _4931_/A vssd1 vssd1 vccd1 vccd1 _4927_/X sky130_fd_sc_hd__or2_1
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4595__A2 _4490_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_309 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_230 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4858_ _5620_/Q _4859_/B _4857_/Y _4840_/X vssd1 vssd1 vccd1 vccd1 _5620_/D sky130_fd_sc_hd__o211a_1
XFILLER_165_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3809_ _5472_/Q _5376_/Q _3813_/S vssd1 vssd1 vccd1 vccd1 _3810_/A sky130_fd_sc_hd__mux2_1
X_4789_ _5591_/Q _4784_/B _4788_/Y _4769_/X vssd1 vssd1 vccd1 vccd1 _5591_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4752__C1 _4745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4837__A _5684_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4556__B _4581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4283__A1 _5450_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4283__B2 _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_322 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_203_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3619__C _4379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4338__A2 _4239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5299__A0 _5067_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3127__S _4651_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater214_A _5769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_258_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4510__A2 _5469_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4747__A _4972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_285_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_331 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5442__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4466__B _4466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3077__A2 _3089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3797__S _3813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5592__CLK _5659_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4482__A _4484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_179_349 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761_ _5761_/A vssd1 vssd1 vccd1 vccd1 _5761_/X sky130_fd_sc_hd__clkbuf_1
X_2973_ _5396_/Q vssd1 vssd1 vccd1 vccd1 _2973_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4712_ input11/X _4689_/X _4690_/X _4711_/Y vssd1 vssd1 vccd1 vccd1 _4981_/A sky130_fd_sc_hd__o2bb2a_4
XFILLER_187_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4982__C1 _4979_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5692_ _5692_/CLK _5692_/D vssd1 vssd1 vccd1 vccd1 _5692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4329__A2 _4033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4643_ input21/X input7/X _4651_/S vssd1 vssd1 vccd1 vccd1 _4643_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4734__C1 _4718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4574_ _5539_/Q _4511_/X _3919_/A _4573_/X vssd1 vssd1 vccd1 vccd1 _5539_/D sky130_fd_sc_hd__o211a_1
XFILLER_155_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3525_ _4987_/A _5331_/B vssd1 vssd1 vccd1 vccd1 _5442_/D sky130_fd_sc_hd__nor2_1
XFILLER_226_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_305 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3456_ _3456_/A vssd1 vssd1 vccd1 vccd1 _5407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_226_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3387_ _3387_/A vssd1 vssd1 vccd1 vccd1 _5373_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5126_ _5518_/Q _3931_/A _5082_/B _5498_/Q vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_284_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5057_ _5460_/Q vssd1 vssd1 vccd1 vccd1 _5071_/B sky130_fd_sc_hd__clkinv_2
XFILLER_242_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3068__A2 _3063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4008_ _4108_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _4008_/X sky130_fd_sc_hd__or2_1
XFILLER_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4973__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4740__A2 _4724_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5465__CLK _5743_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4179__S1 _4449_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4567__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3700__B1 _3606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A i_req_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_275_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4256__A1 _4281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_216_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_231_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4964__C1 _4957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output93_A _3197_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2700__D _5590_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2742__A1 _5554_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3310_ _3310_/A _3310_/B vssd1 vssd1 vccd1 vccd1 _3310_/X sky130_fd_sc_hd__or2_2
X_4290_ _4010_/X _4016_/X _4087_/A _4084_/B vssd1 vssd1 vccd1 vccd1 _4348_/C sky130_fd_sc_hd__o211a_1
XFILLER_112_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_i_clk_A clkbuf_2_0_0_i_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3241_ _5472_/Q _5473_/Q _3860_/B _5471_/Q vssd1 vssd1 vccd1 vccd1 _5094_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__3298__A2 _5366_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_112_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3172_ _5552_/Q _3131_/X _3169_/X _3171_/X vssd1 vssd1 vccd1 vccd1 _3172_/X sky130_fd_sc_hd__o22a_2
XFILLER_239_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_367 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4798__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_281_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__5338__CLK _5686_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5744_ _5747_/CLK _5744_/D vssd1 vssd1 vccd1 vccd1 _5744_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4955__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2956_ _2954_/X _5486_/D _2955_/X vssd1 vssd1 vccd1 vccd1 _5449_/D sky130_fd_sc_hd__o21a_1
XANTENNA__3222__A2 _3131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_5675_ _5675_/CLK _5675_/D vssd1 vssd1 vccd1 vccd1 _5675_/Q sky130_fd_sc_hd__dfxtp_2
X_2887_ _2949_/A _2922_/A vssd1 vssd1 vccd1 vccd1 _2928_/A sky130_fd_sc_hd__or2_2
XANTENNA__5247__S _5253_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3556__A _4030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4626_ _5325_/A _4457_/D _4626_/S vssd1 vssd1 vccd1 vccd1 _4626_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5488__CLK _5722_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_333 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_237_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4557_ _4529_/X _4555_/X _4556_/X _3919_/X vssd1 vssd1 vccd1 vccd1 _5537_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5771__A _5771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3508_ _3508_/A vssd1 vssd1 vccd1 vccd1 _5433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4488_ _5531_/Q _4458_/A _4485_/X _4486_/Y _4487_/X vssd1 vssd1 vccd1 vccd1 _5531_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3439_ _5399_/Q _3064_/X _3451_/S vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4486__A1 _3943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3694__C1 _3693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5109_ _5109_/A _5109_/B vssd1 vssd1 vccd1 vccd1 _5131_/A sky130_fd_sc_hd__or2_1
XFILLER_245_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4789__A2 _4784_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4834__B _4834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4850__A _5617_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4946__C1 _4933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_297 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3213__A2 _3137_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_138 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4174__B1 _4471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput63 _3222_/X vssd1 vssd1 vccd1 vccd1 dbg_out[14] sky130_fd_sc_hd__buf_2
Xoutput74 _5768_/A vssd1 vssd1 vccd1 vccd1 dbg_out[24] sky130_fd_sc_hd__buf_2
XFILLER_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 _3458_/C vssd1 vssd1 vccd1 vccd1 dbg_out[34] sky130_fd_sc_hd__buf_2
XANTENNA__4477__A1 _5529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput96 _5771_/X vssd1 vssd1 vccd1 vccd1 dbg_pc[11] sky130_fd_sc_hd__buf_2
XANTENNA__3405__S _3415_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4744__B _4747_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3988__A0 _5774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_337 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2810_ _5343_/Q vssd1 vssd1 vccd1 vccd1 _3599_/B sky130_fd_sc_hd__buf_4
XFILLER_176_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3204__A2 _3133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3790_ _5464_/Q vssd1 vssd1 vccd1 vccd1 _3790_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_176_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5630__CLK _5653_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _5586_/Q _2635_/Y _2686_/X _2739_/X _2740_/X vssd1 vssd1 vccd1 vccd1 _2741_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_191_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5460_ _5707_/CLK _5460_/D vssd1 vssd1 vccd1 vccd1 _5460_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2672_ _5576_/Q _2644_/X _2664_/X _5608_/Q vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__a22o_1
XFILLER_274_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4165__B1 _4159_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4411_ _4405_/A _4406_/Y _4483_/B vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__a21oi_1
X_5391_ _5404_/CLK _5391_/D vssd1 vssd1 vccd1 vccd1 _5391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_377 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2715__A1 _5572_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2715__B2 _5604_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ _4030_/A _4063_/A _5452_/Q vssd1 vssd1 vccd1 vccd1 _4342_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4919__B _4947_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5741__D _5741_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4273_ _4231_/X _4272_/X _4304_/S vssd1 vssd1 vccd1 vccd1 _4273_/X sky130_fd_sc_hd__mux2_1
XANTENNA__2684__A_N _2757_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3224_ _5611_/Q _3133_/A _3135_/A _5627_/Q _3223_/X vssd1 vssd1 vccd1 vccd1 _3224_/X
+ sky130_fd_sc_hd__a221o_1
.ends

