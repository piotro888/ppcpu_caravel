VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO interconnect_inner
  CLASS BLOCK ;
  FOREIGN interconnect_inner ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 350.000 ;
  PIN c0_dbg_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END c0_dbg_pc[0]
  PIN c0_dbg_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 4.000 ;
    END
  END c0_dbg_pc[10]
  PIN c0_dbg_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 374.080 0.000 374.640 4.000 ;
    END
  END c0_dbg_pc[11]
  PIN c0_dbg_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 0.000 397.040 4.000 ;
    END
  END c0_dbg_pc[12]
  PIN c0_dbg_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END c0_dbg_pc[13]
  PIN c0_dbg_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 441.280 0.000 441.840 4.000 ;
    END
  END c0_dbg_pc[14]
  PIN c0_dbg_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 0.000 464.240 4.000 ;
    END
  END c0_dbg_pc[15]
  PIN c0_dbg_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END c0_dbg_pc[1]
  PIN c0_dbg_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 0.000 146.160 4.000 ;
    END
  END c0_dbg_pc[2]
  PIN c0_dbg_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 0.000 173.040 4.000 ;
    END
  END c0_dbg_pc[3]
  PIN c0_dbg_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 199.360 0.000 199.920 4.000 ;
    END
  END c0_dbg_pc[4]
  PIN c0_dbg_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END c0_dbg_pc[5]
  PIN c0_dbg_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 253.120 0.000 253.680 4.000 ;
    END
  END c0_dbg_pc[6]
  PIN c0_dbg_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END c0_dbg_pc[7]
  PIN c0_dbg_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.880 0.000 307.440 4.000 ;
    END
  END c0_dbg_pc[8]
  PIN c0_dbg_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 0.000 329.840 4.000 ;
    END
  END c0_dbg_pc[9]
  PIN c0_dbg_r0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END c0_dbg_r0[0]
  PIN c0_dbg_r0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 0.000 354.480 4.000 ;
    END
  END c0_dbg_r0[10]
  PIN c0_dbg_r0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 0.000 376.880 4.000 ;
    END
  END c0_dbg_r0[11]
  PIN c0_dbg_r0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 0.000 399.280 4.000 ;
    END
  END c0_dbg_r0[12]
  PIN c0_dbg_r0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 0.000 421.680 4.000 ;
    END
  END c0_dbg_r0[13]
  PIN c0_dbg_r0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 0.000 444.080 4.000 ;
    END
  END c0_dbg_r0[14]
  PIN c0_dbg_r0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 465.920 0.000 466.480 4.000 ;
    END
  END c0_dbg_r0[15]
  PIN c0_dbg_r0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.720 0.000 119.280 4.000 ;
    END
  END c0_dbg_r0[1]
  PIN c0_dbg_r0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END c0_dbg_r0[2]
  PIN c0_dbg_r0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 0.000 175.280 4.000 ;
    END
  END c0_dbg_r0[3]
  PIN c0_dbg_r0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 0.000 202.160 4.000 ;
    END
  END c0_dbg_r0[4]
  PIN c0_dbg_r0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 0.000 229.040 4.000 ;
    END
  END c0_dbg_r0[5]
  PIN c0_dbg_r0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END c0_dbg_r0[6]
  PIN c0_dbg_r0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 0.000 282.800 4.000 ;
    END
  END c0_dbg_r0[7]
  PIN c0_dbg_r0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 0.000 309.680 4.000 ;
    END
  END c0_dbg_r0[8]
  PIN c0_dbg_r0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 0.000 332.080 4.000 ;
    END
  END c0_dbg_r0[9]
  PIN c0_disable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END c0_disable
  PIN c0_i_core_int_sreg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.840 0.000 92.400 4.000 ;
    END
  END c0_i_core_int_sreg[0]
  PIN c0_i_core_int_sreg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 0.000 356.720 4.000 ;
    END
  END c0_i_core_int_sreg[10]
  PIN c0_i_core_int_sreg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END c0_i_core_int_sreg[11]
  PIN c0_i_core_int_sreg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END c0_i_core_int_sreg[12]
  PIN c0_i_core_int_sreg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 0.000 423.920 4.000 ;
    END
  END c0_i_core_int_sreg[13]
  PIN c0_i_core_int_sreg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 0.000 446.320 4.000 ;
    END
  END c0_i_core_int_sreg[14]
  PIN c0_i_core_int_sreg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 0.000 468.720 4.000 ;
    END
  END c0_i_core_int_sreg[15]
  PIN c0_i_core_int_sreg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 0.000 121.520 4.000 ;
    END
  END c0_i_core_int_sreg[1]
  PIN c0_i_core_int_sreg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 4.000 ;
    END
  END c0_i_core_int_sreg[2]
  PIN c0_i_core_int_sreg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END c0_i_core_int_sreg[3]
  PIN c0_i_core_int_sreg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 0.000 204.400 4.000 ;
    END
  END c0_i_core_int_sreg[4]
  PIN c0_i_core_int_sreg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 4.000 ;
    END
  END c0_i_core_int_sreg[5]
  PIN c0_i_core_int_sreg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END c0_i_core_int_sreg[6]
  PIN c0_i_core_int_sreg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END c0_i_core_int_sreg[7]
  PIN c0_i_core_int_sreg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 4.000 ;
    END
  END c0_i_core_int_sreg[8]
  PIN c0_i_core_int_sreg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 333.760 0.000 334.320 4.000 ;
    END
  END c0_i_core_int_sreg[9]
  PIN c0_i_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END c0_i_irq
  PIN c0_i_mc_core_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END c0_i_mc_core_int
  PIN c0_i_mem_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END c0_i_mem_ack
  PIN c0_i_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END c0_i_mem_data[0]
  PIN c0_i_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 358.400 0.000 358.960 4.000 ;
    END
  END c0_i_mem_data[10]
  PIN c0_i_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 0.000 381.360 4.000 ;
    END
  END c0_i_mem_data[11]
  PIN c0_i_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 0.000 403.760 4.000 ;
    END
  END c0_i_mem_data[12]
  PIN c0_i_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 0.000 426.160 4.000 ;
    END
  END c0_i_mem_data[13]
  PIN c0_i_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 0.000 448.560 4.000 ;
    END
  END c0_i_mem_data[14]
  PIN c0_i_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 0.000 470.960 4.000 ;
    END
  END c0_i_mem_data[15]
  PIN c0_i_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END c0_i_mem_data[1]
  PIN c0_i_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 0.000 152.880 4.000 ;
    END
  END c0_i_mem_data[2]
  PIN c0_i_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END c0_i_mem_data[3]
  PIN c0_i_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 0.000 206.640 4.000 ;
    END
  END c0_i_mem_data[4]
  PIN c0_i_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 0.000 233.520 4.000 ;
    END
  END c0_i_mem_data[5]
  PIN c0_i_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 0.000 260.400 4.000 ;
    END
  END c0_i_mem_data[6]
  PIN c0_i_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END c0_i_mem_data[7]
  PIN c0_i_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END c0_i_mem_data[8]
  PIN c0_i_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 0.000 336.560 4.000 ;
    END
  END c0_i_mem_data[9]
  PIN c0_i_mem_exception
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END c0_i_mem_exception
  PIN c0_i_req_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END c0_i_req_data[0]
  PIN c0_i_req_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 0.000 361.200 4.000 ;
    END
  END c0_i_req_data[10]
  PIN c0_i_req_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 0.000 383.600 4.000 ;
    END
  END c0_i_req_data[11]
  PIN c0_i_req_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 0.000 406.000 4.000 ;
    END
  END c0_i_req_data[12]
  PIN c0_i_req_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 427.840 0.000 428.400 4.000 ;
    END
  END c0_i_req_data[13]
  PIN c0_i_req_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 0.000 450.800 4.000 ;
    END
  END c0_i_req_data[14]
  PIN c0_i_req_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 0.000 473.200 4.000 ;
    END
  END c0_i_req_data[15]
  PIN c0_i_req_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 0.000 486.640 4.000 ;
    END
  END c0_i_req_data[16]
  PIN c0_i_req_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 0.000 488.880 4.000 ;
    END
  END c0_i_req_data[17]
  PIN c0_i_req_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 0.000 491.120 4.000 ;
    END
  END c0_i_req_data[18]
  PIN c0_i_req_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 492.800 0.000 493.360 4.000 ;
    END
  END c0_i_req_data[19]
  PIN c0_i_req_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END c0_i_req_data[1]
  PIN c0_i_req_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 495.040 0.000 495.600 4.000 ;
    END
  END c0_i_req_data[20]
  PIN c0_i_req_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 0.000 497.840 4.000 ;
    END
  END c0_i_req_data[21]
  PIN c0_i_req_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END c0_i_req_data[22]
  PIN c0_i_req_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 501.760 0.000 502.320 4.000 ;
    END
  END c0_i_req_data[23]
  PIN c0_i_req_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 0.000 504.560 4.000 ;
    END
  END c0_i_req_data[24]
  PIN c0_i_req_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 506.240 0.000 506.800 4.000 ;
    END
  END c0_i_req_data[25]
  PIN c0_i_req_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 508.480 0.000 509.040 4.000 ;
    END
  END c0_i_req_data[26]
  PIN c0_i_req_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 0.000 511.280 4.000 ;
    END
  END c0_i_req_data[27]
  PIN c0_i_req_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 0.000 513.520 4.000 ;
    END
  END c0_i_req_data[28]
  PIN c0_i_req_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 0.000 515.760 4.000 ;
    END
  END c0_i_req_data[29]
  PIN c0_i_req_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END c0_i_req_data[2]
  PIN c0_i_req_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 0.000 518.000 4.000 ;
    END
  END c0_i_req_data[30]
  PIN c0_i_req_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 0.000 520.240 4.000 ;
    END
  END c0_i_req_data[31]
  PIN c0_i_req_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 0.000 182.000 4.000 ;
    END
  END c0_i_req_data[3]
  PIN c0_i_req_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 0.000 208.880 4.000 ;
    END
  END c0_i_req_data[4]
  PIN c0_i_req_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 0.000 235.760 4.000 ;
    END
  END c0_i_req_data[5]
  PIN c0_i_req_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 0.000 262.640 4.000 ;
    END
  END c0_i_req_data[6]
  PIN c0_i_req_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 0.000 289.520 4.000 ;
    END
  END c0_i_req_data[7]
  PIN c0_i_req_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 0.000 316.400 4.000 ;
    END
  END c0_i_req_data[8]
  PIN c0_i_req_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 4.000 ;
    END
  END c0_i_req_data[9]
  PIN c0_i_req_data_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END c0_i_req_data_valid
  PIN c0_o_c_data_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 4.000 ;
    END
  END c0_o_c_data_page
  PIN c0_o_c_instr_long
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 64.960 0.000 65.520 4.000 ;
    END
  END c0_o_c_instr_long
  PIN c0_o_c_instr_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END c0_o_c_instr_page
  PIN c0_o_icache_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END c0_o_icache_flush
  PIN c0_o_instr_long_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END c0_o_instr_long_addr[0]
  PIN c0_o_instr_long_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 4.000 ;
    END
  END c0_o_instr_long_addr[1]
  PIN c0_o_instr_long_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 0.000 157.360 4.000 ;
    END
  END c0_o_instr_long_addr[2]
  PIN c0_o_instr_long_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 0.000 184.240 4.000 ;
    END
  END c0_o_instr_long_addr[3]
  PIN c0_o_instr_long_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 0.000 211.120 4.000 ;
    END
  END c0_o_instr_long_addr[4]
  PIN c0_o_instr_long_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 0.000 238.000 4.000 ;
    END
  END c0_o_instr_long_addr[5]
  PIN c0_o_instr_long_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 0.000 264.880 4.000 ;
    END
  END c0_o_instr_long_addr[6]
  PIN c0_o_instr_long_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 0.000 291.760 4.000 ;
    END
  END c0_o_instr_long_addr[7]
  PIN c0_o_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END c0_o_mem_addr[0]
  PIN c0_o_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 0.000 363.440 4.000 ;
    END
  END c0_o_mem_addr[10]
  PIN c0_o_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 385.280 0.000 385.840 4.000 ;
    END
  END c0_o_mem_addr[11]
  PIN c0_o_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 0.000 408.240 4.000 ;
    END
  END c0_o_mem_addr[12]
  PIN c0_o_mem_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 0.000 430.640 4.000 ;
    END
  END c0_o_mem_addr[13]
  PIN c0_o_mem_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 452.480 0.000 453.040 4.000 ;
    END
  END c0_o_mem_addr[14]
  PIN c0_o_mem_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 474.880 0.000 475.440 4.000 ;
    END
  END c0_o_mem_addr[15]
  PIN c0_o_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 0.000 130.480 4.000 ;
    END
  END c0_o_mem_addr[1]
  PIN c0_o_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 159.040 0.000 159.600 4.000 ;
    END
  END c0_o_mem_addr[2]
  PIN c0_o_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 185.920 0.000 186.480 4.000 ;
    END
  END c0_o_mem_addr[3]
  PIN c0_o_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 0.000 213.360 4.000 ;
    END
  END c0_o_mem_addr[4]
  PIN c0_o_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 239.680 0.000 240.240 4.000 ;
    END
  END c0_o_mem_addr[5]
  PIN c0_o_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 0.000 267.120 4.000 ;
    END
  END c0_o_mem_addr[6]
  PIN c0_o_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 293.440 0.000 294.000 4.000 ;
    END
  END c0_o_mem_addr[7]
  PIN c0_o_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 0.000 318.640 4.000 ;
    END
  END c0_o_mem_addr[8]
  PIN c0_o_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END c0_o_mem_addr[9]
  PIN c0_o_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 0.000 103.600 4.000 ;
    END
  END c0_o_mem_data[0]
  PIN c0_o_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 0.000 365.680 4.000 ;
    END
  END c0_o_mem_data[10]
  PIN c0_o_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 387.520 0.000 388.080 4.000 ;
    END
  END c0_o_mem_data[11]
  PIN c0_o_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 0.000 410.480 4.000 ;
    END
  END c0_o_mem_data[12]
  PIN c0_o_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 0.000 432.880 4.000 ;
    END
  END c0_o_mem_data[13]
  PIN c0_o_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 454.720 0.000 455.280 4.000 ;
    END
  END c0_o_mem_data[14]
  PIN c0_o_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 0.000 477.680 4.000 ;
    END
  END c0_o_mem_data[15]
  PIN c0_o_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 132.160 0.000 132.720 4.000 ;
    END
  END c0_o_mem_data[1]
  PIN c0_o_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 0.000 161.840 4.000 ;
    END
  END c0_o_mem_data[2]
  PIN c0_o_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 0.000 188.720 4.000 ;
    END
  END c0_o_mem_data[3]
  PIN c0_o_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END c0_o_mem_data[4]
  PIN c0_o_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 0.000 242.480 4.000 ;
    END
  END c0_o_mem_data[5]
  PIN c0_o_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 0.000 269.360 4.000 ;
    END
  END c0_o_mem_data[6]
  PIN c0_o_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 0.000 296.240 4.000 ;
    END
  END c0_o_mem_data[7]
  PIN c0_o_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 0.000 320.880 4.000 ;
    END
  END c0_o_mem_data[8]
  PIN c0_o_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 0.000 343.280 4.000 ;
    END
  END c0_o_mem_data[9]
  PIN c0_o_mem_high_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 105.280 0.000 105.840 4.000 ;
    END
  END c0_o_mem_high_addr[0]
  PIN c0_o_mem_high_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END c0_o_mem_high_addr[1]
  PIN c0_o_mem_high_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 0.000 164.080 4.000 ;
    END
  END c0_o_mem_high_addr[2]
  PIN c0_o_mem_high_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END c0_o_mem_high_addr[3]
  PIN c0_o_mem_high_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END c0_o_mem_high_addr[4]
  PIN c0_o_mem_high_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END c0_o_mem_high_addr[5]
  PIN c0_o_mem_high_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 0.000 271.600 4.000 ;
    END
  END c0_o_mem_high_addr[6]
  PIN c0_o_mem_high_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 0.000 298.480 4.000 ;
    END
  END c0_o_mem_high_addr[7]
  PIN c0_o_mem_long_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 4.000 ;
    END
  END c0_o_mem_long_mode
  PIN c0_o_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END c0_o_mem_req
  PIN c0_o_mem_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END c0_o_mem_sel[0]
  PIN c0_o_mem_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END c0_o_mem_sel[1]
  PIN c0_o_mem_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END c0_o_mem_we
  PIN c0_o_req_active
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 0.000 78.960 4.000 ;
    END
  END c0_o_req_active
  PIN c0_o_req_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END c0_o_req_addr[0]
  PIN c0_o_req_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 0.000 367.920 4.000 ;
    END
  END c0_o_req_addr[10]
  PIN c0_o_req_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 0.000 390.320 4.000 ;
    END
  END c0_o_req_addr[11]
  PIN c0_o_req_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 412.160 0.000 412.720 4.000 ;
    END
  END c0_o_req_addr[12]
  PIN c0_o_req_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 0.000 435.120 4.000 ;
    END
  END c0_o_req_addr[13]
  PIN c0_o_req_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 0.000 457.520 4.000 ;
    END
  END c0_o_req_addr[14]
  PIN c0_o_req_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 0.000 479.920 4.000 ;
    END
  END c0_o_req_addr[15]
  PIN c0_o_req_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END c0_o_req_addr[1]
  PIN c0_o_req_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 0.000 166.320 4.000 ;
    END
  END c0_o_req_addr[2]
  PIN c0_o_req_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END c0_o_req_addr[3]
  PIN c0_o_req_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 0.000 220.080 4.000 ;
    END
  END c0_o_req_addr[4]
  PIN c0_o_req_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END c0_o_req_addr[5]
  PIN c0_o_req_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 0.000 273.840 4.000 ;
    END
  END c0_o_req_addr[6]
  PIN c0_o_req_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 0.000 300.720 4.000 ;
    END
  END c0_o_req_addr[7]
  PIN c0_o_req_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 0.000 323.120 4.000 ;
    END
  END c0_o_req_addr[8]
  PIN c0_o_req_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 0.000 345.520 4.000 ;
    END
  END c0_o_req_addr[9]
  PIN c0_o_req_ppl_submit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END c0_o_req_ppl_submit
  PIN c0_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END c0_rst
  PIN c0_sr_bus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END c0_sr_bus_addr[0]
  PIN c0_sr_bus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 0.000 370.160 4.000 ;
    END
  END c0_sr_bus_addr[10]
  PIN c0_sr_bus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 0.000 392.560 4.000 ;
    END
  END c0_sr_bus_addr[11]
  PIN c0_sr_bus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END c0_sr_bus_addr[12]
  PIN c0_sr_bus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 0.000 437.360 4.000 ;
    END
  END c0_sr_bus_addr[13]
  PIN c0_sr_bus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END c0_sr_bus_addr[14]
  PIN c0_sr_bus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 0.000 482.160 4.000 ;
    END
  END c0_sr_bus_addr[15]
  PIN c0_sr_bus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 0.000 141.680 4.000 ;
    END
  END c0_sr_bus_addr[1]
  PIN c0_sr_bus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END c0_sr_bus_addr[2]
  PIN c0_sr_bus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END c0_sr_bus_addr[3]
  PIN c0_sr_bus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 0.000 222.320 4.000 ;
    END
  END c0_sr_bus_addr[4]
  PIN c0_sr_bus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 0.000 249.200 4.000 ;
    END
  END c0_sr_bus_addr[5]
  PIN c0_sr_bus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 0.000 276.080 4.000 ;
    END
  END c0_sr_bus_addr[6]
  PIN c0_sr_bus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 0.000 302.960 4.000 ;
    END
  END c0_sr_bus_addr[7]
  PIN c0_sr_bus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END c0_sr_bus_addr[8]
  PIN c0_sr_bus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 0.000 347.760 4.000 ;
    END
  END c0_sr_bus_addr[9]
  PIN c0_sr_bus_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END c0_sr_bus_data_o[0]
  PIN c0_sr_bus_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 0.000 372.400 4.000 ;
    END
  END c0_sr_bus_data_o[10]
  PIN c0_sr_bus_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 0.000 394.800 4.000 ;
    END
  END c0_sr_bus_data_o[11]
  PIN c0_sr_bus_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 0.000 417.200 4.000 ;
    END
  END c0_sr_bus_data_o[12]
  PIN c0_sr_bus_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 0.000 439.600 4.000 ;
    END
  END c0_sr_bus_data_o[13]
  PIN c0_sr_bus_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 0.000 462.000 4.000 ;
    END
  END c0_sr_bus_data_o[14]
  PIN c0_sr_bus_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 0.000 484.400 4.000 ;
    END
  END c0_sr_bus_data_o[15]
  PIN c0_sr_bus_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 0.000 143.920 4.000 ;
    END
  END c0_sr_bus_data_o[1]
  PIN c0_sr_bus_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 0.000 170.800 4.000 ;
    END
  END c0_sr_bus_data_o[2]
  PIN c0_sr_bus_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 4.000 ;
    END
  END c0_sr_bus_data_o[3]
  PIN c0_sr_bus_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 0.000 224.560 4.000 ;
    END
  END c0_sr_bus_data_o[4]
  PIN c0_sr_bus_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 0.000 251.440 4.000 ;
    END
  END c0_sr_bus_data_o[5]
  PIN c0_sr_bus_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 0.000 278.320 4.000 ;
    END
  END c0_sr_bus_data_o[6]
  PIN c0_sr_bus_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 0.000 305.200 4.000 ;
    END
  END c0_sr_bus_data_o[7]
  PIN c0_sr_bus_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 0.000 327.600 4.000 ;
    END
  END c0_sr_bus_data_o[8]
  PIN c0_sr_bus_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 0.000 350.000 4.000 ;
    END
  END c0_sr_bus_data_o[9]
  PIN c0_sr_bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END c0_sr_bus_we
  PIN c1_dbg_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 716.800 0.000 717.360 4.000 ;
    END
  END c1_dbg_pc[0]
  PIN c1_dbg_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 0.000 981.680 4.000 ;
    END
  END c1_dbg_pc[10]
  PIN c1_dbg_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1003.520 0.000 1004.080 4.000 ;
    END
  END c1_dbg_pc[11]
  PIN c1_dbg_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1025.920 0.000 1026.480 4.000 ;
    END
  END c1_dbg_pc[12]
  PIN c1_dbg_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1048.320 0.000 1048.880 4.000 ;
    END
  END c1_dbg_pc[13]
  PIN c1_dbg_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1070.720 0.000 1071.280 4.000 ;
    END
  END c1_dbg_pc[14]
  PIN c1_dbg_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1093.120 0.000 1093.680 4.000 ;
    END
  END c1_dbg_pc[15]
  PIN c1_dbg_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 0.000 746.480 4.000 ;
    END
  END c1_dbg_pc[1]
  PIN c1_dbg_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 775.040 0.000 775.600 4.000 ;
    END
  END c1_dbg_pc[2]
  PIN c1_dbg_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 0.000 802.480 4.000 ;
    END
  END c1_dbg_pc[3]
  PIN c1_dbg_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 828.800 0.000 829.360 4.000 ;
    END
  END c1_dbg_pc[4]
  PIN c1_dbg_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 855.680 0.000 856.240 4.000 ;
    END
  END c1_dbg_pc[5]
  PIN c1_dbg_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 882.560 0.000 883.120 4.000 ;
    END
  END c1_dbg_pc[6]
  PIN c1_dbg_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 909.440 0.000 910.000 4.000 ;
    END
  END c1_dbg_pc[7]
  PIN c1_dbg_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 936.320 0.000 936.880 4.000 ;
    END
  END c1_dbg_pc[8]
  PIN c1_dbg_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 958.720 0.000 959.280 4.000 ;
    END
  END c1_dbg_pc[9]
  PIN c1_dbg_r0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 0.000 719.600 4.000 ;
    END
  END c1_dbg_r0[0]
  PIN c1_dbg_r0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 0.000 983.920 4.000 ;
    END
  END c1_dbg_r0[10]
  PIN c1_dbg_r0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1005.760 0.000 1006.320 4.000 ;
    END
  END c1_dbg_r0[11]
  PIN c1_dbg_r0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 0.000 1028.720 4.000 ;
    END
  END c1_dbg_r0[12]
  PIN c1_dbg_r0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1050.560 0.000 1051.120 4.000 ;
    END
  END c1_dbg_r0[13]
  PIN c1_dbg_r0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1072.960 0.000 1073.520 4.000 ;
    END
  END c1_dbg_r0[14]
  PIN c1_dbg_r0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1095.360 0.000 1095.920 4.000 ;
    END
  END c1_dbg_r0[15]
  PIN c1_dbg_r0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 748.160 0.000 748.720 4.000 ;
    END
  END c1_dbg_r0[1]
  PIN c1_dbg_r0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 777.280 0.000 777.840 4.000 ;
    END
  END c1_dbg_r0[2]
  PIN c1_dbg_r0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 804.160 0.000 804.720 4.000 ;
    END
  END c1_dbg_r0[3]
  PIN c1_dbg_r0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 831.040 0.000 831.600 4.000 ;
    END
  END c1_dbg_r0[4]
  PIN c1_dbg_r0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 857.920 0.000 858.480 4.000 ;
    END
  END c1_dbg_r0[5]
  PIN c1_dbg_r0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 884.800 0.000 885.360 4.000 ;
    END
  END c1_dbg_r0[6]
  PIN c1_dbg_r0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 911.680 0.000 912.240 4.000 ;
    END
  END c1_dbg_r0[7]
  PIN c1_dbg_r0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 938.560 0.000 939.120 4.000 ;
    END
  END c1_dbg_r0[8]
  PIN c1_dbg_r0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 0.000 961.520 4.000 ;
    END
  END c1_dbg_r0[9]
  PIN c1_disable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 0.000 679.280 4.000 ;
    END
  END c1_disable
  PIN c1_i_core_int_sreg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 721.280 0.000 721.840 4.000 ;
    END
  END c1_i_core_int_sreg[0]
  PIN c1_i_core_int_sreg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 985.600 0.000 986.160 4.000 ;
    END
  END c1_i_core_int_sreg[10]
  PIN c1_i_core_int_sreg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1008.000 0.000 1008.560 4.000 ;
    END
  END c1_i_core_int_sreg[11]
  PIN c1_i_core_int_sreg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1030.400 0.000 1030.960 4.000 ;
    END
  END c1_i_core_int_sreg[12]
  PIN c1_i_core_int_sreg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1052.800 0.000 1053.360 4.000 ;
    END
  END c1_i_core_int_sreg[13]
  PIN c1_i_core_int_sreg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1075.200 0.000 1075.760 4.000 ;
    END
  END c1_i_core_int_sreg[14]
  PIN c1_i_core_int_sreg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1097.600 0.000 1098.160 4.000 ;
    END
  END c1_i_core_int_sreg[15]
  PIN c1_i_core_int_sreg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 750.400 0.000 750.960 4.000 ;
    END
  END c1_i_core_int_sreg[1]
  PIN c1_i_core_int_sreg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 0.000 780.080 4.000 ;
    END
  END c1_i_core_int_sreg[2]
  PIN c1_i_core_int_sreg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 806.400 0.000 806.960 4.000 ;
    END
  END c1_i_core_int_sreg[3]
  PIN c1_i_core_int_sreg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 833.280 0.000 833.840 4.000 ;
    END
  END c1_i_core_int_sreg[4]
  PIN c1_i_core_int_sreg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 0.000 860.720 4.000 ;
    END
  END c1_i_core_int_sreg[5]
  PIN c1_i_core_int_sreg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 0.000 887.600 4.000 ;
    END
  END c1_i_core_int_sreg[6]
  PIN c1_i_core_int_sreg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 0.000 914.480 4.000 ;
    END
  END c1_i_core_int_sreg[7]
  PIN c1_i_core_int_sreg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 940.800 0.000 941.360 4.000 ;
    END
  END c1_i_core_int_sreg[8]
  PIN c1_i_core_int_sreg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 963.200 0.000 963.760 4.000 ;
    END
  END c1_i_core_int_sreg[9]
  PIN c1_i_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 0.000 681.520 4.000 ;
    END
  END c1_i_irq
  PIN c1_i_mc_core_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 683.200 0.000 683.760 4.000 ;
    END
  END c1_i_mc_core_int
  PIN c1_i_mem_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 0.000 686.000 4.000 ;
    END
  END c1_i_mem_ack
  PIN c1_i_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 723.520 0.000 724.080 4.000 ;
    END
  END c1_i_mem_data[0]
  PIN c1_i_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 987.840 0.000 988.400 4.000 ;
    END
  END c1_i_mem_data[10]
  PIN c1_i_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1010.240 0.000 1010.800 4.000 ;
    END
  END c1_i_mem_data[11]
  PIN c1_i_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1032.640 0.000 1033.200 4.000 ;
    END
  END c1_i_mem_data[12]
  PIN c1_i_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1055.040 0.000 1055.600 4.000 ;
    END
  END c1_i_mem_data[13]
  PIN c1_i_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1077.440 0.000 1078.000 4.000 ;
    END
  END c1_i_mem_data[14]
  PIN c1_i_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1099.840 0.000 1100.400 4.000 ;
    END
  END c1_i_mem_data[15]
  PIN c1_i_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 0.000 753.200 4.000 ;
    END
  END c1_i_mem_data[1]
  PIN c1_i_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 0.000 782.320 4.000 ;
    END
  END c1_i_mem_data[2]
  PIN c1_i_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 0.000 809.200 4.000 ;
    END
  END c1_i_mem_data[3]
  PIN c1_i_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 835.520 0.000 836.080 4.000 ;
    END
  END c1_i_mem_data[4]
  PIN c1_i_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END c1_i_mem_data[5]
  PIN c1_i_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 889.280 0.000 889.840 4.000 ;
    END
  END c1_i_mem_data[6]
  PIN c1_i_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 916.160 0.000 916.720 4.000 ;
    END
  END c1_i_mem_data[7]
  PIN c1_i_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 943.040 0.000 943.600 4.000 ;
    END
  END c1_i_mem_data[8]
  PIN c1_i_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 965.440 0.000 966.000 4.000 ;
    END
  END c1_i_mem_data[9]
  PIN c1_i_mem_exception
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 0.000 688.240 4.000 ;
    END
  END c1_i_mem_exception
  PIN c1_i_req_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 0.000 726.320 4.000 ;
    END
  END c1_i_req_data[0]
  PIN c1_i_req_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 990.080 0.000 990.640 4.000 ;
    END
  END c1_i_req_data[10]
  PIN c1_i_req_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1012.480 0.000 1013.040 4.000 ;
    END
  END c1_i_req_data[11]
  PIN c1_i_req_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1034.880 0.000 1035.440 4.000 ;
    END
  END c1_i_req_data[12]
  PIN c1_i_req_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1057.280 0.000 1057.840 4.000 ;
    END
  END c1_i_req_data[13]
  PIN c1_i_req_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1079.680 0.000 1080.240 4.000 ;
    END
  END c1_i_req_data[14]
  PIN c1_i_req_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1102.080 0.000 1102.640 4.000 ;
    END
  END c1_i_req_data[15]
  PIN c1_i_req_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1115.520 0.000 1116.080 4.000 ;
    END
  END c1_i_req_data[16]
  PIN c1_i_req_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1117.760 0.000 1118.320 4.000 ;
    END
  END c1_i_req_data[17]
  PIN c1_i_req_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1120.000 0.000 1120.560 4.000 ;
    END
  END c1_i_req_data[18]
  PIN c1_i_req_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1122.240 0.000 1122.800 4.000 ;
    END
  END c1_i_req_data[19]
  PIN c1_i_req_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 754.880 0.000 755.440 4.000 ;
    END
  END c1_i_req_data[1]
  PIN c1_i_req_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1124.480 0.000 1125.040 4.000 ;
    END
  END c1_i_req_data[20]
  PIN c1_i_req_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1126.720 0.000 1127.280 4.000 ;
    END
  END c1_i_req_data[21]
  PIN c1_i_req_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1128.960 0.000 1129.520 4.000 ;
    END
  END c1_i_req_data[22]
  PIN c1_i_req_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1131.200 0.000 1131.760 4.000 ;
    END
  END c1_i_req_data[23]
  PIN c1_i_req_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1133.440 0.000 1134.000 4.000 ;
    END
  END c1_i_req_data[24]
  PIN c1_i_req_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1135.680 0.000 1136.240 4.000 ;
    END
  END c1_i_req_data[25]
  PIN c1_i_req_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1137.920 0.000 1138.480 4.000 ;
    END
  END c1_i_req_data[26]
  PIN c1_i_req_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1140.160 0.000 1140.720 4.000 ;
    END
  END c1_i_req_data[27]
  PIN c1_i_req_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1142.400 0.000 1142.960 4.000 ;
    END
  END c1_i_req_data[28]
  PIN c1_i_req_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1144.640 0.000 1145.200 4.000 ;
    END
  END c1_i_req_data[29]
  PIN c1_i_req_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 784.000 0.000 784.560 4.000 ;
    END
  END c1_i_req_data[2]
  PIN c1_i_req_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1146.880 0.000 1147.440 4.000 ;
    END
  END c1_i_req_data[30]
  PIN c1_i_req_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1149.120 0.000 1149.680 4.000 ;
    END
  END c1_i_req_data[31]
  PIN c1_i_req_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 810.880 0.000 811.440 4.000 ;
    END
  END c1_i_req_data[3]
  PIN c1_i_req_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 0.000 838.320 4.000 ;
    END
  END c1_i_req_data[4]
  PIN c1_i_req_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 864.640 0.000 865.200 4.000 ;
    END
  END c1_i_req_data[5]
  PIN c1_i_req_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 891.520 0.000 892.080 4.000 ;
    END
  END c1_i_req_data[6]
  PIN c1_i_req_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 918.400 0.000 918.960 4.000 ;
    END
  END c1_i_req_data[7]
  PIN c1_i_req_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 945.280 0.000 945.840 4.000 ;
    END
  END c1_i_req_data[8]
  PIN c1_i_req_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 967.680 0.000 968.240 4.000 ;
    END
  END c1_i_req_data[9]
  PIN c1_i_req_data_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 689.920 0.000 690.480 4.000 ;
    END
  END c1_i_req_data_valid
  PIN c1_o_c_data_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 0.000 692.720 4.000 ;
    END
  END c1_o_c_data_page
  PIN c1_o_c_instr_long
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 694.400 0.000 694.960 4.000 ;
    END
  END c1_o_c_instr_long
  PIN c1_o_c_instr_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 696.640 0.000 697.200 4.000 ;
    END
  END c1_o_c_instr_page
  PIN c1_o_icache_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 0.000 699.440 4.000 ;
    END
  END c1_o_icache_flush
  PIN c1_o_instr_long_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 728.000 0.000 728.560 4.000 ;
    END
  END c1_o_instr_long_addr[0]
  PIN c1_o_instr_long_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 757.120 0.000 757.680 4.000 ;
    END
  END c1_o_instr_long_addr[1]
  PIN c1_o_instr_long_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 0.000 786.800 4.000 ;
    END
  END c1_o_instr_long_addr[2]
  PIN c1_o_instr_long_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 0.000 813.680 4.000 ;
    END
  END c1_o_instr_long_addr[3]
  PIN c1_o_instr_long_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 0.000 840.560 4.000 ;
    END
  END c1_o_instr_long_addr[4]
  PIN c1_o_instr_long_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 0.000 867.440 4.000 ;
    END
  END c1_o_instr_long_addr[5]
  PIN c1_o_instr_long_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 0.000 894.320 4.000 ;
    END
  END c1_o_instr_long_addr[6]
  PIN c1_o_instr_long_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 0.000 921.200 4.000 ;
    END
  END c1_o_instr_long_addr[7]
  PIN c1_o_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 730.240 0.000 730.800 4.000 ;
    END
  END c1_o_mem_addr[0]
  PIN c1_o_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 992.320 0.000 992.880 4.000 ;
    END
  END c1_o_mem_addr[10]
  PIN c1_o_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 0.000 1015.280 4.000 ;
    END
  END c1_o_mem_addr[11]
  PIN c1_o_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1037.120 0.000 1037.680 4.000 ;
    END
  END c1_o_mem_addr[12]
  PIN c1_o_mem_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1059.520 0.000 1060.080 4.000 ;
    END
  END c1_o_mem_addr[13]
  PIN c1_o_mem_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1081.920 0.000 1082.480 4.000 ;
    END
  END c1_o_mem_addr[14]
  PIN c1_o_mem_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1104.320 0.000 1104.880 4.000 ;
    END
  END c1_o_mem_addr[15]
  PIN c1_o_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 0.000 759.920 4.000 ;
    END
  END c1_o_mem_addr[1]
  PIN c1_o_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 788.480 0.000 789.040 4.000 ;
    END
  END c1_o_mem_addr[2]
  PIN c1_o_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 815.360 0.000 815.920 4.000 ;
    END
  END c1_o_mem_addr[3]
  PIN c1_o_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 842.240 0.000 842.800 4.000 ;
    END
  END c1_o_mem_addr[4]
  PIN c1_o_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 869.120 0.000 869.680 4.000 ;
    END
  END c1_o_mem_addr[5]
  PIN c1_o_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 896.000 0.000 896.560 4.000 ;
    END
  END c1_o_mem_addr[6]
  PIN c1_o_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 922.880 0.000 923.440 4.000 ;
    END
  END c1_o_mem_addr[7]
  PIN c1_o_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 0.000 948.080 4.000 ;
    END
  END c1_o_mem_addr[8]
  PIN c1_o_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 969.920 0.000 970.480 4.000 ;
    END
  END c1_o_mem_addr[9]
  PIN c1_o_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 0.000 733.040 4.000 ;
    END
  END c1_o_mem_data[0]
  PIN c1_o_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 0.000 995.120 4.000 ;
    END
  END c1_o_mem_data[10]
  PIN c1_o_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1016.960 0.000 1017.520 4.000 ;
    END
  END c1_o_mem_data[11]
  PIN c1_o_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1039.360 0.000 1039.920 4.000 ;
    END
  END c1_o_mem_data[12]
  PIN c1_o_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1061.760 0.000 1062.320 4.000 ;
    END
  END c1_o_mem_data[13]
  PIN c1_o_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1084.160 0.000 1084.720 4.000 ;
    END
  END c1_o_mem_data[14]
  PIN c1_o_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1106.560 0.000 1107.120 4.000 ;
    END
  END c1_o_mem_data[15]
  PIN c1_o_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 761.600 0.000 762.160 4.000 ;
    END
  END c1_o_mem_data[1]
  PIN c1_o_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 790.720 0.000 791.280 4.000 ;
    END
  END c1_o_mem_data[2]
  PIN c1_o_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 817.600 0.000 818.160 4.000 ;
    END
  END c1_o_mem_data[3]
  PIN c1_o_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 844.480 0.000 845.040 4.000 ;
    END
  END c1_o_mem_data[4]
  PIN c1_o_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 871.360 0.000 871.920 4.000 ;
    END
  END c1_o_mem_data[5]
  PIN c1_o_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 898.240 0.000 898.800 4.000 ;
    END
  END c1_o_mem_data[6]
  PIN c1_o_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 925.120 0.000 925.680 4.000 ;
    END
  END c1_o_mem_data[7]
  PIN c1_o_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 949.760 0.000 950.320 4.000 ;
    END
  END c1_o_mem_data[8]
  PIN c1_o_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 972.160 0.000 972.720 4.000 ;
    END
  END c1_o_mem_data[9]
  PIN c1_o_mem_high_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 734.720 0.000 735.280 4.000 ;
    END
  END c1_o_mem_high_addr[0]
  PIN c1_o_mem_high_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 0.000 764.400 4.000 ;
    END
  END c1_o_mem_high_addr[1]
  PIN c1_o_mem_high_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 0.000 793.520 4.000 ;
    END
  END c1_o_mem_high_addr[2]
  PIN c1_o_mem_high_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 819.840 0.000 820.400 4.000 ;
    END
  END c1_o_mem_high_addr[3]
  PIN c1_o_mem_high_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 846.720 0.000 847.280 4.000 ;
    END
  END c1_o_mem_high_addr[4]
  PIN c1_o_mem_high_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 873.600 0.000 874.160 4.000 ;
    END
  END c1_o_mem_high_addr[5]
  PIN c1_o_mem_high_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 900.480 0.000 901.040 4.000 ;
    END
  END c1_o_mem_high_addr[6]
  PIN c1_o_mem_high_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 0.000 927.920 4.000 ;
    END
  END c1_o_mem_high_addr[7]
  PIN c1_o_mem_long_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 0.000 701.680 4.000 ;
    END
  END c1_o_mem_long_mode
  PIN c1_o_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 703.360 0.000 703.920 4.000 ;
    END
  END c1_o_mem_req
  PIN c1_o_mem_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 736.960 0.000 737.520 4.000 ;
    END
  END c1_o_mem_sel[0]
  PIN c1_o_mem_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 766.080 0.000 766.640 4.000 ;
    END
  END c1_o_mem_sel[1]
  PIN c1_o_mem_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 0.000 706.160 4.000 ;
    END
  END c1_o_mem_we
  PIN c1_o_req_active
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 707.840 0.000 708.400 4.000 ;
    END
  END c1_o_req_active
  PIN c1_o_req_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 0.000 739.760 4.000 ;
    END
  END c1_o_req_addr[0]
  PIN c1_o_req_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 996.800 0.000 997.360 4.000 ;
    END
  END c1_o_req_addr[10]
  PIN c1_o_req_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1019.200 0.000 1019.760 4.000 ;
    END
  END c1_o_req_addr[11]
  PIN c1_o_req_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1041.600 0.000 1042.160 4.000 ;
    END
  END c1_o_req_addr[12]
  PIN c1_o_req_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1064.000 0.000 1064.560 4.000 ;
    END
  END c1_o_req_addr[13]
  PIN c1_o_req_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1086.400 0.000 1086.960 4.000 ;
    END
  END c1_o_req_addr[14]
  PIN c1_o_req_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1108.800 0.000 1109.360 4.000 ;
    END
  END c1_o_req_addr[15]
  PIN c1_o_req_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 768.320 0.000 768.880 4.000 ;
    END
  END c1_o_req_addr[1]
  PIN c1_o_req_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 795.200 0.000 795.760 4.000 ;
    END
  END c1_o_req_addr[2]
  PIN c1_o_req_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 0.000 822.640 4.000 ;
    END
  END c1_o_req_addr[3]
  PIN c1_o_req_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 848.960 0.000 849.520 4.000 ;
    END
  END c1_o_req_addr[4]
  PIN c1_o_req_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 875.840 0.000 876.400 4.000 ;
    END
  END c1_o_req_addr[5]
  PIN c1_o_req_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 902.720 0.000 903.280 4.000 ;
    END
  END c1_o_req_addr[6]
  PIN c1_o_req_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 929.600 0.000 930.160 4.000 ;
    END
  END c1_o_req_addr[7]
  PIN c1_o_req_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 952.000 0.000 952.560 4.000 ;
    END
  END c1_o_req_addr[8]
  PIN c1_o_req_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 0.000 974.960 4.000 ;
    END
  END c1_o_req_addr[9]
  PIN c1_o_req_ppl_submit
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 710.080 0.000 710.640 4.000 ;
    END
  END c1_o_req_ppl_submit
  PIN c1_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 0.000 712.880 4.000 ;
    END
  END c1_rst
  PIN c1_sr_bus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 0.000 742.000 4.000 ;
    END
  END c1_sr_bus_addr[0]
  PIN c1_sr_bus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 999.040 0.000 999.600 4.000 ;
    END
  END c1_sr_bus_addr[10]
  PIN c1_sr_bus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1021.440 0.000 1022.000 4.000 ;
    END
  END c1_sr_bus_addr[11]
  PIN c1_sr_bus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1043.840 0.000 1044.400 4.000 ;
    END
  END c1_sr_bus_addr[12]
  PIN c1_sr_bus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1066.240 0.000 1066.800 4.000 ;
    END
  END c1_sr_bus_addr[13]
  PIN c1_sr_bus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1088.640 0.000 1089.200 4.000 ;
    END
  END c1_sr_bus_addr[14]
  PIN c1_sr_bus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1111.040 0.000 1111.600 4.000 ;
    END
  END c1_sr_bus_addr[15]
  PIN c1_sr_bus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 770.560 0.000 771.120 4.000 ;
    END
  END c1_sr_bus_addr[1]
  PIN c1_sr_bus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 797.440 0.000 798.000 4.000 ;
    END
  END c1_sr_bus_addr[2]
  PIN c1_sr_bus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 824.320 0.000 824.880 4.000 ;
    END
  END c1_sr_bus_addr[3]
  PIN c1_sr_bus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 851.200 0.000 851.760 4.000 ;
    END
  END c1_sr_bus_addr[4]
  PIN c1_sr_bus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 878.080 0.000 878.640 4.000 ;
    END
  END c1_sr_bus_addr[5]
  PIN c1_sr_bus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 904.960 0.000 905.520 4.000 ;
    END
  END c1_sr_bus_addr[6]
  PIN c1_sr_bus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 931.840 0.000 932.400 4.000 ;
    END
  END c1_sr_bus_addr[7]
  PIN c1_sr_bus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 0.000 954.800 4.000 ;
    END
  END c1_sr_bus_addr[8]
  PIN c1_sr_bus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 976.640 0.000 977.200 4.000 ;
    END
  END c1_sr_bus_addr[9]
  PIN c1_sr_bus_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 0.000 744.240 4.000 ;
    END
  END c1_sr_bus_data_o[0]
  PIN c1_sr_bus_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1001.280 0.000 1001.840 4.000 ;
    END
  END c1_sr_bus_data_o[10]
  PIN c1_sr_bus_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1023.680 0.000 1024.240 4.000 ;
    END
  END c1_sr_bus_data_o[11]
  PIN c1_sr_bus_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1046.080 0.000 1046.640 4.000 ;
    END
  END c1_sr_bus_data_o[12]
  PIN c1_sr_bus_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1068.480 0.000 1069.040 4.000 ;
    END
  END c1_sr_bus_data_o[13]
  PIN c1_sr_bus_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1090.880 0.000 1091.440 4.000 ;
    END
  END c1_sr_bus_data_o[14]
  PIN c1_sr_bus_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1113.280 0.000 1113.840 4.000 ;
    END
  END c1_sr_bus_data_o[15]
  PIN c1_sr_bus_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 0.000 773.360 4.000 ;
    END
  END c1_sr_bus_data_o[1]
  PIN c1_sr_bus_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 0.000 800.240 4.000 ;
    END
  END c1_sr_bus_data_o[2]
  PIN c1_sr_bus_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 0.000 827.120 4.000 ;
    END
  END c1_sr_bus_data_o[3]
  PIN c1_sr_bus_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 0.000 854.000 4.000 ;
    END
  END c1_sr_bus_data_o[4]
  PIN c1_sr_bus_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 0.000 880.880 4.000 ;
    END
  END c1_sr_bus_data_o[5]
  PIN c1_sr_bus_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 0.000 907.760 4.000 ;
    END
  END c1_sr_bus_data_o[6]
  PIN c1_sr_bus_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 0.000 934.640 4.000 ;
    END
  END c1_sr_bus_data_o[7]
  PIN c1_sr_bus_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 956.480 0.000 957.040 4.000 ;
    END
  END c1_sr_bus_data_o[8]
  PIN c1_sr_bus_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 978.880 0.000 979.440 4.000 ;
    END
  END c1_sr_bus_data_o[9]
  PIN c1_sr_bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 0.000 715.120 4.000 ;
    END
  END c1_sr_bus_we
  PIN core_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 521.920 0.000 522.480 4.000 ;
    END
  END core_clock
  PIN core_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 0.000 524.720 4.000 ;
    END
  END core_reset
  PIN dcache_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 346.000 30.800 350.000 ;
    END
  END dcache_mem_ack
  PIN dcache_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 346.000 138.320 350.000 ;
    END
  END dcache_mem_addr[0]
  PIN dcache_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 346.000 711.760 350.000 ;
    END
  END dcache_mem_addr[10]
  PIN dcache_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 764.960 346.000 765.520 350.000 ;
    END
  END dcache_mem_addr[11]
  PIN dcache_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 818.720 346.000 819.280 350.000 ;
    END
  END dcache_mem_addr[12]
  PIN dcache_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 346.000 873.040 350.000 ;
    END
  END dcache_mem_addr[13]
  PIN dcache_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 926.240 346.000 926.800 350.000 ;
    END
  END dcache_mem_addr[14]
  PIN dcache_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 980.000 346.000 980.560 350.000 ;
    END
  END dcache_mem_addr[15]
  PIN dcache_mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1033.760 346.000 1034.320 350.000 ;
    END
  END dcache_mem_addr[16]
  PIN dcache_mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1051.680 346.000 1052.240 350.000 ;
    END
  END dcache_mem_addr[17]
  PIN dcache_mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1069.600 346.000 1070.160 350.000 ;
    END
  END dcache_mem_addr[18]
  PIN dcache_mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1087.520 346.000 1088.080 350.000 ;
    END
  END dcache_mem_addr[19]
  PIN dcache_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 346.000 210.000 350.000 ;
    END
  END dcache_mem_addr[1]
  PIN dcache_mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 1105.440 346.000 1106.000 350.000 ;
    END
  END dcache_mem_addr[20]
  PIN dcache_mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1123.360 346.000 1123.920 350.000 ;
    END
  END dcache_mem_addr[21]
  PIN dcache_mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1141.280 346.000 1141.840 350.000 ;
    END
  END dcache_mem_addr[22]
  PIN dcache_mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1159.200 346.000 1159.760 350.000 ;
    END
  END dcache_mem_addr[23]
  PIN dcache_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 346.000 281.680 350.000 ;
    END
  END dcache_mem_addr[2]
  PIN dcache_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 346.000 335.440 350.000 ;
    END
  END dcache_mem_addr[3]
  PIN dcache_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 346.000 389.200 350.000 ;
    END
  END dcache_mem_addr[4]
  PIN dcache_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 442.400 346.000 442.960 350.000 ;
    END
  END dcache_mem_addr[5]
  PIN dcache_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 346.000 496.720 350.000 ;
    END
  END dcache_mem_addr[6]
  PIN dcache_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 346.000 550.480 350.000 ;
    END
  END dcache_mem_addr[7]
  PIN dcache_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 346.000 604.240 350.000 ;
    END
  END dcache_mem_addr[8]
  PIN dcache_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 657.440 346.000 658.000 350.000 ;
    END
  END dcache_mem_addr[9]
  PIN dcache_mem_cache_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 346.000 39.760 350.000 ;
    END
  END dcache_mem_cache_enable
  PIN dcache_mem_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 48.160 346.000 48.720 350.000 ;
    END
  END dcache_mem_exception
  PIN dcache_mem_i_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 346.000 147.280 350.000 ;
    END
  END dcache_mem_i_data[0]
  PIN dcache_mem_i_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 346.000 720.720 350.000 ;
    END
  END dcache_mem_i_data[10]
  PIN dcache_mem_i_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 773.920 346.000 774.480 350.000 ;
    END
  END dcache_mem_i_data[11]
  PIN dcache_mem_i_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 827.680 346.000 828.240 350.000 ;
    END
  END dcache_mem_i_data[12]
  PIN dcache_mem_i_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 881.440 346.000 882.000 350.000 ;
    END
  END dcache_mem_i_data[13]
  PIN dcache_mem_i_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 935.200 346.000 935.760 350.000 ;
    END
  END dcache_mem_i_data[14]
  PIN dcache_mem_i_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 988.960 346.000 989.520 350.000 ;
    END
  END dcache_mem_i_data[15]
  PIN dcache_mem_i_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 346.000 218.960 350.000 ;
    END
  END dcache_mem_i_data[1]
  PIN dcache_mem_i_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 290.080 346.000 290.640 350.000 ;
    END
  END dcache_mem_i_data[2]
  PIN dcache_mem_i_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 343.840 346.000 344.400 350.000 ;
    END
  END dcache_mem_i_data[3]
  PIN dcache_mem_i_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 346.000 398.160 350.000 ;
    END
  END dcache_mem_i_data[4]
  PIN dcache_mem_i_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 451.360 346.000 451.920 350.000 ;
    END
  END dcache_mem_i_data[5]
  PIN dcache_mem_i_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 346.000 505.680 350.000 ;
    END
  END dcache_mem_i_data[6]
  PIN dcache_mem_i_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 346.000 559.440 350.000 ;
    END
  END dcache_mem_i_data[7]
  PIN dcache_mem_i_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 612.640 346.000 613.200 350.000 ;
    END
  END dcache_mem_i_data[8]
  PIN dcache_mem_i_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 666.400 346.000 666.960 350.000 ;
    END
  END dcache_mem_i_data[9]
  PIN dcache_mem_o_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 346.000 156.240 350.000 ;
    END
  END dcache_mem_o_data[0]
  PIN dcache_mem_o_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 729.120 346.000 729.680 350.000 ;
    END
  END dcache_mem_o_data[10]
  PIN dcache_mem_o_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 346.000 783.440 350.000 ;
    END
  END dcache_mem_o_data[11]
  PIN dcache_mem_o_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 346.000 837.200 350.000 ;
    END
  END dcache_mem_o_data[12]
  PIN dcache_mem_o_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 890.400 346.000 890.960 350.000 ;
    END
  END dcache_mem_o_data[13]
  PIN dcache_mem_o_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 346.000 944.720 350.000 ;
    END
  END dcache_mem_o_data[14]
  PIN dcache_mem_o_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 997.920 346.000 998.480 350.000 ;
    END
  END dcache_mem_o_data[15]
  PIN dcache_mem_o_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 346.000 227.920 350.000 ;
    END
  END dcache_mem_o_data[1]
  PIN dcache_mem_o_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 346.000 299.600 350.000 ;
    END
  END dcache_mem_o_data[2]
  PIN dcache_mem_o_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 352.800 346.000 353.360 350.000 ;
    END
  END dcache_mem_o_data[3]
  PIN dcache_mem_o_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 346.000 407.120 350.000 ;
    END
  END dcache_mem_o_data[4]
  PIN dcache_mem_o_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 346.000 460.880 350.000 ;
    END
  END dcache_mem_o_data[5]
  PIN dcache_mem_o_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 514.080 346.000 514.640 350.000 ;
    END
  END dcache_mem_o_data[6]
  PIN dcache_mem_o_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 346.000 568.400 350.000 ;
    END
  END dcache_mem_o_data[7]
  PIN dcache_mem_o_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 621.600 346.000 622.160 350.000 ;
    END
  END dcache_mem_o_data[8]
  PIN dcache_mem_o_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 346.000 675.920 350.000 ;
    END
  END dcache_mem_o_data[9]
  PIN dcache_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 346.000 57.680 350.000 ;
    END
  END dcache_mem_req
  PIN dcache_mem_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 346.000 165.200 350.000 ;
    END
  END dcache_mem_sel[0]
  PIN dcache_mem_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 346.000 236.880 350.000 ;
    END
  END dcache_mem_sel[1]
  PIN dcache_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 346.000 66.640 350.000 ;
    END
  END dcache_mem_we
  PIN dcache_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 346.000 75.600 350.000 ;
    END
  END dcache_rst
  PIN dcache_wb_4_burst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 346.000 84.560 350.000 ;
    END
  END dcache_wb_4_burst
  PIN dcache_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 346.000 93.520 350.000 ;
    END
  END dcache_wb_ack
  PIN dcache_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 346.000 174.160 350.000 ;
    END
  END dcache_wb_adr[0]
  PIN dcache_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 738.080 346.000 738.640 350.000 ;
    END
  END dcache_wb_adr[10]
  PIN dcache_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 791.840 346.000 792.400 350.000 ;
    END
  END dcache_wb_adr[11]
  PIN dcache_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 845.600 346.000 846.160 350.000 ;
    END
  END dcache_wb_adr[12]
  PIN dcache_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 899.360 346.000 899.920 350.000 ;
    END
  END dcache_wb_adr[13]
  PIN dcache_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 953.120 346.000 953.680 350.000 ;
    END
  END dcache_wb_adr[14]
  PIN dcache_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1006.880 346.000 1007.440 350.000 ;
    END
  END dcache_wb_adr[15]
  PIN dcache_wb_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1042.720 346.000 1043.280 350.000 ;
    END
  END dcache_wb_adr[16]
  PIN dcache_wb_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1060.640 346.000 1061.200 350.000 ;
    END
  END dcache_wb_adr[17]
  PIN dcache_wb_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1078.560 346.000 1079.120 350.000 ;
    END
  END dcache_wb_adr[18]
  PIN dcache_wb_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1096.480 346.000 1097.040 350.000 ;
    END
  END dcache_wb_adr[19]
  PIN dcache_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 346.000 245.840 350.000 ;
    END
  END dcache_wb_adr[1]
  PIN dcache_wb_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1114.400 346.000 1114.960 350.000 ;
    END
  END dcache_wb_adr[20]
  PIN dcache_wb_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1132.320 346.000 1132.880 350.000 ;
    END
  END dcache_wb_adr[21]
  PIN dcache_wb_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1150.240 346.000 1150.800 350.000 ;
    END
  END dcache_wb_adr[22]
  PIN dcache_wb_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1168.160 346.000 1168.720 350.000 ;
    END
  END dcache_wb_adr[23]
  PIN dcache_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 346.000 308.560 350.000 ;
    END
  END dcache_wb_adr[2]
  PIN dcache_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 346.000 362.320 350.000 ;
    END
  END dcache_wb_adr[3]
  PIN dcache_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 346.000 416.080 350.000 ;
    END
  END dcache_wb_adr[4]
  PIN dcache_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 346.000 469.840 350.000 ;
    END
  END dcache_wb_adr[5]
  PIN dcache_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 523.040 346.000 523.600 350.000 ;
    END
  END dcache_wb_adr[6]
  PIN dcache_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 576.800 346.000 577.360 350.000 ;
    END
  END dcache_wb_adr[7]
  PIN dcache_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 346.000 631.120 350.000 ;
    END
  END dcache_wb_adr[8]
  PIN dcache_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 684.320 346.000 684.880 350.000 ;
    END
  END dcache_wb_adr[9]
  PIN dcache_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.920 346.000 102.480 350.000 ;
    END
  END dcache_wb_cyc
  PIN dcache_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 346.000 111.440 350.000 ;
    END
  END dcache_wb_err
  PIN dcache_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 346.000 183.120 350.000 ;
    END
  END dcache_wb_i_dat[0]
  PIN dcache_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 747.040 346.000 747.600 350.000 ;
    END
  END dcache_wb_i_dat[10]
  PIN dcache_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 800.800 346.000 801.360 350.000 ;
    END
  END dcache_wb_i_dat[11]
  PIN dcache_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 854.560 346.000 855.120 350.000 ;
    END
  END dcache_wb_i_dat[12]
  PIN dcache_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 908.320 346.000 908.880 350.000 ;
    END
  END dcache_wb_i_dat[13]
  PIN dcache_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 346.000 962.640 350.000 ;
    END
  END dcache_wb_i_dat[14]
  PIN dcache_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 1015.840 346.000 1016.400 350.000 ;
    END
  END dcache_wb_i_dat[15]
  PIN dcache_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 346.000 254.800 350.000 ;
    END
  END dcache_wb_i_dat[1]
  PIN dcache_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 346.000 317.520 350.000 ;
    END
  END dcache_wb_i_dat[2]
  PIN dcache_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 370.720 346.000 371.280 350.000 ;
    END
  END dcache_wb_i_dat[3]
  PIN dcache_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 424.480 346.000 425.040 350.000 ;
    END
  END dcache_wb_i_dat[4]
  PIN dcache_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 346.000 478.800 350.000 ;
    END
  END dcache_wb_i_dat[5]
  PIN dcache_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 346.000 532.560 350.000 ;
    END
  END dcache_wb_i_dat[6]
  PIN dcache_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 585.760 346.000 586.320 350.000 ;
    END
  END dcache_wb_i_dat[7]
  PIN dcache_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 346.000 640.080 350.000 ;
    END
  END dcache_wb_i_dat[8]
  PIN dcache_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 693.280 346.000 693.840 350.000 ;
    END
  END dcache_wb_i_dat[9]
  PIN dcache_wb_o_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 346.000 192.080 350.000 ;
    END
  END dcache_wb_o_dat[0]
  PIN dcache_wb_o_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 756.000 346.000 756.560 350.000 ;
    END
  END dcache_wb_o_dat[10]
  PIN dcache_wb_o_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 346.000 810.320 350.000 ;
    END
  END dcache_wb_o_dat[11]
  PIN dcache_wb_o_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 863.520 346.000 864.080 350.000 ;
    END
  END dcache_wb_o_dat[12]
  PIN dcache_wb_o_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 346.000 917.840 350.000 ;
    END
  END dcache_wb_o_dat[13]
  PIN dcache_wb_o_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 971.040 346.000 971.600 350.000 ;
    END
  END dcache_wb_o_dat[14]
  PIN dcache_wb_o_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1024.800 346.000 1025.360 350.000 ;
    END
  END dcache_wb_o_dat[15]
  PIN dcache_wb_o_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 346.000 263.760 350.000 ;
    END
  END dcache_wb_o_dat[1]
  PIN dcache_wb_o_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 346.000 326.480 350.000 ;
    END
  END dcache_wb_o_dat[2]
  PIN dcache_wb_o_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 379.680 346.000 380.240 350.000 ;
    END
  END dcache_wb_o_dat[3]
  PIN dcache_wb_o_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 346.000 434.000 350.000 ;
    END
  END dcache_wb_o_dat[4]
  PIN dcache_wb_o_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 487.200 346.000 487.760 350.000 ;
    END
  END dcache_wb_o_dat[5]
  PIN dcache_wb_o_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 346.000 541.520 350.000 ;
    END
  END dcache_wb_o_dat[6]
  PIN dcache_wb_o_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 594.720 346.000 595.280 350.000 ;
    END
  END dcache_wb_o_dat[7]
  PIN dcache_wb_o_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 346.000 649.040 350.000 ;
    END
  END dcache_wb_o_dat[8]
  PIN dcache_wb_o_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 346.000 702.800 350.000 ;
    END
  END dcache_wb_o_dat[9]
  PIN dcache_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 346.000 201.040 350.000 ;
    END
  END dcache_wb_sel[0]
  PIN dcache_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 346.000 272.720 350.000 ;
    END
  END dcache_wb_sel[1]
  PIN dcache_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 346.000 120.400 350.000 ;
    END
  END dcache_wb_stb
  PIN dcache_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 346.000 129.360 350.000 ;
    END
  END dcache_wb_we
  PIN ic0_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.280 4.000 21.840 ;
    END
  END ic0_mem_ack
  PIN ic0_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 54.880 4.000 55.440 ;
    END
  END ic0_mem_addr[0]
  PIN ic0_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.000 4.000 196.560 ;
    END
  END ic0_mem_addr[10]
  PIN ic0_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 209.440 4.000 210.000 ;
    END
  END ic0_mem_addr[11]
  PIN ic0_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 222.880 4.000 223.440 ;
    END
  END ic0_mem_addr[12]
  PIN ic0_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 236.320 4.000 236.880 ;
    END
  END ic0_mem_addr[13]
  PIN ic0_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.760 4.000 250.320 ;
    END
  END ic0_mem_addr[14]
  PIN ic0_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END ic0_mem_addr[15]
  PIN ic0_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 71.680 4.000 72.240 ;
    END
  END ic0_mem_addr[1]
  PIN ic0_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 4.000 89.040 ;
    END
  END ic0_mem_addr[2]
  PIN ic0_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 4.000 102.480 ;
    END
  END ic0_mem_addr[3]
  PIN ic0_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END ic0_mem_addr[4]
  PIN ic0_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 4.000 129.360 ;
    END
  END ic0_mem_addr[5]
  PIN ic0_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 4.000 142.800 ;
    END
  END ic0_mem_addr[6]
  PIN ic0_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 4.000 156.240 ;
    END
  END ic0_mem_addr[7]
  PIN ic0_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 4.000 169.680 ;
    END
  END ic0_mem_addr[8]
  PIN ic0_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 4.000 183.120 ;
    END
  END ic0_mem_addr[9]
  PIN ic0_mem_cache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 24.640 4.000 25.200 ;
    END
  END ic0_mem_cache_flush
  PIN ic0_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 58.240 4.000 58.800 ;
    END
  END ic0_mem_data[0]
  PIN ic0_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END ic0_mem_data[10]
  PIN ic0_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 212.800 4.000 213.360 ;
    END
  END ic0_mem_data[11]
  PIN ic0_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.240 4.000 226.800 ;
    END
  END ic0_mem_data[12]
  PIN ic0_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 239.680 4.000 240.240 ;
    END
  END ic0_mem_data[13]
  PIN ic0_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.120 4.000 253.680 ;
    END
  END ic0_mem_data[14]
  PIN ic0_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 4.000 267.120 ;
    END
  END ic0_mem_data[15]
  PIN ic0_mem_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 276.640 4.000 277.200 ;
    END
  END ic0_mem_data[16]
  PIN ic0_mem_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.000 4.000 280.560 ;
    END
  END ic0_mem_data[17]
  PIN ic0_mem_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 283.360 4.000 283.920 ;
    END
  END ic0_mem_data[18]
  PIN ic0_mem_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.720 4.000 287.280 ;
    END
  END ic0_mem_data[19]
  PIN ic0_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.040 4.000 75.600 ;
    END
  END ic0_mem_data[1]
  PIN ic0_mem_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.080 4.000 290.640 ;
    END
  END ic0_mem_data[20]
  PIN ic0_mem_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 293.440 4.000 294.000 ;
    END
  END ic0_mem_data[21]
  PIN ic0_mem_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 296.800 4.000 297.360 ;
    END
  END ic0_mem_data[22]
  PIN ic0_mem_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 300.160 4.000 300.720 ;
    END
  END ic0_mem_data[23]
  PIN ic0_mem_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 303.520 4.000 304.080 ;
    END
  END ic0_mem_data[24]
  PIN ic0_mem_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.880 4.000 307.440 ;
    END
  END ic0_mem_data[25]
  PIN ic0_mem_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.240 4.000 310.800 ;
    END
  END ic0_mem_data[26]
  PIN ic0_mem_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 313.600 4.000 314.160 ;
    END
  END ic0_mem_data[27]
  PIN ic0_mem_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 316.960 4.000 317.520 ;
    END
  END ic0_mem_data[28]
  PIN ic0_mem_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 320.320 4.000 320.880 ;
    END
  END ic0_mem_data[29]
  PIN ic0_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 91.840 4.000 92.400 ;
    END
  END ic0_mem_data[2]
  PIN ic0_mem_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 323.680 4.000 324.240 ;
    END
  END ic0_mem_data[30]
  PIN ic0_mem_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 327.040 4.000 327.600 ;
    END
  END ic0_mem_data[31]
  PIN ic0_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.280 4.000 105.840 ;
    END
  END ic0_mem_data[3]
  PIN ic0_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.720 4.000 119.280 ;
    END
  END ic0_mem_data[4]
  PIN ic0_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END ic0_mem_data[5]
  PIN ic0_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 145.600 4.000 146.160 ;
    END
  END ic0_mem_data[6]
  PIN ic0_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.040 4.000 159.600 ;
    END
  END ic0_mem_data[7]
  PIN ic0_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 172.480 4.000 173.040 ;
    END
  END ic0_mem_data[8]
  PIN ic0_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.920 4.000 186.480 ;
    END
  END ic0_mem_data[9]
  PIN ic0_mem_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.000 4.000 28.560 ;
    END
  END ic0_mem_ppl_submit
  PIN ic0_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.360 4.000 31.920 ;
    END
  END ic0_mem_req
  PIN ic0_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 4.000 35.280 ;
    END
  END ic0_rst
  PIN ic0_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.080 4.000 38.640 ;
    END
  END ic0_wb_ack
  PIN ic0_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 4.000 62.160 ;
    END
  END ic0_wb_adr[0]
  PIN ic0_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 202.720 4.000 203.280 ;
    END
  END ic0_wb_adr[10]
  PIN ic0_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 4.000 216.720 ;
    END
  END ic0_wb_adr[11]
  PIN ic0_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 229.600 4.000 230.160 ;
    END
  END ic0_wb_adr[12]
  PIN ic0_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.040 4.000 243.600 ;
    END
  END ic0_wb_adr[13]
  PIN ic0_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 256.480 4.000 257.040 ;
    END
  END ic0_wb_adr[14]
  PIN ic0_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.920 4.000 270.480 ;
    END
  END ic0_wb_adr[15]
  PIN ic0_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END ic0_wb_adr[1]
  PIN ic0_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.200 4.000 95.760 ;
    END
  END ic0_wb_adr[2]
  PIN ic0_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 108.640 4.000 109.200 ;
    END
  END ic0_wb_adr[3]
  PIN ic0_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.080 4.000 122.640 ;
    END
  END ic0_wb_adr[4]
  PIN ic0_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 135.520 4.000 136.080 ;
    END
  END ic0_wb_adr[5]
  PIN ic0_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 4.000 149.520 ;
    END
  END ic0_wb_adr[6]
  PIN ic0_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 4.000 162.960 ;
    END
  END ic0_wb_adr[7]
  PIN ic0_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 175.840 4.000 176.400 ;
    END
  END ic0_wb_adr[8]
  PIN ic0_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END ic0_wb_adr[9]
  PIN ic0_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 4.000 42.000 ;
    END
  END ic0_wb_cyc
  PIN ic0_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 44.800 4.000 45.360 ;
    END
  END ic0_wb_err
  PIN ic0_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 4.000 65.520 ;
    END
  END ic0_wb_i_dat[0]
  PIN ic0_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.080 4.000 206.640 ;
    END
  END ic0_wb_i_dat[10]
  PIN ic0_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 219.520 4.000 220.080 ;
    END
  END ic0_wb_i_dat[11]
  PIN ic0_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.960 4.000 233.520 ;
    END
  END ic0_wb_i_dat[12]
  PIN ic0_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.400 4.000 246.960 ;
    END
  END ic0_wb_i_dat[13]
  PIN ic0_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 259.840 4.000 260.400 ;
    END
  END ic0_wb_i_dat[14]
  PIN ic0_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 273.280 4.000 273.840 ;
    END
  END ic0_wb_i_dat[15]
  PIN ic0_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 4.000 82.320 ;
    END
  END ic0_wb_i_dat[1]
  PIN ic0_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 98.560 4.000 99.120 ;
    END
  END ic0_wb_i_dat[2]
  PIN ic0_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.000 4.000 112.560 ;
    END
  END ic0_wb_i_dat[3]
  PIN ic0_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 125.440 4.000 126.000 ;
    END
  END ic0_wb_i_dat[4]
  PIN ic0_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 138.880 4.000 139.440 ;
    END
  END ic0_wb_i_dat[5]
  PIN ic0_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END ic0_wb_i_dat[6]
  PIN ic0_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 165.760 4.000 166.320 ;
    END
  END ic0_wb_i_dat[7]
  PIN ic0_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.200 4.000 179.760 ;
    END
  END ic0_wb_i_dat[8]
  PIN ic0_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 192.640 4.000 193.200 ;
    END
  END ic0_wb_i_dat[9]
  PIN ic0_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.320 4.000 68.880 ;
    END
  END ic0_wb_sel[0]
  PIN ic0_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.120 4.000 85.680 ;
    END
  END ic0_wb_sel[1]
  PIN ic0_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 4.000 48.720 ;
    END
  END ic0_wb_stb
  PIN ic0_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 51.520 4.000 52.080 ;
    END
  END ic0_wb_we
  PIN ic1_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 21.280 1200.000 21.840 ;
    END
  END ic1_mem_ack
  PIN ic1_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 54.880 1200.000 55.440 ;
    END
  END ic1_mem_addr[0]
  PIN ic1_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 196.000 1200.000 196.560 ;
    END
  END ic1_mem_addr[10]
  PIN ic1_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 209.440 1200.000 210.000 ;
    END
  END ic1_mem_addr[11]
  PIN ic1_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 222.880 1200.000 223.440 ;
    END
  END ic1_mem_addr[12]
  PIN ic1_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 236.320 1200.000 236.880 ;
    END
  END ic1_mem_addr[13]
  PIN ic1_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 249.760 1200.000 250.320 ;
    END
  END ic1_mem_addr[14]
  PIN ic1_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 263.200 1200.000 263.760 ;
    END
  END ic1_mem_addr[15]
  PIN ic1_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 71.680 1200.000 72.240 ;
    END
  END ic1_mem_addr[1]
  PIN ic1_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 88.480 1200.000 89.040 ;
    END
  END ic1_mem_addr[2]
  PIN ic1_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 101.920 1200.000 102.480 ;
    END
  END ic1_mem_addr[3]
  PIN ic1_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 115.360 1200.000 115.920 ;
    END
  END ic1_mem_addr[4]
  PIN ic1_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 128.800 1200.000 129.360 ;
    END
  END ic1_mem_addr[5]
  PIN ic1_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 142.240 1200.000 142.800 ;
    END
  END ic1_mem_addr[6]
  PIN ic1_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 155.680 1200.000 156.240 ;
    END
  END ic1_mem_addr[7]
  PIN ic1_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 169.120 1200.000 169.680 ;
    END
  END ic1_mem_addr[8]
  PIN ic1_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 182.560 1200.000 183.120 ;
    END
  END ic1_mem_addr[9]
  PIN ic1_mem_cache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 24.640 1200.000 25.200 ;
    END
  END ic1_mem_cache_flush
  PIN ic1_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 58.240 1200.000 58.800 ;
    END
  END ic1_mem_data[0]
  PIN ic1_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 199.360 1200.000 199.920 ;
    END
  END ic1_mem_data[10]
  PIN ic1_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 212.800 1200.000 213.360 ;
    END
  END ic1_mem_data[11]
  PIN ic1_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 226.240 1200.000 226.800 ;
    END
  END ic1_mem_data[12]
  PIN ic1_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 239.680 1200.000 240.240 ;
    END
  END ic1_mem_data[13]
  PIN ic1_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 253.120 1200.000 253.680 ;
    END
  END ic1_mem_data[14]
  PIN ic1_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 266.560 1200.000 267.120 ;
    END
  END ic1_mem_data[15]
  PIN ic1_mem_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 276.640 1200.000 277.200 ;
    END
  END ic1_mem_data[16]
  PIN ic1_mem_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 280.000 1200.000 280.560 ;
    END
  END ic1_mem_data[17]
  PIN ic1_mem_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 283.360 1200.000 283.920 ;
    END
  END ic1_mem_data[18]
  PIN ic1_mem_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 286.720 1200.000 287.280 ;
    END
  END ic1_mem_data[19]
  PIN ic1_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 75.040 1200.000 75.600 ;
    END
  END ic1_mem_data[1]
  PIN ic1_mem_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 290.080 1200.000 290.640 ;
    END
  END ic1_mem_data[20]
  PIN ic1_mem_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 293.440 1200.000 294.000 ;
    END
  END ic1_mem_data[21]
  PIN ic1_mem_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 296.800 1200.000 297.360 ;
    END
  END ic1_mem_data[22]
  PIN ic1_mem_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 300.160 1200.000 300.720 ;
    END
  END ic1_mem_data[23]
  PIN ic1_mem_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 303.520 1200.000 304.080 ;
    END
  END ic1_mem_data[24]
  PIN ic1_mem_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 306.880 1200.000 307.440 ;
    END
  END ic1_mem_data[25]
  PIN ic1_mem_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 310.240 1200.000 310.800 ;
    END
  END ic1_mem_data[26]
  PIN ic1_mem_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 313.600 1200.000 314.160 ;
    END
  END ic1_mem_data[27]
  PIN ic1_mem_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 316.960 1200.000 317.520 ;
    END
  END ic1_mem_data[28]
  PIN ic1_mem_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 320.320 1200.000 320.880 ;
    END
  END ic1_mem_data[29]
  PIN ic1_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 91.840 1200.000 92.400 ;
    END
  END ic1_mem_data[2]
  PIN ic1_mem_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 323.680 1200.000 324.240 ;
    END
  END ic1_mem_data[30]
  PIN ic1_mem_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 327.040 1200.000 327.600 ;
    END
  END ic1_mem_data[31]
  PIN ic1_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 105.280 1200.000 105.840 ;
    END
  END ic1_mem_data[3]
  PIN ic1_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 118.720 1200.000 119.280 ;
    END
  END ic1_mem_data[4]
  PIN ic1_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 132.160 1200.000 132.720 ;
    END
  END ic1_mem_data[5]
  PIN ic1_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 145.600 1200.000 146.160 ;
    END
  END ic1_mem_data[6]
  PIN ic1_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 159.040 1200.000 159.600 ;
    END
  END ic1_mem_data[7]
  PIN ic1_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 172.480 1200.000 173.040 ;
    END
  END ic1_mem_data[8]
  PIN ic1_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 185.920 1200.000 186.480 ;
    END
  END ic1_mem_data[9]
  PIN ic1_mem_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 28.000 1200.000 28.560 ;
    END
  END ic1_mem_ppl_submit
  PIN ic1_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 31.360 1200.000 31.920 ;
    END
  END ic1_mem_req
  PIN ic1_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 34.720 1200.000 35.280 ;
    END
  END ic1_rst
  PIN ic1_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 38.080 1200.000 38.640 ;
    END
  END ic1_wb_ack
  PIN ic1_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 61.600 1200.000 62.160 ;
    END
  END ic1_wb_adr[0]
  PIN ic1_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 202.720 1200.000 203.280 ;
    END
  END ic1_wb_adr[10]
  PIN ic1_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 216.160 1200.000 216.720 ;
    END
  END ic1_wb_adr[11]
  PIN ic1_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 229.600 1200.000 230.160 ;
    END
  END ic1_wb_adr[12]
  PIN ic1_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 243.040 1200.000 243.600 ;
    END
  END ic1_wb_adr[13]
  PIN ic1_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 256.480 1200.000 257.040 ;
    END
  END ic1_wb_adr[14]
  PIN ic1_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 269.920 1200.000 270.480 ;
    END
  END ic1_wb_adr[15]
  PIN ic1_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 78.400 1200.000 78.960 ;
    END
  END ic1_wb_adr[1]
  PIN ic1_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 95.200 1200.000 95.760 ;
    END
  END ic1_wb_adr[2]
  PIN ic1_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 108.640 1200.000 109.200 ;
    END
  END ic1_wb_adr[3]
  PIN ic1_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 122.080 1200.000 122.640 ;
    END
  END ic1_wb_adr[4]
  PIN ic1_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 135.520 1200.000 136.080 ;
    END
  END ic1_wb_adr[5]
  PIN ic1_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 148.960 1200.000 149.520 ;
    END
  END ic1_wb_adr[6]
  PIN ic1_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 162.400 1200.000 162.960 ;
    END
  END ic1_wb_adr[7]
  PIN ic1_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 175.840 1200.000 176.400 ;
    END
  END ic1_wb_adr[8]
  PIN ic1_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 189.280 1200.000 189.840 ;
    END
  END ic1_wb_adr[9]
  PIN ic1_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 41.440 1200.000 42.000 ;
    END
  END ic1_wb_cyc
  PIN ic1_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 44.800 1200.000 45.360 ;
    END
  END ic1_wb_err
  PIN ic1_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 64.960 1200.000 65.520 ;
    END
  END ic1_wb_i_dat[0]
  PIN ic1_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 206.080 1200.000 206.640 ;
    END
  END ic1_wb_i_dat[10]
  PIN ic1_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 219.520 1200.000 220.080 ;
    END
  END ic1_wb_i_dat[11]
  PIN ic1_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 232.960 1200.000 233.520 ;
    END
  END ic1_wb_i_dat[12]
  PIN ic1_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 246.400 1200.000 246.960 ;
    END
  END ic1_wb_i_dat[13]
  PIN ic1_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 259.840 1200.000 260.400 ;
    END
  END ic1_wb_i_dat[14]
  PIN ic1_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 273.280 1200.000 273.840 ;
    END
  END ic1_wb_i_dat[15]
  PIN ic1_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 81.760 1200.000 82.320 ;
    END
  END ic1_wb_i_dat[1]
  PIN ic1_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 98.560 1200.000 99.120 ;
    END
  END ic1_wb_i_dat[2]
  PIN ic1_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 112.000 1200.000 112.560 ;
    END
  END ic1_wb_i_dat[3]
  PIN ic1_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 125.440 1200.000 126.000 ;
    END
  END ic1_wb_i_dat[4]
  PIN ic1_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 138.880 1200.000 139.440 ;
    END
  END ic1_wb_i_dat[5]
  PIN ic1_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 152.320 1200.000 152.880 ;
    END
  END ic1_wb_i_dat[6]
  PIN ic1_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 165.760 1200.000 166.320 ;
    END
  END ic1_wb_i_dat[7]
  PIN ic1_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 179.200 1200.000 179.760 ;
    END
  END ic1_wb_i_dat[8]
  PIN ic1_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 192.640 1200.000 193.200 ;
    END
  END ic1_wb_i_dat[9]
  PIN ic1_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 68.320 1200.000 68.880 ;
    END
  END ic1_wb_sel[0]
  PIN ic1_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 85.120 1200.000 85.680 ;
    END
  END ic1_wb_sel[1]
  PIN ic1_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 48.160 1200.000 48.720 ;
    END
  END ic1_wb_stb
  PIN ic1_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1196.000 51.520 1200.000 52.080 ;
    END
  END ic1_wb_we
  PIN inner_disable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 0.000 526.960 4.000 ;
    END
  END inner_disable
  PIN inner_embed_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 0.000 529.200 4.000 ;
    END
  END inner_embed_mode
  PIN inner_ext_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 0.000 531.440 4.000 ;
    END
  END inner_ext_irq
  PIN inner_wb_4_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 533.120 0.000 533.680 4.000 ;
    END
  END inner_wb_4_burst
  PIN inner_wb_8_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 535.360 0.000 535.920 4.000 ;
    END
  END inner_wb_8_burst
  PIN inner_wb_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 0.000 538.160 4.000 ;
    END
  END inner_wb_ack
  PIN inner_wb_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 0.000 549.360 4.000 ;
    END
  END inner_wb_adr[0]
  PIN inner_wb_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 0.000 621.040 4.000 ;
    END
  END inner_wb_adr[10]
  PIN inner_wb_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 627.200 0.000 627.760 4.000 ;
    END
  END inner_wb_adr[11]
  PIN inner_wb_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 0.000 634.480 4.000 ;
    END
  END inner_wb_adr[12]
  PIN inner_wb_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 640.640 0.000 641.200 4.000 ;
    END
  END inner_wb_adr[13]
  PIN inner_wb_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 0.000 647.920 4.000 ;
    END
  END inner_wb_adr[14]
  PIN inner_wb_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 654.080 0.000 654.640 4.000 ;
    END
  END inner_wb_adr[15]
  PIN inner_wb_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 0.000 661.360 4.000 ;
    END
  END inner_wb_adr[16]
  PIN inner_wb_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 663.040 0.000 663.600 4.000 ;
    END
  END inner_wb_adr[17]
  PIN inner_wb_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 0.000 665.840 4.000 ;
    END
  END inner_wb_adr[18]
  PIN inner_wb_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 667.520 0.000 668.080 4.000 ;
    END
  END inner_wb_adr[19]
  PIN inner_wb_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 0.000 558.320 4.000 ;
    END
  END inner_wb_adr[1]
  PIN inner_wb_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 669.760 0.000 670.320 4.000 ;
    END
  END inner_wb_adr[20]
  PIN inner_wb_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 0.000 672.560 4.000 ;
    END
  END inner_wb_adr[21]
  PIN inner_wb_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 674.240 0.000 674.800 4.000 ;
    END
  END inner_wb_adr[22]
  PIN inner_wb_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 676.480 0.000 677.040 4.000 ;
    END
  END inner_wb_adr[23]
  PIN inner_wb_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 0.000 567.280 4.000 ;
    END
  END inner_wb_adr[2]
  PIN inner_wb_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 573.440 0.000 574.000 4.000 ;
    END
  END inner_wb_adr[3]
  PIN inner_wb_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 0.000 580.720 4.000 ;
    END
  END inner_wb_adr[4]
  PIN inner_wb_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 586.880 0.000 587.440 4.000 ;
    END
  END inner_wb_adr[5]
  PIN inner_wb_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 0.000 594.160 4.000 ;
    END
  END inner_wb_adr[6]
  PIN inner_wb_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 600.320 0.000 600.880 4.000 ;
    END
  END inner_wb_adr[7]
  PIN inner_wb_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 0.000 607.600 4.000 ;
    END
  END inner_wb_adr[8]
  PIN inner_wb_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 613.760 0.000 614.320 4.000 ;
    END
  END inner_wb_adr[9]
  PIN inner_wb_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END inner_wb_cyc
  PIN inner_wb_err
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 542.080 0.000 542.640 4.000 ;
    END
  END inner_wb_err
  PIN inner_wb_i_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 0.000 551.600 4.000 ;
    END
  END inner_wb_i_dat[0]
  PIN inner_wb_i_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 0.000 623.280 4.000 ;
    END
  END inner_wb_i_dat[10]
  PIN inner_wb_i_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 629.440 0.000 630.000 4.000 ;
    END
  END inner_wb_i_dat[11]
  PIN inner_wb_i_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 636.160 0.000 636.720 4.000 ;
    END
  END inner_wb_i_dat[12]
  PIN inner_wb_i_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 642.880 0.000 643.440 4.000 ;
    END
  END inner_wb_i_dat[13]
  PIN inner_wb_i_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 0.000 650.160 4.000 ;
    END
  END inner_wb_i_dat[14]
  PIN inner_wb_i_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 656.320 0.000 656.880 4.000 ;
    END
  END inner_wb_i_dat[15]
  PIN inner_wb_i_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 0.000 560.560 4.000 ;
    END
  END inner_wb_i_dat[1]
  PIN inner_wb_i_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 568.960 0.000 569.520 4.000 ;
    END
  END inner_wb_i_dat[2]
  PIN inner_wb_i_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END inner_wb_i_dat[3]
  PIN inner_wb_i_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 582.400 0.000 582.960 4.000 ;
    END
  END inner_wb_i_dat[4]
  PIN inner_wb_i_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 589.120 0.000 589.680 4.000 ;
    END
  END inner_wb_i_dat[5]
  PIN inner_wb_i_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 595.840 0.000 596.400 4.000 ;
    END
  END inner_wb_i_dat[6]
  PIN inner_wb_i_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 602.560 0.000 603.120 4.000 ;
    END
  END inner_wb_i_dat[7]
  PIN inner_wb_i_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 609.280 0.000 609.840 4.000 ;
    END
  END inner_wb_i_dat[8]
  PIN inner_wb_i_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 0.000 616.560 4.000 ;
    END
  END inner_wb_i_dat[9]
  PIN inner_wb_o_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 0.000 553.840 4.000 ;
    END
  END inner_wb_o_dat[0]
  PIN inner_wb_o_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 0.000 625.520 4.000 ;
    END
  END inner_wb_o_dat[10]
  PIN inner_wb_o_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 0.000 632.240 4.000 ;
    END
  END inner_wb_o_dat[11]
  PIN inner_wb_o_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 0.000 638.960 4.000 ;
    END
  END inner_wb_o_dat[12]
  PIN inner_wb_o_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 0.000 645.680 4.000 ;
    END
  END inner_wb_o_dat[13]
  PIN inner_wb_o_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 0.000 652.400 4.000 ;
    END
  END inner_wb_o_dat[14]
  PIN inner_wb_o_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 0.000 659.120 4.000 ;
    END
  END inner_wb_o_dat[15]
  PIN inner_wb_o_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 562.240 0.000 562.800 4.000 ;
    END
  END inner_wb_o_dat[1]
  PIN inner_wb_o_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 0.000 571.760 4.000 ;
    END
  END inner_wb_o_dat[2]
  PIN inner_wb_o_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 0.000 578.480 4.000 ;
    END
  END inner_wb_o_dat[3]
  PIN inner_wb_o_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 0.000 585.200 4.000 ;
    END
  END inner_wb_o_dat[4]
  PIN inner_wb_o_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 0.000 591.920 4.000 ;
    END
  END inner_wb_o_dat[5]
  PIN inner_wb_o_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 0.000 598.640 4.000 ;
    END
  END inner_wb_o_dat[6]
  PIN inner_wb_o_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 0.000 605.360 4.000 ;
    END
  END inner_wb_o_dat[7]
  PIN inner_wb_o_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 0.000 612.080 4.000 ;
    END
  END inner_wb_o_dat[8]
  PIN inner_wb_o_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 0.000 618.800 4.000 ;
    END
  END inner_wb_o_dat[9]
  PIN inner_wb_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 0.000 556.080 4.000 ;
    END
  END inner_wb_sel[0]
  PIN inner_wb_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 0.000 565.040 4.000 ;
    END
  END inner_wb_sel[1]
  PIN inner_wb_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 0.000 544.880 4.000 ;
    END
  END inner_wb_stb
  PIN inner_wb_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 0.000 547.120 4.000 ;
    END
  END inner_wb_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 333.500 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 333.500 ;
    END
  END vssd1
  OBS
      LAYER Metal1 ;
        RECT 6.720 9.110 1192.800 335.850 ;
      LAYER Metal2 ;
        RECT 6.300 345.700 29.940 346.500 ;
        RECT 31.100 345.700 38.900 346.500 ;
        RECT 40.060 345.700 47.860 346.500 ;
        RECT 49.020 345.700 56.820 346.500 ;
        RECT 57.980 345.700 65.780 346.500 ;
        RECT 66.940 345.700 74.740 346.500 ;
        RECT 75.900 345.700 83.700 346.500 ;
        RECT 84.860 345.700 92.660 346.500 ;
        RECT 93.820 345.700 101.620 346.500 ;
        RECT 102.780 345.700 110.580 346.500 ;
        RECT 111.740 345.700 119.540 346.500 ;
        RECT 120.700 345.700 128.500 346.500 ;
        RECT 129.660 345.700 137.460 346.500 ;
        RECT 138.620 345.700 146.420 346.500 ;
        RECT 147.580 345.700 155.380 346.500 ;
        RECT 156.540 345.700 164.340 346.500 ;
        RECT 165.500 345.700 173.300 346.500 ;
        RECT 174.460 345.700 182.260 346.500 ;
        RECT 183.420 345.700 191.220 346.500 ;
        RECT 192.380 345.700 200.180 346.500 ;
        RECT 201.340 345.700 209.140 346.500 ;
        RECT 210.300 345.700 218.100 346.500 ;
        RECT 219.260 345.700 227.060 346.500 ;
        RECT 228.220 345.700 236.020 346.500 ;
        RECT 237.180 345.700 244.980 346.500 ;
        RECT 246.140 345.700 253.940 346.500 ;
        RECT 255.100 345.700 262.900 346.500 ;
        RECT 264.060 345.700 271.860 346.500 ;
        RECT 273.020 345.700 280.820 346.500 ;
        RECT 281.980 345.700 289.780 346.500 ;
        RECT 290.940 345.700 298.740 346.500 ;
        RECT 299.900 345.700 307.700 346.500 ;
        RECT 308.860 345.700 316.660 346.500 ;
        RECT 317.820 345.700 325.620 346.500 ;
        RECT 326.780 345.700 334.580 346.500 ;
        RECT 335.740 345.700 343.540 346.500 ;
        RECT 344.700 345.700 352.500 346.500 ;
        RECT 353.660 345.700 361.460 346.500 ;
        RECT 362.620 345.700 370.420 346.500 ;
        RECT 371.580 345.700 379.380 346.500 ;
        RECT 380.540 345.700 388.340 346.500 ;
        RECT 389.500 345.700 397.300 346.500 ;
        RECT 398.460 345.700 406.260 346.500 ;
        RECT 407.420 345.700 415.220 346.500 ;
        RECT 416.380 345.700 424.180 346.500 ;
        RECT 425.340 345.700 433.140 346.500 ;
        RECT 434.300 345.700 442.100 346.500 ;
        RECT 443.260 345.700 451.060 346.500 ;
        RECT 452.220 345.700 460.020 346.500 ;
        RECT 461.180 345.700 468.980 346.500 ;
        RECT 470.140 345.700 477.940 346.500 ;
        RECT 479.100 345.700 486.900 346.500 ;
        RECT 488.060 345.700 495.860 346.500 ;
        RECT 497.020 345.700 504.820 346.500 ;
        RECT 505.980 345.700 513.780 346.500 ;
        RECT 514.940 345.700 522.740 346.500 ;
        RECT 523.900 345.700 531.700 346.500 ;
        RECT 532.860 345.700 540.660 346.500 ;
        RECT 541.820 345.700 549.620 346.500 ;
        RECT 550.780 345.700 558.580 346.500 ;
        RECT 559.740 345.700 567.540 346.500 ;
        RECT 568.700 345.700 576.500 346.500 ;
        RECT 577.660 345.700 585.460 346.500 ;
        RECT 586.620 345.700 594.420 346.500 ;
        RECT 595.580 345.700 603.380 346.500 ;
        RECT 604.540 345.700 612.340 346.500 ;
        RECT 613.500 345.700 621.300 346.500 ;
        RECT 622.460 345.700 630.260 346.500 ;
        RECT 631.420 345.700 639.220 346.500 ;
        RECT 640.380 345.700 648.180 346.500 ;
        RECT 649.340 345.700 657.140 346.500 ;
        RECT 658.300 345.700 666.100 346.500 ;
        RECT 667.260 345.700 675.060 346.500 ;
        RECT 676.220 345.700 684.020 346.500 ;
        RECT 685.180 345.700 692.980 346.500 ;
        RECT 694.140 345.700 701.940 346.500 ;
        RECT 703.100 345.700 710.900 346.500 ;
        RECT 712.060 345.700 719.860 346.500 ;
        RECT 721.020 345.700 728.820 346.500 ;
        RECT 729.980 345.700 737.780 346.500 ;
        RECT 738.940 345.700 746.740 346.500 ;
        RECT 747.900 345.700 755.700 346.500 ;
        RECT 756.860 345.700 764.660 346.500 ;
        RECT 765.820 345.700 773.620 346.500 ;
        RECT 774.780 345.700 782.580 346.500 ;
        RECT 783.740 345.700 791.540 346.500 ;
        RECT 792.700 345.700 800.500 346.500 ;
        RECT 801.660 345.700 809.460 346.500 ;
        RECT 810.620 345.700 818.420 346.500 ;
        RECT 819.580 345.700 827.380 346.500 ;
        RECT 828.540 345.700 836.340 346.500 ;
        RECT 837.500 345.700 845.300 346.500 ;
        RECT 846.460 345.700 854.260 346.500 ;
        RECT 855.420 345.700 863.220 346.500 ;
        RECT 864.380 345.700 872.180 346.500 ;
        RECT 873.340 345.700 881.140 346.500 ;
        RECT 882.300 345.700 890.100 346.500 ;
        RECT 891.260 345.700 899.060 346.500 ;
        RECT 900.220 345.700 908.020 346.500 ;
        RECT 909.180 345.700 916.980 346.500 ;
        RECT 918.140 345.700 925.940 346.500 ;
        RECT 927.100 345.700 934.900 346.500 ;
        RECT 936.060 345.700 943.860 346.500 ;
        RECT 945.020 345.700 952.820 346.500 ;
        RECT 953.980 345.700 961.780 346.500 ;
        RECT 962.940 345.700 970.740 346.500 ;
        RECT 971.900 345.700 979.700 346.500 ;
        RECT 980.860 345.700 988.660 346.500 ;
        RECT 989.820 345.700 997.620 346.500 ;
        RECT 998.780 345.700 1006.580 346.500 ;
        RECT 1007.740 345.700 1015.540 346.500 ;
        RECT 1016.700 345.700 1024.500 346.500 ;
        RECT 1025.660 345.700 1033.460 346.500 ;
        RECT 1034.620 345.700 1042.420 346.500 ;
        RECT 1043.580 345.700 1051.380 346.500 ;
        RECT 1052.540 345.700 1060.340 346.500 ;
        RECT 1061.500 345.700 1069.300 346.500 ;
        RECT 1070.460 345.700 1078.260 346.500 ;
        RECT 1079.420 345.700 1087.220 346.500 ;
        RECT 1088.380 345.700 1096.180 346.500 ;
        RECT 1097.340 345.700 1105.140 346.500 ;
        RECT 1106.300 345.700 1114.100 346.500 ;
        RECT 1115.260 345.700 1123.060 346.500 ;
        RECT 1124.220 345.700 1132.020 346.500 ;
        RECT 1133.180 345.700 1140.980 346.500 ;
        RECT 1142.140 345.700 1149.940 346.500 ;
        RECT 1151.100 345.700 1158.900 346.500 ;
        RECT 1160.060 345.700 1167.860 346.500 ;
        RECT 1169.020 345.700 1193.220 346.500 ;
        RECT 6.300 4.300 1193.220 345.700 ;
        RECT 6.300 1.770 48.980 4.300 ;
        RECT 50.140 1.770 51.220 4.300 ;
        RECT 52.380 1.770 53.460 4.300 ;
        RECT 54.620 1.770 55.700 4.300 ;
        RECT 56.860 1.770 57.940 4.300 ;
        RECT 59.100 1.770 60.180 4.300 ;
        RECT 61.340 1.770 62.420 4.300 ;
        RECT 63.580 1.770 64.660 4.300 ;
        RECT 65.820 1.770 66.900 4.300 ;
        RECT 68.060 1.770 69.140 4.300 ;
        RECT 70.300 1.770 71.380 4.300 ;
        RECT 72.540 1.770 73.620 4.300 ;
        RECT 74.780 1.770 75.860 4.300 ;
        RECT 77.020 1.770 78.100 4.300 ;
        RECT 79.260 1.770 80.340 4.300 ;
        RECT 81.500 1.770 82.580 4.300 ;
        RECT 83.740 1.770 84.820 4.300 ;
        RECT 85.980 1.770 87.060 4.300 ;
        RECT 88.220 1.770 89.300 4.300 ;
        RECT 90.460 1.770 91.540 4.300 ;
        RECT 92.700 1.770 93.780 4.300 ;
        RECT 94.940 1.770 96.020 4.300 ;
        RECT 97.180 1.770 98.260 4.300 ;
        RECT 99.420 1.770 100.500 4.300 ;
        RECT 101.660 1.770 102.740 4.300 ;
        RECT 103.900 1.770 104.980 4.300 ;
        RECT 106.140 1.770 107.220 4.300 ;
        RECT 108.380 1.770 109.460 4.300 ;
        RECT 110.620 1.770 111.700 4.300 ;
        RECT 112.860 1.770 113.940 4.300 ;
        RECT 115.100 1.770 116.180 4.300 ;
        RECT 117.340 1.770 118.420 4.300 ;
        RECT 119.580 1.770 120.660 4.300 ;
        RECT 121.820 1.770 122.900 4.300 ;
        RECT 124.060 1.770 125.140 4.300 ;
        RECT 126.300 1.770 127.380 4.300 ;
        RECT 128.540 1.770 129.620 4.300 ;
        RECT 130.780 1.770 131.860 4.300 ;
        RECT 133.020 1.770 134.100 4.300 ;
        RECT 135.260 1.770 136.340 4.300 ;
        RECT 137.500 1.770 138.580 4.300 ;
        RECT 139.740 1.770 140.820 4.300 ;
        RECT 141.980 1.770 143.060 4.300 ;
        RECT 144.220 1.770 145.300 4.300 ;
        RECT 146.460 1.770 147.540 4.300 ;
        RECT 148.700 1.770 149.780 4.300 ;
        RECT 150.940 1.770 152.020 4.300 ;
        RECT 153.180 1.770 154.260 4.300 ;
        RECT 155.420 1.770 156.500 4.300 ;
        RECT 157.660 1.770 158.740 4.300 ;
        RECT 159.900 1.770 160.980 4.300 ;
        RECT 162.140 1.770 163.220 4.300 ;
        RECT 164.380 1.770 165.460 4.300 ;
        RECT 166.620 1.770 167.700 4.300 ;
        RECT 168.860 1.770 169.940 4.300 ;
        RECT 171.100 1.770 172.180 4.300 ;
        RECT 173.340 1.770 174.420 4.300 ;
        RECT 175.580 1.770 176.660 4.300 ;
        RECT 177.820 1.770 178.900 4.300 ;
        RECT 180.060 1.770 181.140 4.300 ;
        RECT 182.300 1.770 183.380 4.300 ;
        RECT 184.540 1.770 185.620 4.300 ;
        RECT 186.780 1.770 187.860 4.300 ;
        RECT 189.020 1.770 190.100 4.300 ;
        RECT 191.260 1.770 192.340 4.300 ;
        RECT 193.500 1.770 194.580 4.300 ;
        RECT 195.740 1.770 196.820 4.300 ;
        RECT 197.980 1.770 199.060 4.300 ;
        RECT 200.220 1.770 201.300 4.300 ;
        RECT 202.460 1.770 203.540 4.300 ;
        RECT 204.700 1.770 205.780 4.300 ;
        RECT 206.940 1.770 208.020 4.300 ;
        RECT 209.180 1.770 210.260 4.300 ;
        RECT 211.420 1.770 212.500 4.300 ;
        RECT 213.660 1.770 214.740 4.300 ;
        RECT 215.900 1.770 216.980 4.300 ;
        RECT 218.140 1.770 219.220 4.300 ;
        RECT 220.380 1.770 221.460 4.300 ;
        RECT 222.620 1.770 223.700 4.300 ;
        RECT 224.860 1.770 225.940 4.300 ;
        RECT 227.100 1.770 228.180 4.300 ;
        RECT 229.340 1.770 230.420 4.300 ;
        RECT 231.580 1.770 232.660 4.300 ;
        RECT 233.820 1.770 234.900 4.300 ;
        RECT 236.060 1.770 237.140 4.300 ;
        RECT 238.300 1.770 239.380 4.300 ;
        RECT 240.540 1.770 241.620 4.300 ;
        RECT 242.780 1.770 243.860 4.300 ;
        RECT 245.020 1.770 246.100 4.300 ;
        RECT 247.260 1.770 248.340 4.300 ;
        RECT 249.500 1.770 250.580 4.300 ;
        RECT 251.740 1.770 252.820 4.300 ;
        RECT 253.980 1.770 255.060 4.300 ;
        RECT 256.220 1.770 257.300 4.300 ;
        RECT 258.460 1.770 259.540 4.300 ;
        RECT 260.700 1.770 261.780 4.300 ;
        RECT 262.940 1.770 264.020 4.300 ;
        RECT 265.180 1.770 266.260 4.300 ;
        RECT 267.420 1.770 268.500 4.300 ;
        RECT 269.660 1.770 270.740 4.300 ;
        RECT 271.900 1.770 272.980 4.300 ;
        RECT 274.140 1.770 275.220 4.300 ;
        RECT 276.380 1.770 277.460 4.300 ;
        RECT 278.620 1.770 279.700 4.300 ;
        RECT 280.860 1.770 281.940 4.300 ;
        RECT 283.100 1.770 284.180 4.300 ;
        RECT 285.340 1.770 286.420 4.300 ;
        RECT 287.580 1.770 288.660 4.300 ;
        RECT 289.820 1.770 290.900 4.300 ;
        RECT 292.060 1.770 293.140 4.300 ;
        RECT 294.300 1.770 295.380 4.300 ;
        RECT 296.540 1.770 297.620 4.300 ;
        RECT 298.780 1.770 299.860 4.300 ;
        RECT 301.020 1.770 302.100 4.300 ;
        RECT 303.260 1.770 304.340 4.300 ;
        RECT 305.500 1.770 306.580 4.300 ;
        RECT 307.740 1.770 308.820 4.300 ;
        RECT 309.980 1.770 311.060 4.300 ;
        RECT 312.220 1.770 313.300 4.300 ;
        RECT 314.460 1.770 315.540 4.300 ;
        RECT 316.700 1.770 317.780 4.300 ;
        RECT 318.940 1.770 320.020 4.300 ;
        RECT 321.180 1.770 322.260 4.300 ;
        RECT 323.420 1.770 324.500 4.300 ;
        RECT 325.660 1.770 326.740 4.300 ;
        RECT 327.900 1.770 328.980 4.300 ;
        RECT 330.140 1.770 331.220 4.300 ;
        RECT 332.380 1.770 333.460 4.300 ;
        RECT 334.620 1.770 335.700 4.300 ;
        RECT 336.860 1.770 337.940 4.300 ;
        RECT 339.100 1.770 340.180 4.300 ;
        RECT 341.340 1.770 342.420 4.300 ;
        RECT 343.580 1.770 344.660 4.300 ;
        RECT 345.820 1.770 346.900 4.300 ;
        RECT 348.060 1.770 349.140 4.300 ;
        RECT 350.300 1.770 351.380 4.300 ;
        RECT 352.540 1.770 353.620 4.300 ;
        RECT 354.780 1.770 355.860 4.300 ;
        RECT 357.020 1.770 358.100 4.300 ;
        RECT 359.260 1.770 360.340 4.300 ;
        RECT 361.500 1.770 362.580 4.300 ;
        RECT 363.740 1.770 364.820 4.300 ;
        RECT 365.980 1.770 367.060 4.300 ;
        RECT 368.220 1.770 369.300 4.300 ;
        RECT 370.460 1.770 371.540 4.300 ;
        RECT 372.700 1.770 373.780 4.300 ;
        RECT 374.940 1.770 376.020 4.300 ;
        RECT 377.180 1.770 378.260 4.300 ;
        RECT 379.420 1.770 380.500 4.300 ;
        RECT 381.660 1.770 382.740 4.300 ;
        RECT 383.900 1.770 384.980 4.300 ;
        RECT 386.140 1.770 387.220 4.300 ;
        RECT 388.380 1.770 389.460 4.300 ;
        RECT 390.620 1.770 391.700 4.300 ;
        RECT 392.860 1.770 393.940 4.300 ;
        RECT 395.100 1.770 396.180 4.300 ;
        RECT 397.340 1.770 398.420 4.300 ;
        RECT 399.580 1.770 400.660 4.300 ;
        RECT 401.820 1.770 402.900 4.300 ;
        RECT 404.060 1.770 405.140 4.300 ;
        RECT 406.300 1.770 407.380 4.300 ;
        RECT 408.540 1.770 409.620 4.300 ;
        RECT 410.780 1.770 411.860 4.300 ;
        RECT 413.020 1.770 414.100 4.300 ;
        RECT 415.260 1.770 416.340 4.300 ;
        RECT 417.500 1.770 418.580 4.300 ;
        RECT 419.740 1.770 420.820 4.300 ;
        RECT 421.980 1.770 423.060 4.300 ;
        RECT 424.220 1.770 425.300 4.300 ;
        RECT 426.460 1.770 427.540 4.300 ;
        RECT 428.700 1.770 429.780 4.300 ;
        RECT 430.940 1.770 432.020 4.300 ;
        RECT 433.180 1.770 434.260 4.300 ;
        RECT 435.420 1.770 436.500 4.300 ;
        RECT 437.660 1.770 438.740 4.300 ;
        RECT 439.900 1.770 440.980 4.300 ;
        RECT 442.140 1.770 443.220 4.300 ;
        RECT 444.380 1.770 445.460 4.300 ;
        RECT 446.620 1.770 447.700 4.300 ;
        RECT 448.860 1.770 449.940 4.300 ;
        RECT 451.100 1.770 452.180 4.300 ;
        RECT 453.340 1.770 454.420 4.300 ;
        RECT 455.580 1.770 456.660 4.300 ;
        RECT 457.820 1.770 458.900 4.300 ;
        RECT 460.060 1.770 461.140 4.300 ;
        RECT 462.300 1.770 463.380 4.300 ;
        RECT 464.540 1.770 465.620 4.300 ;
        RECT 466.780 1.770 467.860 4.300 ;
        RECT 469.020 1.770 470.100 4.300 ;
        RECT 471.260 1.770 472.340 4.300 ;
        RECT 473.500 1.770 474.580 4.300 ;
        RECT 475.740 1.770 476.820 4.300 ;
        RECT 477.980 1.770 479.060 4.300 ;
        RECT 480.220 1.770 481.300 4.300 ;
        RECT 482.460 1.770 483.540 4.300 ;
        RECT 484.700 1.770 485.780 4.300 ;
        RECT 486.940 1.770 488.020 4.300 ;
        RECT 489.180 1.770 490.260 4.300 ;
        RECT 491.420 1.770 492.500 4.300 ;
        RECT 493.660 1.770 494.740 4.300 ;
        RECT 495.900 1.770 496.980 4.300 ;
        RECT 498.140 1.770 499.220 4.300 ;
        RECT 500.380 1.770 501.460 4.300 ;
        RECT 502.620 1.770 503.700 4.300 ;
        RECT 504.860 1.770 505.940 4.300 ;
        RECT 507.100 1.770 508.180 4.300 ;
        RECT 509.340 1.770 510.420 4.300 ;
        RECT 511.580 1.770 512.660 4.300 ;
        RECT 513.820 1.770 514.900 4.300 ;
        RECT 516.060 1.770 517.140 4.300 ;
        RECT 518.300 1.770 519.380 4.300 ;
        RECT 520.540 1.770 521.620 4.300 ;
        RECT 522.780 1.770 523.860 4.300 ;
        RECT 525.020 1.770 526.100 4.300 ;
        RECT 527.260 1.770 528.340 4.300 ;
        RECT 529.500 1.770 530.580 4.300 ;
        RECT 531.740 1.770 532.820 4.300 ;
        RECT 533.980 1.770 535.060 4.300 ;
        RECT 536.220 1.770 537.300 4.300 ;
        RECT 538.460 1.770 539.540 4.300 ;
        RECT 540.700 1.770 541.780 4.300 ;
        RECT 542.940 1.770 544.020 4.300 ;
        RECT 545.180 1.770 546.260 4.300 ;
        RECT 547.420 1.770 548.500 4.300 ;
        RECT 549.660 1.770 550.740 4.300 ;
        RECT 551.900 1.770 552.980 4.300 ;
        RECT 554.140 1.770 555.220 4.300 ;
        RECT 556.380 1.770 557.460 4.300 ;
        RECT 558.620 1.770 559.700 4.300 ;
        RECT 560.860 1.770 561.940 4.300 ;
        RECT 563.100 1.770 564.180 4.300 ;
        RECT 565.340 1.770 566.420 4.300 ;
        RECT 567.580 1.770 568.660 4.300 ;
        RECT 569.820 1.770 570.900 4.300 ;
        RECT 572.060 1.770 573.140 4.300 ;
        RECT 574.300 1.770 575.380 4.300 ;
        RECT 576.540 1.770 577.620 4.300 ;
        RECT 578.780 1.770 579.860 4.300 ;
        RECT 581.020 1.770 582.100 4.300 ;
        RECT 583.260 1.770 584.340 4.300 ;
        RECT 585.500 1.770 586.580 4.300 ;
        RECT 587.740 1.770 588.820 4.300 ;
        RECT 589.980 1.770 591.060 4.300 ;
        RECT 592.220 1.770 593.300 4.300 ;
        RECT 594.460 1.770 595.540 4.300 ;
        RECT 596.700 1.770 597.780 4.300 ;
        RECT 598.940 1.770 600.020 4.300 ;
        RECT 601.180 1.770 602.260 4.300 ;
        RECT 603.420 1.770 604.500 4.300 ;
        RECT 605.660 1.770 606.740 4.300 ;
        RECT 607.900 1.770 608.980 4.300 ;
        RECT 610.140 1.770 611.220 4.300 ;
        RECT 612.380 1.770 613.460 4.300 ;
        RECT 614.620 1.770 615.700 4.300 ;
        RECT 616.860 1.770 617.940 4.300 ;
        RECT 619.100 1.770 620.180 4.300 ;
        RECT 621.340 1.770 622.420 4.300 ;
        RECT 623.580 1.770 624.660 4.300 ;
        RECT 625.820 1.770 626.900 4.300 ;
        RECT 628.060 1.770 629.140 4.300 ;
        RECT 630.300 1.770 631.380 4.300 ;
        RECT 632.540 1.770 633.620 4.300 ;
        RECT 634.780 1.770 635.860 4.300 ;
        RECT 637.020 1.770 638.100 4.300 ;
        RECT 639.260 1.770 640.340 4.300 ;
        RECT 641.500 1.770 642.580 4.300 ;
        RECT 643.740 1.770 644.820 4.300 ;
        RECT 645.980 1.770 647.060 4.300 ;
        RECT 648.220 1.770 649.300 4.300 ;
        RECT 650.460 1.770 651.540 4.300 ;
        RECT 652.700 1.770 653.780 4.300 ;
        RECT 654.940 1.770 656.020 4.300 ;
        RECT 657.180 1.770 658.260 4.300 ;
        RECT 659.420 1.770 660.500 4.300 ;
        RECT 661.660 1.770 662.740 4.300 ;
        RECT 663.900 1.770 664.980 4.300 ;
        RECT 666.140 1.770 667.220 4.300 ;
        RECT 668.380 1.770 669.460 4.300 ;
        RECT 670.620 1.770 671.700 4.300 ;
        RECT 672.860 1.770 673.940 4.300 ;
        RECT 675.100 1.770 676.180 4.300 ;
        RECT 677.340 1.770 678.420 4.300 ;
        RECT 679.580 1.770 680.660 4.300 ;
        RECT 681.820 1.770 682.900 4.300 ;
        RECT 684.060 1.770 685.140 4.300 ;
        RECT 686.300 1.770 687.380 4.300 ;
        RECT 688.540 1.770 689.620 4.300 ;
        RECT 690.780 1.770 691.860 4.300 ;
        RECT 693.020 1.770 694.100 4.300 ;
        RECT 695.260 1.770 696.340 4.300 ;
        RECT 697.500 1.770 698.580 4.300 ;
        RECT 699.740 1.770 700.820 4.300 ;
        RECT 701.980 1.770 703.060 4.300 ;
        RECT 704.220 1.770 705.300 4.300 ;
        RECT 706.460 1.770 707.540 4.300 ;
        RECT 708.700 1.770 709.780 4.300 ;
        RECT 710.940 1.770 712.020 4.300 ;
        RECT 713.180 1.770 714.260 4.300 ;
        RECT 715.420 1.770 716.500 4.300 ;
        RECT 717.660 1.770 718.740 4.300 ;
        RECT 719.900 1.770 720.980 4.300 ;
        RECT 722.140 1.770 723.220 4.300 ;
        RECT 724.380 1.770 725.460 4.300 ;
        RECT 726.620 1.770 727.700 4.300 ;
        RECT 728.860 1.770 729.940 4.300 ;
        RECT 731.100 1.770 732.180 4.300 ;
        RECT 733.340 1.770 734.420 4.300 ;
        RECT 735.580 1.770 736.660 4.300 ;
        RECT 737.820 1.770 738.900 4.300 ;
        RECT 740.060 1.770 741.140 4.300 ;
        RECT 742.300 1.770 743.380 4.300 ;
        RECT 744.540 1.770 745.620 4.300 ;
        RECT 746.780 1.770 747.860 4.300 ;
        RECT 749.020 1.770 750.100 4.300 ;
        RECT 751.260 1.770 752.340 4.300 ;
        RECT 753.500 1.770 754.580 4.300 ;
        RECT 755.740 1.770 756.820 4.300 ;
        RECT 757.980 1.770 759.060 4.300 ;
        RECT 760.220 1.770 761.300 4.300 ;
        RECT 762.460 1.770 763.540 4.300 ;
        RECT 764.700 1.770 765.780 4.300 ;
        RECT 766.940 1.770 768.020 4.300 ;
        RECT 769.180 1.770 770.260 4.300 ;
        RECT 771.420 1.770 772.500 4.300 ;
        RECT 773.660 1.770 774.740 4.300 ;
        RECT 775.900 1.770 776.980 4.300 ;
        RECT 778.140 1.770 779.220 4.300 ;
        RECT 780.380 1.770 781.460 4.300 ;
        RECT 782.620 1.770 783.700 4.300 ;
        RECT 784.860 1.770 785.940 4.300 ;
        RECT 787.100 1.770 788.180 4.300 ;
        RECT 789.340 1.770 790.420 4.300 ;
        RECT 791.580 1.770 792.660 4.300 ;
        RECT 793.820 1.770 794.900 4.300 ;
        RECT 796.060 1.770 797.140 4.300 ;
        RECT 798.300 1.770 799.380 4.300 ;
        RECT 800.540 1.770 801.620 4.300 ;
        RECT 802.780 1.770 803.860 4.300 ;
        RECT 805.020 1.770 806.100 4.300 ;
        RECT 807.260 1.770 808.340 4.300 ;
        RECT 809.500 1.770 810.580 4.300 ;
        RECT 811.740 1.770 812.820 4.300 ;
        RECT 813.980 1.770 815.060 4.300 ;
        RECT 816.220 1.770 817.300 4.300 ;
        RECT 818.460 1.770 819.540 4.300 ;
        RECT 820.700 1.770 821.780 4.300 ;
        RECT 822.940 1.770 824.020 4.300 ;
        RECT 825.180 1.770 826.260 4.300 ;
        RECT 827.420 1.770 828.500 4.300 ;
        RECT 829.660 1.770 830.740 4.300 ;
        RECT 831.900 1.770 832.980 4.300 ;
        RECT 834.140 1.770 835.220 4.300 ;
        RECT 836.380 1.770 837.460 4.300 ;
        RECT 838.620 1.770 839.700 4.300 ;
        RECT 840.860 1.770 841.940 4.300 ;
        RECT 843.100 1.770 844.180 4.300 ;
        RECT 845.340 1.770 846.420 4.300 ;
        RECT 847.580 1.770 848.660 4.300 ;
        RECT 849.820 1.770 850.900 4.300 ;
        RECT 852.060 1.770 853.140 4.300 ;
        RECT 854.300 1.770 855.380 4.300 ;
        RECT 856.540 1.770 857.620 4.300 ;
        RECT 858.780 1.770 859.860 4.300 ;
        RECT 861.020 1.770 862.100 4.300 ;
        RECT 863.260 1.770 864.340 4.300 ;
        RECT 865.500 1.770 866.580 4.300 ;
        RECT 867.740 1.770 868.820 4.300 ;
        RECT 869.980 1.770 871.060 4.300 ;
        RECT 872.220 1.770 873.300 4.300 ;
        RECT 874.460 1.770 875.540 4.300 ;
        RECT 876.700 1.770 877.780 4.300 ;
        RECT 878.940 1.770 880.020 4.300 ;
        RECT 881.180 1.770 882.260 4.300 ;
        RECT 883.420 1.770 884.500 4.300 ;
        RECT 885.660 1.770 886.740 4.300 ;
        RECT 887.900 1.770 888.980 4.300 ;
        RECT 890.140 1.770 891.220 4.300 ;
        RECT 892.380 1.770 893.460 4.300 ;
        RECT 894.620 1.770 895.700 4.300 ;
        RECT 896.860 1.770 897.940 4.300 ;
        RECT 899.100 1.770 900.180 4.300 ;
        RECT 901.340 1.770 902.420 4.300 ;
        RECT 903.580 1.770 904.660 4.300 ;
        RECT 905.820 1.770 906.900 4.300 ;
        RECT 908.060 1.770 909.140 4.300 ;
        RECT 910.300 1.770 911.380 4.300 ;
        RECT 912.540 1.770 913.620 4.300 ;
        RECT 914.780 1.770 915.860 4.300 ;
        RECT 917.020 1.770 918.100 4.300 ;
        RECT 919.260 1.770 920.340 4.300 ;
        RECT 921.500 1.770 922.580 4.300 ;
        RECT 923.740 1.770 924.820 4.300 ;
        RECT 925.980 1.770 927.060 4.300 ;
        RECT 928.220 1.770 929.300 4.300 ;
        RECT 930.460 1.770 931.540 4.300 ;
        RECT 932.700 1.770 933.780 4.300 ;
        RECT 934.940 1.770 936.020 4.300 ;
        RECT 937.180 1.770 938.260 4.300 ;
        RECT 939.420 1.770 940.500 4.300 ;
        RECT 941.660 1.770 942.740 4.300 ;
        RECT 943.900 1.770 944.980 4.300 ;
        RECT 946.140 1.770 947.220 4.300 ;
        RECT 948.380 1.770 949.460 4.300 ;
        RECT 950.620 1.770 951.700 4.300 ;
        RECT 952.860 1.770 953.940 4.300 ;
        RECT 955.100 1.770 956.180 4.300 ;
        RECT 957.340 1.770 958.420 4.300 ;
        RECT 959.580 1.770 960.660 4.300 ;
        RECT 961.820 1.770 962.900 4.300 ;
        RECT 964.060 1.770 965.140 4.300 ;
        RECT 966.300 1.770 967.380 4.300 ;
        RECT 968.540 1.770 969.620 4.300 ;
        RECT 970.780 1.770 971.860 4.300 ;
        RECT 973.020 1.770 974.100 4.300 ;
        RECT 975.260 1.770 976.340 4.300 ;
        RECT 977.500 1.770 978.580 4.300 ;
        RECT 979.740 1.770 980.820 4.300 ;
        RECT 981.980 1.770 983.060 4.300 ;
        RECT 984.220 1.770 985.300 4.300 ;
        RECT 986.460 1.770 987.540 4.300 ;
        RECT 988.700 1.770 989.780 4.300 ;
        RECT 990.940 1.770 992.020 4.300 ;
        RECT 993.180 1.770 994.260 4.300 ;
        RECT 995.420 1.770 996.500 4.300 ;
        RECT 997.660 1.770 998.740 4.300 ;
        RECT 999.900 1.770 1000.980 4.300 ;
        RECT 1002.140 1.770 1003.220 4.300 ;
        RECT 1004.380 1.770 1005.460 4.300 ;
        RECT 1006.620 1.770 1007.700 4.300 ;
        RECT 1008.860 1.770 1009.940 4.300 ;
        RECT 1011.100 1.770 1012.180 4.300 ;
        RECT 1013.340 1.770 1014.420 4.300 ;
        RECT 1015.580 1.770 1016.660 4.300 ;
        RECT 1017.820 1.770 1018.900 4.300 ;
        RECT 1020.060 1.770 1021.140 4.300 ;
        RECT 1022.300 1.770 1023.380 4.300 ;
        RECT 1024.540 1.770 1025.620 4.300 ;
        RECT 1026.780 1.770 1027.860 4.300 ;
        RECT 1029.020 1.770 1030.100 4.300 ;
        RECT 1031.260 1.770 1032.340 4.300 ;
        RECT 1033.500 1.770 1034.580 4.300 ;
        RECT 1035.740 1.770 1036.820 4.300 ;
        RECT 1037.980 1.770 1039.060 4.300 ;
        RECT 1040.220 1.770 1041.300 4.300 ;
        RECT 1042.460 1.770 1043.540 4.300 ;
        RECT 1044.700 1.770 1045.780 4.300 ;
        RECT 1046.940 1.770 1048.020 4.300 ;
        RECT 1049.180 1.770 1050.260 4.300 ;
        RECT 1051.420 1.770 1052.500 4.300 ;
        RECT 1053.660 1.770 1054.740 4.300 ;
        RECT 1055.900 1.770 1056.980 4.300 ;
        RECT 1058.140 1.770 1059.220 4.300 ;
        RECT 1060.380 1.770 1061.460 4.300 ;
        RECT 1062.620 1.770 1063.700 4.300 ;
        RECT 1064.860 1.770 1065.940 4.300 ;
        RECT 1067.100 1.770 1068.180 4.300 ;
        RECT 1069.340 1.770 1070.420 4.300 ;
        RECT 1071.580 1.770 1072.660 4.300 ;
        RECT 1073.820 1.770 1074.900 4.300 ;
        RECT 1076.060 1.770 1077.140 4.300 ;
        RECT 1078.300 1.770 1079.380 4.300 ;
        RECT 1080.540 1.770 1081.620 4.300 ;
        RECT 1082.780 1.770 1083.860 4.300 ;
        RECT 1085.020 1.770 1086.100 4.300 ;
        RECT 1087.260 1.770 1088.340 4.300 ;
        RECT 1089.500 1.770 1090.580 4.300 ;
        RECT 1091.740 1.770 1092.820 4.300 ;
        RECT 1093.980 1.770 1095.060 4.300 ;
        RECT 1096.220 1.770 1097.300 4.300 ;
        RECT 1098.460 1.770 1099.540 4.300 ;
        RECT 1100.700 1.770 1101.780 4.300 ;
        RECT 1102.940 1.770 1104.020 4.300 ;
        RECT 1105.180 1.770 1106.260 4.300 ;
        RECT 1107.420 1.770 1108.500 4.300 ;
        RECT 1109.660 1.770 1110.740 4.300 ;
        RECT 1111.900 1.770 1112.980 4.300 ;
        RECT 1114.140 1.770 1115.220 4.300 ;
        RECT 1116.380 1.770 1117.460 4.300 ;
        RECT 1118.620 1.770 1119.700 4.300 ;
        RECT 1120.860 1.770 1121.940 4.300 ;
        RECT 1123.100 1.770 1124.180 4.300 ;
        RECT 1125.340 1.770 1126.420 4.300 ;
        RECT 1127.580 1.770 1128.660 4.300 ;
        RECT 1129.820 1.770 1130.900 4.300 ;
        RECT 1132.060 1.770 1133.140 4.300 ;
        RECT 1134.300 1.770 1135.380 4.300 ;
        RECT 1136.540 1.770 1137.620 4.300 ;
        RECT 1138.780 1.770 1139.860 4.300 ;
        RECT 1141.020 1.770 1142.100 4.300 ;
        RECT 1143.260 1.770 1144.340 4.300 ;
        RECT 1145.500 1.770 1146.580 4.300 ;
        RECT 1147.740 1.770 1148.820 4.300 ;
        RECT 1149.980 1.770 1193.220 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 327.900 1196.000 340.340 ;
        RECT 4.300 326.740 1195.700 327.900 ;
        RECT 4.000 324.540 1196.000 326.740 ;
        RECT 4.300 323.380 1195.700 324.540 ;
        RECT 4.000 321.180 1196.000 323.380 ;
        RECT 4.300 320.020 1195.700 321.180 ;
        RECT 4.000 317.820 1196.000 320.020 ;
        RECT 4.300 316.660 1195.700 317.820 ;
        RECT 4.000 314.460 1196.000 316.660 ;
        RECT 4.300 313.300 1195.700 314.460 ;
        RECT 4.000 311.100 1196.000 313.300 ;
        RECT 4.300 309.940 1195.700 311.100 ;
        RECT 4.000 307.740 1196.000 309.940 ;
        RECT 4.300 306.580 1195.700 307.740 ;
        RECT 4.000 304.380 1196.000 306.580 ;
        RECT 4.300 303.220 1195.700 304.380 ;
        RECT 4.000 301.020 1196.000 303.220 ;
        RECT 4.300 299.860 1195.700 301.020 ;
        RECT 4.000 297.660 1196.000 299.860 ;
        RECT 4.300 296.500 1195.700 297.660 ;
        RECT 4.000 294.300 1196.000 296.500 ;
        RECT 4.300 293.140 1195.700 294.300 ;
        RECT 4.000 290.940 1196.000 293.140 ;
        RECT 4.300 289.780 1195.700 290.940 ;
        RECT 4.000 287.580 1196.000 289.780 ;
        RECT 4.300 286.420 1195.700 287.580 ;
        RECT 4.000 284.220 1196.000 286.420 ;
        RECT 4.300 283.060 1195.700 284.220 ;
        RECT 4.000 280.860 1196.000 283.060 ;
        RECT 4.300 279.700 1195.700 280.860 ;
        RECT 4.000 277.500 1196.000 279.700 ;
        RECT 4.300 276.340 1195.700 277.500 ;
        RECT 4.000 274.140 1196.000 276.340 ;
        RECT 4.300 272.980 1195.700 274.140 ;
        RECT 4.000 270.780 1196.000 272.980 ;
        RECT 4.300 269.620 1195.700 270.780 ;
        RECT 4.000 267.420 1196.000 269.620 ;
        RECT 4.300 266.260 1195.700 267.420 ;
        RECT 4.000 264.060 1196.000 266.260 ;
        RECT 4.300 262.900 1195.700 264.060 ;
        RECT 4.000 260.700 1196.000 262.900 ;
        RECT 4.300 259.540 1195.700 260.700 ;
        RECT 4.000 257.340 1196.000 259.540 ;
        RECT 4.300 256.180 1195.700 257.340 ;
        RECT 4.000 253.980 1196.000 256.180 ;
        RECT 4.300 252.820 1195.700 253.980 ;
        RECT 4.000 250.620 1196.000 252.820 ;
        RECT 4.300 249.460 1195.700 250.620 ;
        RECT 4.000 247.260 1196.000 249.460 ;
        RECT 4.300 246.100 1195.700 247.260 ;
        RECT 4.000 243.900 1196.000 246.100 ;
        RECT 4.300 242.740 1195.700 243.900 ;
        RECT 4.000 240.540 1196.000 242.740 ;
        RECT 4.300 239.380 1195.700 240.540 ;
        RECT 4.000 237.180 1196.000 239.380 ;
        RECT 4.300 236.020 1195.700 237.180 ;
        RECT 4.000 233.820 1196.000 236.020 ;
        RECT 4.300 232.660 1195.700 233.820 ;
        RECT 4.000 230.460 1196.000 232.660 ;
        RECT 4.300 229.300 1195.700 230.460 ;
        RECT 4.000 227.100 1196.000 229.300 ;
        RECT 4.300 225.940 1195.700 227.100 ;
        RECT 4.000 223.740 1196.000 225.940 ;
        RECT 4.300 222.580 1195.700 223.740 ;
        RECT 4.000 220.380 1196.000 222.580 ;
        RECT 4.300 219.220 1195.700 220.380 ;
        RECT 4.000 217.020 1196.000 219.220 ;
        RECT 4.300 215.860 1195.700 217.020 ;
        RECT 4.000 213.660 1196.000 215.860 ;
        RECT 4.300 212.500 1195.700 213.660 ;
        RECT 4.000 210.300 1196.000 212.500 ;
        RECT 4.300 209.140 1195.700 210.300 ;
        RECT 4.000 206.940 1196.000 209.140 ;
        RECT 4.300 205.780 1195.700 206.940 ;
        RECT 4.000 203.580 1196.000 205.780 ;
        RECT 4.300 202.420 1195.700 203.580 ;
        RECT 4.000 200.220 1196.000 202.420 ;
        RECT 4.300 199.060 1195.700 200.220 ;
        RECT 4.000 196.860 1196.000 199.060 ;
        RECT 4.300 195.700 1195.700 196.860 ;
        RECT 4.000 193.500 1196.000 195.700 ;
        RECT 4.300 192.340 1195.700 193.500 ;
        RECT 4.000 190.140 1196.000 192.340 ;
        RECT 4.300 188.980 1195.700 190.140 ;
        RECT 4.000 186.780 1196.000 188.980 ;
        RECT 4.300 185.620 1195.700 186.780 ;
        RECT 4.000 183.420 1196.000 185.620 ;
        RECT 4.300 182.260 1195.700 183.420 ;
        RECT 4.000 180.060 1196.000 182.260 ;
        RECT 4.300 178.900 1195.700 180.060 ;
        RECT 4.000 176.700 1196.000 178.900 ;
        RECT 4.300 175.540 1195.700 176.700 ;
        RECT 4.000 173.340 1196.000 175.540 ;
        RECT 4.300 172.180 1195.700 173.340 ;
        RECT 4.000 169.980 1196.000 172.180 ;
        RECT 4.300 168.820 1195.700 169.980 ;
        RECT 4.000 166.620 1196.000 168.820 ;
        RECT 4.300 165.460 1195.700 166.620 ;
        RECT 4.000 163.260 1196.000 165.460 ;
        RECT 4.300 162.100 1195.700 163.260 ;
        RECT 4.000 159.900 1196.000 162.100 ;
        RECT 4.300 158.740 1195.700 159.900 ;
        RECT 4.000 156.540 1196.000 158.740 ;
        RECT 4.300 155.380 1195.700 156.540 ;
        RECT 4.000 153.180 1196.000 155.380 ;
        RECT 4.300 152.020 1195.700 153.180 ;
        RECT 4.000 149.820 1196.000 152.020 ;
        RECT 4.300 148.660 1195.700 149.820 ;
        RECT 4.000 146.460 1196.000 148.660 ;
        RECT 4.300 145.300 1195.700 146.460 ;
        RECT 4.000 143.100 1196.000 145.300 ;
        RECT 4.300 141.940 1195.700 143.100 ;
        RECT 4.000 139.740 1196.000 141.940 ;
        RECT 4.300 138.580 1195.700 139.740 ;
        RECT 4.000 136.380 1196.000 138.580 ;
        RECT 4.300 135.220 1195.700 136.380 ;
        RECT 4.000 133.020 1196.000 135.220 ;
        RECT 4.300 131.860 1195.700 133.020 ;
        RECT 4.000 129.660 1196.000 131.860 ;
        RECT 4.300 128.500 1195.700 129.660 ;
        RECT 4.000 126.300 1196.000 128.500 ;
        RECT 4.300 125.140 1195.700 126.300 ;
        RECT 4.000 122.940 1196.000 125.140 ;
        RECT 4.300 121.780 1195.700 122.940 ;
        RECT 4.000 119.580 1196.000 121.780 ;
        RECT 4.300 118.420 1195.700 119.580 ;
        RECT 4.000 116.220 1196.000 118.420 ;
        RECT 4.300 115.060 1195.700 116.220 ;
        RECT 4.000 112.860 1196.000 115.060 ;
        RECT 4.300 111.700 1195.700 112.860 ;
        RECT 4.000 109.500 1196.000 111.700 ;
        RECT 4.300 108.340 1195.700 109.500 ;
        RECT 4.000 106.140 1196.000 108.340 ;
        RECT 4.300 104.980 1195.700 106.140 ;
        RECT 4.000 102.780 1196.000 104.980 ;
        RECT 4.300 101.620 1195.700 102.780 ;
        RECT 4.000 99.420 1196.000 101.620 ;
        RECT 4.300 98.260 1195.700 99.420 ;
        RECT 4.000 96.060 1196.000 98.260 ;
        RECT 4.300 94.900 1195.700 96.060 ;
        RECT 4.000 92.700 1196.000 94.900 ;
        RECT 4.300 91.540 1195.700 92.700 ;
        RECT 4.000 89.340 1196.000 91.540 ;
        RECT 4.300 88.180 1195.700 89.340 ;
        RECT 4.000 85.980 1196.000 88.180 ;
        RECT 4.300 84.820 1195.700 85.980 ;
        RECT 4.000 82.620 1196.000 84.820 ;
        RECT 4.300 81.460 1195.700 82.620 ;
        RECT 4.000 79.260 1196.000 81.460 ;
        RECT 4.300 78.100 1195.700 79.260 ;
        RECT 4.000 75.900 1196.000 78.100 ;
        RECT 4.300 74.740 1195.700 75.900 ;
        RECT 4.000 72.540 1196.000 74.740 ;
        RECT 4.300 71.380 1195.700 72.540 ;
        RECT 4.000 69.180 1196.000 71.380 ;
        RECT 4.300 68.020 1195.700 69.180 ;
        RECT 4.000 65.820 1196.000 68.020 ;
        RECT 4.300 64.660 1195.700 65.820 ;
        RECT 4.000 62.460 1196.000 64.660 ;
        RECT 4.300 61.300 1195.700 62.460 ;
        RECT 4.000 59.100 1196.000 61.300 ;
        RECT 4.300 57.940 1195.700 59.100 ;
        RECT 4.000 55.740 1196.000 57.940 ;
        RECT 4.300 54.580 1195.700 55.740 ;
        RECT 4.000 52.380 1196.000 54.580 ;
        RECT 4.300 51.220 1195.700 52.380 ;
        RECT 4.000 49.020 1196.000 51.220 ;
        RECT 4.300 47.860 1195.700 49.020 ;
        RECT 4.000 45.660 1196.000 47.860 ;
        RECT 4.300 44.500 1195.700 45.660 ;
        RECT 4.000 42.300 1196.000 44.500 ;
        RECT 4.300 41.140 1195.700 42.300 ;
        RECT 4.000 38.940 1196.000 41.140 ;
        RECT 4.300 37.780 1195.700 38.940 ;
        RECT 4.000 35.580 1196.000 37.780 ;
        RECT 4.300 34.420 1195.700 35.580 ;
        RECT 4.000 32.220 1196.000 34.420 ;
        RECT 4.300 31.060 1195.700 32.220 ;
        RECT 4.000 28.860 1196.000 31.060 ;
        RECT 4.300 27.700 1195.700 28.860 ;
        RECT 4.000 25.500 1196.000 27.700 ;
        RECT 4.300 24.340 1195.700 25.500 ;
        RECT 4.000 22.140 1196.000 24.340 ;
        RECT 4.300 20.980 1195.700 22.140 ;
        RECT 4.000 1.820 1196.000 20.980 ;
      LAYER Metal4 ;
        RECT 9.100 333.800 1182.020 337.590 ;
        RECT 9.100 15.080 21.940 333.800 ;
        RECT 24.140 15.080 98.740 333.800 ;
        RECT 100.940 15.080 175.540 333.800 ;
        RECT 177.740 15.080 252.340 333.800 ;
        RECT 254.540 15.080 329.140 333.800 ;
        RECT 331.340 15.080 405.940 333.800 ;
        RECT 408.140 15.080 482.740 333.800 ;
        RECT 484.940 15.080 559.540 333.800 ;
        RECT 561.740 15.080 636.340 333.800 ;
        RECT 638.540 15.080 713.140 333.800 ;
        RECT 715.340 15.080 789.940 333.800 ;
        RECT 792.140 15.080 866.740 333.800 ;
        RECT 868.940 15.080 943.540 333.800 ;
        RECT 945.740 15.080 1020.340 333.800 ;
        RECT 1022.540 15.080 1097.140 333.800 ;
        RECT 1099.340 15.080 1173.940 333.800 ;
        RECT 1176.140 15.080 1182.020 333.800 ;
        RECT 9.100 4.570 1182.020 15.080 ;
  END
END interconnect_inner
END LIBRARY

