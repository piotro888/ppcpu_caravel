magic
tech sky130B
magscale 1 2
timestamp 1663070773
<< viali >>
rect 8401 37417 8435 37451
rect 16129 37417 16163 37451
rect 31493 37281 31527 37315
rect 1869 37213 1903 37247
rect 2973 37213 3007 37247
rect 4077 37213 4111 37247
rect 5365 37213 5399 37247
rect 6561 37213 6595 37247
rect 7573 37213 7607 37247
rect 9137 37213 9171 37247
rect 9781 37213 9815 37247
rect 10885 37213 10919 37247
rect 11989 37213 12023 37247
rect 13093 37213 13127 37247
rect 14289 37213 14323 37247
rect 15301 37213 15335 37247
rect 16865 37213 16899 37247
rect 17509 37213 17543 37247
rect 18613 37213 18647 37247
rect 19717 37213 19751 37247
rect 20821 37213 20855 37247
rect 21833 37213 21867 37247
rect 23121 37213 23155 37247
rect 23857 37213 23891 37247
rect 24409 37213 24443 37247
rect 25145 37213 25179 37247
rect 26157 37213 26191 37247
rect 27261 37213 27295 37247
rect 28365 37213 28399 37247
rect 29561 37213 29595 37247
rect 30573 37213 30607 37247
rect 32137 37213 32171 37247
rect 32873 37213 32907 37247
rect 33885 37213 33919 37247
rect 34989 37213 35023 37247
rect 36093 37213 36127 37247
rect 37289 37213 37323 37247
rect 1961 37077 1995 37111
rect 3157 37077 3191 37111
rect 4261 37077 4295 37111
rect 5181 37077 5215 37111
rect 6377 37077 6411 37111
rect 7389 37077 7423 37111
rect 8953 37077 8987 37111
rect 9597 37077 9631 37111
rect 10701 37077 10735 37111
rect 11805 37077 11839 37111
rect 12909 37077 12943 37111
rect 14105 37077 14139 37111
rect 15117 37077 15151 37111
rect 16681 37077 16715 37111
rect 17325 37077 17359 37111
rect 18429 37077 18463 37111
rect 19533 37077 19567 37111
rect 20637 37077 20671 37111
rect 22017 37077 22051 37111
rect 22937 37077 22971 37111
rect 24593 37077 24627 37111
rect 25329 37077 25363 37111
rect 26341 37077 26375 37111
rect 27445 37077 27479 37111
rect 28549 37077 28583 37111
rect 29745 37077 29779 37111
rect 30757 37077 30791 37111
rect 32321 37077 32355 37111
rect 33057 37077 33091 37111
rect 34069 37077 34103 37111
rect 35173 37077 35207 37111
rect 36277 37077 36311 37111
rect 37473 37077 37507 37111
rect 38025 37077 38059 37111
rect 1961 36873 1995 36907
rect 2881 36873 2915 36907
rect 3985 36873 4019 36907
rect 5089 36873 5123 36907
rect 6377 36873 6411 36907
rect 7297 36873 7331 36907
rect 9505 36873 9539 36907
rect 10609 36873 10643 36907
rect 11713 36873 11747 36907
rect 12817 36873 12851 36907
rect 13921 36873 13955 36907
rect 15025 36873 15059 36907
rect 17233 36873 17267 36907
rect 18337 36873 18371 36907
rect 19349 36873 19383 36907
rect 20545 36873 20579 36907
rect 38025 36873 38059 36907
rect 2145 36737 2179 36771
rect 37841 36737 37875 36771
rect 21833 36533 21867 36567
rect 22753 36533 22787 36567
rect 25053 36533 25087 36567
rect 26065 36533 26099 36567
rect 27169 36533 27203 36567
rect 28181 36533 28215 36567
rect 29377 36533 29411 36567
rect 30389 36533 30423 36567
rect 32781 36533 32815 36567
rect 33793 36533 33827 36567
rect 34805 36533 34839 36567
rect 35909 36533 35943 36567
rect 37381 36533 37415 36567
rect 1593 36329 1627 36363
rect 38025 36329 38059 36363
rect 37841 36125 37875 36159
rect 2329 35989 2363 36023
rect 37289 35989 37323 36023
rect 1869 30209 1903 30243
rect 2053 30073 2087 30107
rect 1593 29801 1627 29835
rect 10517 20825 10551 20859
rect 11069 20757 11103 20791
rect 11805 20757 11839 20791
rect 12725 20757 12759 20791
rect 13369 20757 13403 20791
rect 16589 20757 16623 20791
rect 10885 20553 10919 20587
rect 13277 20553 13311 20587
rect 14197 20553 14231 20587
rect 17049 20553 17083 20587
rect 17969 20553 18003 20587
rect 10057 20417 10091 20451
rect 12265 20417 12299 20451
rect 13369 20349 13403 20383
rect 13461 20349 13495 20383
rect 16037 20349 16071 20383
rect 17141 20349 17175 20383
rect 17233 20349 17267 20383
rect 9873 20213 9907 20247
rect 11989 20213 12023 20247
rect 12909 20213 12943 20247
rect 16681 20213 16715 20247
rect 4353 20009 4387 20043
rect 7849 20009 7883 20043
rect 14749 20009 14783 20043
rect 18153 20009 18187 20043
rect 10609 19873 10643 19907
rect 11713 19873 11747 19907
rect 13001 19873 13035 19907
rect 14105 19873 14139 19907
rect 17417 19873 17451 19907
rect 10333 19805 10367 19839
rect 11529 19805 11563 19839
rect 15393 19805 15427 19839
rect 17233 19805 17267 19839
rect 9505 19737 9539 19771
rect 11621 19737 11655 19771
rect 12725 19737 12759 19771
rect 17325 19737 17359 19771
rect 8309 19669 8343 19703
rect 9965 19669 9999 19703
rect 10425 19669 10459 19703
rect 11161 19669 11195 19703
rect 12357 19669 12391 19703
rect 12817 19669 12851 19703
rect 15209 19669 15243 19703
rect 16313 19669 16347 19703
rect 16865 19669 16899 19703
rect 3433 19465 3467 19499
rect 3801 19465 3835 19499
rect 7665 19465 7699 19499
rect 10241 19465 10275 19499
rect 10609 19465 10643 19499
rect 15761 19465 15795 19499
rect 16957 19465 16991 19499
rect 17325 19465 17359 19499
rect 18245 19465 18279 19499
rect 9781 19397 9815 19431
rect 13277 19397 13311 19431
rect 7757 19329 7791 19363
rect 8861 19329 8895 19363
rect 12265 19329 12299 19363
rect 15945 19329 15979 19363
rect 3893 19261 3927 19295
rect 4077 19261 4111 19295
rect 5089 19261 5123 19295
rect 7849 19261 7883 19295
rect 8953 19261 8987 19295
rect 9137 19261 9171 19295
rect 10701 19261 10735 19295
rect 10793 19261 10827 19295
rect 12357 19261 12391 19295
rect 12449 19261 12483 19295
rect 17417 19261 17451 19295
rect 17509 19261 17543 19295
rect 2973 19125 3007 19159
rect 7297 19125 7331 19159
rect 8493 19125 8527 19159
rect 11897 19125 11931 19159
rect 13829 19125 13863 19159
rect 6653 18921 6687 18955
rect 11621 18921 11655 18955
rect 12725 18921 12759 18955
rect 16773 18921 16807 18955
rect 17233 18921 17267 18955
rect 10333 18853 10367 18887
rect 4813 18785 4847 18819
rect 5917 18785 5951 18819
rect 7941 18785 7975 18819
rect 9229 18785 9263 18819
rect 4537 18717 4571 18751
rect 5733 18717 5767 18751
rect 7665 18717 7699 18751
rect 9873 18717 9907 18751
rect 10517 18717 10551 18751
rect 11161 18717 11195 18751
rect 11805 18717 11839 18751
rect 15853 18717 15887 18751
rect 3249 18649 3283 18683
rect 4629 18649 4663 18683
rect 5825 18649 5859 18683
rect 4169 18581 4203 18615
rect 5365 18581 5399 18615
rect 7297 18581 7331 18615
rect 7757 18581 7791 18615
rect 9689 18581 9723 18615
rect 10977 18581 11011 18615
rect 15669 18581 15703 18615
rect 3893 18377 3927 18411
rect 4261 18377 4295 18411
rect 8401 18377 8435 18411
rect 8861 18309 8895 18343
rect 2789 18241 2823 18275
rect 3433 18241 3467 18275
rect 6837 18241 6871 18275
rect 7481 18241 7515 18275
rect 9965 18241 9999 18275
rect 4353 18173 4387 18207
rect 4537 18173 4571 18207
rect 2605 18037 2639 18071
rect 3249 18037 3283 18071
rect 5181 18037 5215 18071
rect 6653 18037 6687 18071
rect 7297 18037 7331 18071
rect 10149 18037 10183 18071
rect 10885 18037 10919 18071
rect 11713 18037 11747 18071
rect 12265 18037 12299 18071
rect 16773 18037 16807 18071
rect 4813 17833 4847 17867
rect 8217 17833 8251 17867
rect 2973 17629 3007 17663
rect 4353 17629 4387 17663
rect 6745 17629 6779 17663
rect 2789 17493 2823 17527
rect 4169 17493 4203 17527
rect 6561 17493 6595 17527
rect 3801 17289 3835 17323
rect 14556 17153 14590 17187
rect 14289 17085 14323 17119
rect 15669 16949 15703 16983
rect 5641 16609 5675 16643
rect 5549 16541 5583 16575
rect 5733 16541 5767 16575
rect 8953 16541 8987 16575
rect 12173 16541 12207 16575
rect 14381 16541 14415 16575
rect 9220 16473 9254 16507
rect 12440 16473 12474 16507
rect 14648 16473 14682 16507
rect 10333 16405 10367 16439
rect 13553 16405 13587 16439
rect 15761 16405 15795 16439
rect 19901 16405 19935 16439
rect 13921 16201 13955 16235
rect 19257 16201 19291 16235
rect 20085 16201 20119 16235
rect 2688 16133 2722 16167
rect 6644 16133 6678 16167
rect 9474 16133 9508 16167
rect 12808 16133 12842 16167
rect 14648 16133 14682 16167
rect 9229 16065 9263 16099
rect 19441 16065 19475 16099
rect 20453 16065 20487 16099
rect 2421 15997 2455 16031
rect 6377 15997 6411 16031
rect 12541 15997 12575 16031
rect 14381 15997 14415 16031
rect 20545 15997 20579 16031
rect 20729 15997 20763 16031
rect 15761 15929 15795 15963
rect 3801 15861 3835 15895
rect 7757 15861 7791 15895
rect 10609 15861 10643 15895
rect 10701 15657 10735 15691
rect 21741 15589 21775 15623
rect 9321 15521 9355 15555
rect 19901 15521 19935 15555
rect 21005 15521 21039 15555
rect 21097 15521 21131 15555
rect 1869 15453 1903 15487
rect 3801 15453 3835 15487
rect 4068 15453 4102 15487
rect 6193 15453 6227 15487
rect 6460 15453 6494 15487
rect 12173 15453 12207 15487
rect 14289 15453 14323 15487
rect 16129 15453 16163 15487
rect 18705 15453 18739 15487
rect 19809 15453 19843 15487
rect 2136 15385 2170 15419
rect 9588 15385 9622 15419
rect 12440 15385 12474 15419
rect 14556 15385 14590 15419
rect 16396 15385 16430 15419
rect 19717 15385 19751 15419
rect 20913 15385 20947 15419
rect 3249 15317 3283 15351
rect 5181 15317 5215 15351
rect 7573 15317 7607 15351
rect 13553 15317 13587 15351
rect 15669 15317 15703 15351
rect 17509 15317 17543 15351
rect 19349 15317 19383 15351
rect 20545 15317 20579 15351
rect 22385 15317 22419 15351
rect 18061 15113 18095 15147
rect 18705 15113 18739 15147
rect 21833 15113 21867 15147
rect 22293 15113 22327 15147
rect 6644 15045 6678 15079
rect 9588 15045 9622 15079
rect 14648 15045 14682 15079
rect 19809 15045 19843 15079
rect 2513 14977 2547 15011
rect 2780 14977 2814 15011
rect 9321 14977 9355 15011
rect 12808 14977 12842 15011
rect 18245 14977 18279 15011
rect 18889 14977 18923 15011
rect 19717 14977 19751 15011
rect 20913 14977 20947 15011
rect 22201 14977 22235 15011
rect 6377 14909 6411 14943
rect 12541 14909 12575 14943
rect 14381 14909 14415 14943
rect 17601 14909 17635 14943
rect 19901 14909 19935 14943
rect 21005 14909 21039 14943
rect 21097 14909 21131 14943
rect 22385 14909 22419 14943
rect 3893 14773 3927 14807
rect 7757 14773 7791 14807
rect 10701 14773 10735 14807
rect 13921 14773 13955 14807
rect 15761 14773 15795 14807
rect 19349 14773 19383 14807
rect 20545 14773 20579 14807
rect 23029 14773 23063 14807
rect 18521 14569 18555 14603
rect 20545 14569 20579 14603
rect 19257 14501 19291 14535
rect 21741 14501 21775 14535
rect 14105 14433 14139 14467
rect 21005 14433 21039 14467
rect 21097 14433 21131 14467
rect 22293 14433 22327 14467
rect 4629 14365 4663 14399
rect 5457 14365 5491 14399
rect 10425 14365 10459 14399
rect 14372 14365 14406 14399
rect 18705 14365 18739 14399
rect 19441 14365 19475 14399
rect 20085 14365 20119 14399
rect 5724 14297 5758 14331
rect 10158 14297 10192 14331
rect 20913 14297 20947 14331
rect 22109 14297 22143 14331
rect 4445 14229 4479 14263
rect 6837 14229 6871 14263
rect 9045 14229 9079 14263
rect 15485 14229 15519 14263
rect 19901 14229 19935 14263
rect 22201 14229 22235 14263
rect 2421 14025 2455 14059
rect 19073 14025 19107 14059
rect 19717 14025 19751 14059
rect 21005 14025 21039 14059
rect 21925 14025 21959 14059
rect 3556 13957 3590 13991
rect 14648 13957 14682 13991
rect 3801 13889 3835 13923
rect 9137 13889 9171 13923
rect 14381 13889 14415 13923
rect 19257 13889 19291 13923
rect 19901 13889 19935 13923
rect 20913 13889 20947 13923
rect 8585 13821 8619 13855
rect 21097 13821 21131 13855
rect 15761 13753 15795 13787
rect 10425 13685 10459 13719
rect 20545 13685 20579 13719
rect 19993 13481 20027 13515
rect 20729 13481 20763 13515
rect 21189 13481 21223 13515
rect 12173 13345 12207 13379
rect 20177 13277 20211 13311
rect 5273 13209 5307 13243
rect 10425 13209 10459 13243
rect 6745 13141 6779 13175
rect 10333 12937 10367 12971
rect 9220 12869 9254 12903
rect 2421 12801 2455 12835
rect 2688 12801 2722 12835
rect 7380 12801 7414 12835
rect 8953 12801 8987 12835
rect 14648 12801 14682 12835
rect 7113 12733 7147 12767
rect 14381 12733 14415 12767
rect 3801 12597 3835 12631
rect 8493 12597 8527 12631
rect 15761 12597 15795 12631
rect 19625 12393 19659 12427
rect 20637 12393 20671 12427
rect 1869 12189 1903 12223
rect 6285 12189 6319 12223
rect 10057 12189 10091 12223
rect 14289 12189 14323 12223
rect 19809 12189 19843 12223
rect 20729 12189 20763 12223
rect 2136 12121 2170 12155
rect 6552 12121 6586 12155
rect 10324 12121 10358 12155
rect 14556 12121 14590 12155
rect 3249 12053 3283 12087
rect 7665 12053 7699 12087
rect 11437 12053 11471 12087
rect 15669 12053 15703 12087
rect 18797 11849 18831 11883
rect 19809 11849 19843 11883
rect 20361 11849 20395 11883
rect 9772 11781 9806 11815
rect 2881 11713 2915 11747
rect 3148 11713 3182 11747
rect 6377 11713 6411 11747
rect 6644 11713 6678 11747
rect 14556 11713 14590 11747
rect 18981 11713 19015 11747
rect 20729 11713 20763 11747
rect 9505 11645 9539 11679
rect 14289 11645 14323 11679
rect 20821 11645 20855 11679
rect 20913 11645 20947 11679
rect 15669 11577 15703 11611
rect 4261 11509 4295 11543
rect 7757 11509 7791 11543
rect 10885 11509 10919 11543
rect 18245 11509 18279 11543
rect 5181 11305 5215 11339
rect 8401 11305 8435 11339
rect 15669 11305 15703 11339
rect 20453 11305 20487 11339
rect 3249 11237 3283 11271
rect 11437 11237 11471 11271
rect 17601 11237 17635 11271
rect 18521 11237 18555 11271
rect 10057 11169 10091 11203
rect 19901 11169 19935 11203
rect 1869 11101 1903 11135
rect 6561 11101 6595 11135
rect 7021 11101 7055 11135
rect 14289 11101 14323 11135
rect 16221 11101 16255 11135
rect 18705 11101 18739 11135
rect 19625 11101 19659 11135
rect 2136 11033 2170 11067
rect 6294 11033 6328 11067
rect 7288 11033 7322 11067
rect 10324 11033 10358 11067
rect 14556 11033 14590 11067
rect 16488 11033 16522 11067
rect 19717 11033 19751 11067
rect 19257 10965 19291 10999
rect 2881 10761 2915 10795
rect 17509 10761 17543 10795
rect 18797 10761 18831 10795
rect 19257 10761 19291 10795
rect 19993 10761 20027 10795
rect 20453 10761 20487 10795
rect 4353 10693 4387 10727
rect 14556 10693 14590 10727
rect 19165 10693 19199 10727
rect 10445 10625 10479 10659
rect 10701 10625 10735 10659
rect 17693 10625 17727 10659
rect 18337 10625 18371 10659
rect 20361 10625 20395 10659
rect 14289 10557 14323 10591
rect 19441 10557 19475 10591
rect 20545 10557 20579 10591
rect 15669 10489 15703 10523
rect 9321 10421 9355 10455
rect 18153 10421 18187 10455
rect 11713 10217 11747 10251
rect 17877 10217 17911 10251
rect 18521 10217 18555 10251
rect 19533 10217 19567 10251
rect 20729 10149 20763 10183
rect 14289 10081 14323 10115
rect 20085 10081 20119 10115
rect 21281 10081 21315 10115
rect 1869 10013 1903 10047
rect 10425 10013 10459 10047
rect 14556 10013 14590 10047
rect 18061 10013 18095 10047
rect 18705 10013 18739 10047
rect 21097 10013 21131 10047
rect 2136 9945 2170 9979
rect 19901 9945 19935 9979
rect 3249 9877 3283 9911
rect 15669 9877 15703 9911
rect 19993 9877 20027 9911
rect 21189 9877 21223 9911
rect 19165 9673 19199 9707
rect 20637 9605 20671 9639
rect 2973 9537 3007 9571
rect 8953 9537 8987 9571
rect 10977 9537 11011 9571
rect 14289 9537 14323 9571
rect 14556 9537 14590 9571
rect 18705 9537 18739 9571
rect 19533 9537 19567 9571
rect 18153 9469 18187 9503
rect 19625 9469 19659 9503
rect 19809 9469 19843 9503
rect 2789 9401 2823 9435
rect 8769 9401 8803 9435
rect 10793 9401 10827 9435
rect 15669 9401 15703 9435
rect 2421 9129 2455 9163
rect 3801 9129 3835 9163
rect 5641 9129 5675 9163
rect 9873 9129 9907 9163
rect 11437 9129 11471 9163
rect 5089 9061 5123 9095
rect 19441 9061 19475 9095
rect 4261 8993 4295 9027
rect 6101 8993 6135 9027
rect 6285 8993 6319 9027
rect 2605 8925 2639 8959
rect 3065 8925 3099 8959
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 4169 8925 4203 8959
rect 10057 8925 10091 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 10425 8925 10459 8959
rect 11621 8925 11655 8959
rect 3249 8789 3283 8823
rect 6009 8789 6043 8823
rect 2605 8585 2639 8619
rect 3065 8585 3099 8619
rect 4169 8585 4203 8619
rect 4721 8585 4755 8619
rect 6561 8585 6595 8619
rect 7849 8585 7883 8619
rect 8953 8585 8987 8619
rect 10977 8585 11011 8619
rect 11529 8585 11563 8619
rect 11713 8585 11747 8619
rect 15577 8585 15611 8619
rect 9413 8517 9447 8551
rect 10793 8517 10827 8551
rect 2697 8449 2731 8483
rect 3525 8449 3559 8483
rect 3618 8449 3652 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 3990 8449 4024 8483
rect 4905 8449 4939 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 6837 8449 6871 8483
rect 8033 8449 8067 8483
rect 8309 8449 8343 8483
rect 8493 8449 8527 8483
rect 12081 8449 12115 8483
rect 15761 8449 15795 8483
rect 17417 8449 17451 8483
rect 18061 8449 18095 8483
rect 2513 8381 2547 8415
rect 6745 8381 6779 8415
rect 6929 8381 6963 8415
rect 7021 8381 7055 8415
rect 18153 8381 18187 8415
rect 9045 8313 9079 8347
rect 10425 8313 10459 8347
rect 10793 8245 10827 8279
rect 11713 8245 11747 8279
rect 12541 8245 12575 8279
rect 18705 8245 18739 8279
rect 3801 8041 3835 8075
rect 5089 8041 5123 8075
rect 5273 8041 5307 8075
rect 5917 8041 5951 8075
rect 6837 8041 6871 8075
rect 7481 8041 7515 8075
rect 9965 8041 9999 8075
rect 11805 8041 11839 8075
rect 14105 8041 14139 8075
rect 14657 8041 14691 8075
rect 3249 7973 3283 8007
rect 10425 7973 10459 8007
rect 10149 7905 10183 7939
rect 14381 7905 14415 7939
rect 17049 7905 17083 7939
rect 17141 7905 17175 7939
rect 17969 7905 18003 7939
rect 2881 7837 2915 7871
rect 3065 7837 3099 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4445 7837 4479 7871
rect 6101 7837 6135 7871
rect 6193 7837 6227 7871
rect 6745 7837 6779 7871
rect 7573 7837 7607 7871
rect 10241 7837 10275 7871
rect 11897 7837 11931 7871
rect 14289 7837 14323 7871
rect 17233 7837 17267 7871
rect 17325 7837 17359 7871
rect 18061 7837 18095 7871
rect 5457 7769 5491 7803
rect 9965 7769 9999 7803
rect 10885 7769 10919 7803
rect 11069 7769 11103 7803
rect 14749 7769 14783 7803
rect 16405 7769 16439 7803
rect 5257 7701 5291 7735
rect 9505 7701 9539 7735
rect 11253 7701 11287 7735
rect 16865 7701 16899 7735
rect 2421 7497 2455 7531
rect 3801 7497 3835 7531
rect 5181 7497 5215 7531
rect 6653 7497 6687 7531
rect 7849 7497 7883 7531
rect 9137 7497 9171 7531
rect 10701 7497 10735 7531
rect 14933 7497 14967 7531
rect 16037 7497 16071 7531
rect 16957 7497 16991 7531
rect 20269 7497 20303 7531
rect 2789 7429 2823 7463
rect 9045 7429 9079 7463
rect 9689 7429 9723 7463
rect 15853 7429 15887 7463
rect 20085 7429 20119 7463
rect 3709 7361 3743 7395
rect 3893 7361 3927 7395
rect 4445 7361 4479 7395
rect 4537 7361 4571 7395
rect 4721 7361 4755 7395
rect 5641 7361 5675 7395
rect 8033 7361 8067 7395
rect 10517 7361 10551 7395
rect 13737 7361 13771 7395
rect 13921 7361 13955 7395
rect 14565 7361 14599 7395
rect 14749 7361 14783 7395
rect 16865 7361 16899 7395
rect 19901 7361 19935 7395
rect 20729 7361 20763 7395
rect 2881 7293 2915 7327
rect 3065 7293 3099 7327
rect 5273 7293 5307 7327
rect 5365 7293 5399 7327
rect 8217 7293 8251 7327
rect 8309 7293 8343 7327
rect 19349 7293 19383 7327
rect 15485 7225 15519 7259
rect 5549 7157 5583 7191
rect 13277 7157 13311 7191
rect 14105 7157 14139 7191
rect 14565 7157 14599 7191
rect 15853 7157 15887 7191
rect 20913 7157 20947 7191
rect 3065 6953 3099 6987
rect 6009 6953 6043 6987
rect 14105 6953 14139 6987
rect 14473 6953 14507 6987
rect 15025 6953 15059 6987
rect 15577 6953 15611 6987
rect 16129 6953 16163 6987
rect 19809 6953 19843 6987
rect 6561 6885 6595 6919
rect 8953 6817 8987 6851
rect 9321 6817 9355 6851
rect 13001 6817 13035 6851
rect 15209 6817 15243 6851
rect 16221 6817 16255 6851
rect 19441 6817 19475 6851
rect 20453 6817 20487 6851
rect 21005 6817 21039 6851
rect 2789 6749 2823 6783
rect 5917 6749 5951 6783
rect 6101 6749 6135 6783
rect 6745 6749 6779 6783
rect 9137 6749 9171 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 14105 6749 14139 6783
rect 14289 6749 14323 6783
rect 14933 6749 14967 6783
rect 15393 6749 15427 6783
rect 16129 6749 16163 6783
rect 16957 6749 16991 6783
rect 17693 6749 17727 6783
rect 17877 6749 17911 6783
rect 21189 6749 21223 6783
rect 21373 6749 21407 6783
rect 21465 6749 21499 6783
rect 6929 6681 6963 6715
rect 7113 6681 7147 6715
rect 12817 6681 12851 6715
rect 17785 6681 17819 6715
rect 19809 6681 19843 6715
rect 3249 6613 3283 6647
rect 3801 6613 3835 6647
rect 6837 6613 6871 6647
rect 12357 6613 12391 6647
rect 12725 6613 12759 6647
rect 16497 6613 16531 6647
rect 17141 6613 17175 6647
rect 18613 6613 18647 6647
rect 19993 6613 20027 6647
rect 2697 6409 2731 6443
rect 8217 6409 8251 6443
rect 9781 6409 9815 6443
rect 10977 6409 11011 6443
rect 18981 6409 19015 6443
rect 19349 6409 19383 6443
rect 20453 6409 20487 6443
rect 22385 6409 22419 6443
rect 10241 6341 10275 6375
rect 11897 6341 11931 6375
rect 15025 6341 15059 6375
rect 17233 6341 17267 6375
rect 18337 6341 18371 6375
rect 20729 6341 20763 6375
rect 20821 6341 20855 6375
rect 22753 6341 22787 6375
rect 2881 6273 2915 6307
rect 3157 6273 3191 6307
rect 8677 6273 8711 6307
rect 8861 6273 8895 6307
rect 9413 6273 9447 6307
rect 9597 6273 9631 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 12015 6273 12049 6307
rect 13369 6273 13403 6307
rect 13737 6273 13771 6307
rect 14565 6273 14599 6307
rect 14933 6273 14967 6307
rect 18245 6273 18279 6307
rect 18429 6273 18463 6307
rect 18889 6273 18923 6307
rect 19165 6273 19199 6307
rect 19993 6273 20027 6307
rect 20591 6273 20625 6307
rect 20949 6273 20983 6307
rect 21097 6273 21131 6307
rect 22569 6273 22603 6307
rect 22845 6273 22879 6307
rect 2973 6205 3007 6239
rect 8769 6205 8803 6239
rect 12173 6205 12207 6239
rect 13277 6205 13311 6239
rect 14657 6205 14691 6239
rect 19901 6205 19935 6239
rect 3065 6137 3099 6171
rect 4261 6137 4295 6171
rect 13921 6137 13955 6171
rect 3801 6069 3835 6103
rect 9597 6069 9631 6103
rect 11529 6069 11563 6103
rect 13737 6069 13771 6103
rect 14749 6069 14783 6103
rect 17325 6069 17359 6103
rect 23397 6069 23431 6103
rect 7389 5865 7423 5899
rect 9045 5865 9079 5899
rect 12633 5865 12667 5899
rect 14381 5865 14415 5899
rect 19717 5865 19751 5899
rect 20453 5865 20487 5899
rect 10425 5797 10459 5831
rect 10517 5729 10551 5763
rect 12357 5729 12391 5763
rect 12541 5729 12575 5763
rect 7665 5661 7699 5695
rect 7757 5661 7791 5695
rect 7849 5661 7883 5695
rect 8033 5661 8067 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 10241 5661 10275 5695
rect 11161 5661 11195 5695
rect 11437 5661 11471 5695
rect 11621 5661 11655 5695
rect 12633 5661 12667 5695
rect 19257 5661 19291 5695
rect 19533 5661 19567 5695
rect 20269 5661 20303 5695
rect 10977 5593 11011 5627
rect 10057 5525 10091 5559
rect 19349 5525 19383 5559
rect 6377 5321 6411 5355
rect 7297 5321 7331 5355
rect 8309 5321 8343 5355
rect 18245 5321 18279 5355
rect 21833 5321 21867 5355
rect 17509 5253 17543 5287
rect 6561 5185 6595 5219
rect 7573 5185 7607 5219
rect 7757 5185 7791 5219
rect 19901 5185 19935 5219
rect 22017 5185 22051 5219
rect 22201 5185 22235 5219
rect 22293 5185 22327 5219
rect 7481 5117 7515 5151
rect 7665 5117 7699 5151
rect 20085 5049 20119 5083
rect 9965 4981 9999 5015
rect 16773 4981 16807 5015
rect 6101 4777 6135 4811
rect 9597 4777 9631 4811
rect 10149 4777 10183 4811
rect 17785 4777 17819 4811
rect 20177 4777 20211 4811
rect 21833 4777 21867 4811
rect 23489 4777 23523 4811
rect 24409 4777 24443 4811
rect 18705 4709 18739 4743
rect 7941 4641 7975 4675
rect 6653 4573 6687 4607
rect 6837 4573 6871 4607
rect 7021 4573 7055 4607
rect 7849 4573 7883 4607
rect 8033 4573 8067 4607
rect 10333 4573 10367 4607
rect 10517 4573 10551 4607
rect 10609 4573 10643 4607
rect 15393 4573 15427 4607
rect 17325 4573 17359 4607
rect 17601 4573 17635 4607
rect 18245 4573 18279 4607
rect 18337 4573 18371 4607
rect 18521 4573 18555 4607
rect 19717 4573 19751 4607
rect 19809 4573 19843 4607
rect 19993 4573 20027 4607
rect 21373 4573 21407 4607
rect 21649 4573 21683 4607
rect 24593 4573 24627 4607
rect 24869 4573 24903 4607
rect 6929 4505 6963 4539
rect 11161 4505 11195 4539
rect 7205 4437 7239 4471
rect 11713 4437 11747 4471
rect 15853 4437 15887 4471
rect 16773 4437 16807 4471
rect 17417 4437 17451 4471
rect 21465 4437 21499 4471
rect 22937 4437 22971 4471
rect 24777 4437 24811 4471
rect 6745 4233 6779 4267
rect 12173 4233 12207 4267
rect 22109 4233 22143 4267
rect 17601 4165 17635 4199
rect 18797 4165 18831 4199
rect 23489 4165 23523 4199
rect 6929 4097 6963 4131
rect 9321 4097 9355 4131
rect 10057 4097 10091 4131
rect 10149 4097 10183 4131
rect 10241 4097 10275 4131
rect 10425 4097 10459 4131
rect 12014 4097 12048 4131
rect 15117 4097 15151 4131
rect 15301 4097 15335 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 17509 4097 17543 4131
rect 17693 4097 17727 4131
rect 17877 4097 17911 4131
rect 18521 4097 18555 4131
rect 18705 4097 18739 4131
rect 18889 4097 18923 4131
rect 19625 4097 19659 4131
rect 22293 4097 22327 4131
rect 22385 4097 22419 4131
rect 22477 4097 22511 4131
rect 22661 4097 22695 4131
rect 23259 4097 23293 4131
rect 23373 4097 23407 4131
rect 23673 4097 23707 4131
rect 24133 4097 24167 4131
rect 24317 4097 24351 4131
rect 24501 4097 24535 4131
rect 24593 4097 24627 4131
rect 25605 4097 25639 4131
rect 26249 4097 26283 4131
rect 7113 4029 7147 4063
rect 9781 4029 9815 4063
rect 11529 4029 11563 4063
rect 11805 4029 11839 4063
rect 11897 4029 11931 4063
rect 12725 4029 12759 4063
rect 8769 3961 8803 3995
rect 13185 3961 13219 3995
rect 14657 3961 14691 3995
rect 15393 3961 15427 3995
rect 15485 3961 15519 3995
rect 16865 3961 16899 3995
rect 17325 3961 17359 3995
rect 19073 3961 19107 3995
rect 23121 3961 23155 3995
rect 5365 3893 5399 3927
rect 8217 3893 8251 3927
rect 10977 3893 11011 3927
rect 14105 3893 14139 3927
rect 20085 3893 20119 3927
rect 25053 3893 25087 3927
rect 9505 3689 9539 3723
rect 11989 3689 12023 3723
rect 15393 3689 15427 3723
rect 15577 3689 15611 3723
rect 16129 3689 16163 3723
rect 16497 3689 16531 3723
rect 17141 3689 17175 3723
rect 18705 3689 18739 3723
rect 19993 3689 20027 3723
rect 21005 3689 21039 3723
rect 21557 3689 21591 3723
rect 23581 3689 23615 3723
rect 24961 3689 24995 3723
rect 26525 3689 26559 3723
rect 27077 3689 27111 3723
rect 27629 3689 27663 3723
rect 36645 3689 36679 3723
rect 19349 3621 19383 3655
rect 22569 3621 22603 3655
rect 7849 3553 7883 3587
rect 10977 3553 11011 3587
rect 11529 3553 11563 3587
rect 15301 3553 15335 3587
rect 16497 3553 16531 3587
rect 25421 3553 25455 3587
rect 6193 3485 6227 3519
rect 10425 3485 10459 3519
rect 10701 3485 10735 3519
rect 11253 3485 11287 3519
rect 15117 3485 15151 3519
rect 15393 3485 15427 3519
rect 16313 3485 16347 3519
rect 16589 3485 16623 3519
rect 17325 3485 17359 3519
rect 17509 3485 17543 3519
rect 17693 3485 17727 3519
rect 18153 3485 18187 3519
rect 18337 3485 18371 3519
rect 18521 3485 18555 3519
rect 20177 3485 20211 3519
rect 20545 3485 20579 3519
rect 21741 3485 21775 3519
rect 22089 3485 22123 3519
rect 22753 3485 22787 3519
rect 22845 3485 22879 3519
rect 23121 3485 23155 3519
rect 24409 3485 24443 3519
rect 24777 3485 24811 3519
rect 36829 3485 36863 3519
rect 37289 3485 37323 3519
rect 7297 3417 7331 3451
rect 8401 3417 8435 3451
rect 17417 3417 17451 3451
rect 18429 3417 18463 3451
rect 20269 3417 20303 3451
rect 20361 3417 20395 3451
rect 21833 3417 21867 3451
rect 21925 3417 21959 3451
rect 22937 3417 22971 3451
rect 24593 3417 24627 3451
rect 24685 3417 24719 3451
rect 25973 3417 26007 3451
rect 3985 3349 4019 3383
rect 4537 3349 4571 3383
rect 5089 3349 5123 3383
rect 5641 3349 5675 3383
rect 6745 3349 6779 3383
rect 12817 3349 12851 3383
rect 13369 3349 13403 3383
rect 14657 3349 14691 3383
rect 28181 3349 28215 3383
rect 28733 3349 28767 3383
rect 29561 3349 29595 3383
rect 30481 3349 30515 3383
rect 31125 3349 31159 3383
rect 33241 3349 33275 3383
rect 33701 3349 33735 3383
rect 34713 3349 34747 3383
rect 35449 3349 35483 3383
rect 36001 3349 36035 3383
rect 38025 3349 38059 3383
rect 3157 3145 3191 3179
rect 4721 3145 4755 3179
rect 7021 3145 7055 3179
rect 10609 3145 10643 3179
rect 13645 3145 13679 3179
rect 14381 3145 14415 3179
rect 15209 3145 15243 3179
rect 16129 3145 16163 3179
rect 16865 3145 16899 3179
rect 17785 3145 17819 3179
rect 18245 3145 18279 3179
rect 19809 3145 19843 3179
rect 21833 3145 21867 3179
rect 22845 3145 22879 3179
rect 24409 3145 24443 3179
rect 28365 3145 28399 3179
rect 29009 3145 29043 3179
rect 31217 3145 31251 3179
rect 33333 3145 33367 3179
rect 34437 3145 34471 3179
rect 36093 3145 36127 3179
rect 13001 3077 13035 3111
rect 17417 3077 17451 3111
rect 19441 3077 19475 3111
rect 23121 3077 23155 3111
rect 24041 3077 24075 3111
rect 26341 3077 26375 3111
rect 2513 3009 2547 3043
rect 3065 3009 3099 3043
rect 3893 3009 3927 3043
rect 4537 3009 4571 3043
rect 5181 3009 5215 3043
rect 6837 3009 6871 3043
rect 8493 3009 8527 3043
rect 9597 3009 9631 3043
rect 10609 3009 10643 3043
rect 10793 3009 10827 3043
rect 11805 3009 11839 3043
rect 13461 3009 13495 3043
rect 14197 3009 14231 3043
rect 14841 3009 14875 3043
rect 15025 3009 15059 3043
rect 15945 3009 15979 3043
rect 16681 3009 16715 3043
rect 17325 3009 17359 3043
rect 17601 3009 17635 3043
rect 18429 3009 18463 3043
rect 18521 3009 18555 3043
rect 18613 3009 18647 3043
rect 18797 3009 18831 3043
rect 19257 3009 19291 3043
rect 19533 3009 19567 3043
rect 19625 3009 19659 3043
rect 20545 3009 20579 3043
rect 21005 3009 21039 3043
rect 22017 3009 22051 3043
rect 22109 3009 22143 3043
rect 22201 3009 22235 3043
rect 22385 3009 22419 3043
rect 23005 3009 23039 3043
rect 23213 3009 23247 3043
rect 23397 3009 23431 3043
rect 23857 3009 23891 3043
rect 24133 3009 24167 3043
rect 24225 3009 24259 3043
rect 25145 3009 25179 3043
rect 25605 3009 25639 3043
rect 26985 3009 27019 3043
rect 27905 3009 27939 3043
rect 28549 3009 28583 3043
rect 30757 3009 30791 3043
rect 31401 3009 31435 3043
rect 33517 3009 33551 3043
rect 34621 3009 34655 3043
rect 35081 3009 35115 3043
rect 36277 3009 36311 3043
rect 37565 3009 37599 3043
rect 38025 3009 38059 3043
rect 4077 2873 4111 2907
rect 5365 2873 5399 2907
rect 8677 2873 8711 2907
rect 11989 2873 12023 2907
rect 20361 2873 20395 2907
rect 27169 2873 27203 2907
rect 29561 2873 29595 2907
rect 30573 2873 30607 2907
rect 37381 2873 37415 2907
rect 8033 2805 8067 2839
rect 9781 2805 9815 2839
rect 14933 2805 14967 2839
rect 24961 2805 24995 2839
rect 25789 2805 25823 2839
rect 27721 2805 27755 2839
rect 32137 2805 32171 2839
rect 32689 2805 32723 2839
rect 9689 2601 9723 2635
rect 19441 2601 19475 2635
rect 25237 2601 25271 2635
rect 28457 2601 28491 2635
rect 35357 2601 35391 2635
rect 5825 2533 5859 2567
rect 10333 2533 10367 2567
rect 12265 2533 12299 2567
rect 14749 2533 14783 2567
rect 15393 2533 15427 2567
rect 22661 2533 22695 2567
rect 25973 2533 26007 2567
rect 27813 2533 27847 2567
rect 30849 2533 30883 2567
rect 2697 2465 2731 2499
rect 15853 2465 15887 2499
rect 38117 2465 38151 2499
rect 1961 2397 1995 2431
rect 2421 2397 2455 2431
rect 4077 2397 4111 2431
rect 4997 2397 5031 2431
rect 5641 2397 5675 2431
rect 6929 2397 6963 2431
rect 7573 2397 7607 2431
rect 8217 2397 8251 2431
rect 9505 2397 9539 2431
rect 10149 2397 10183 2431
rect 10793 2397 10827 2431
rect 12081 2397 12115 2431
rect 12725 2397 12759 2431
rect 13369 2397 13403 2431
rect 14565 2397 14599 2431
rect 15209 2397 15243 2431
rect 16957 2397 16991 2431
rect 17693 2397 17727 2431
rect 18429 2397 18463 2431
rect 20177 2397 20211 2431
rect 20637 2397 20671 2431
rect 21833 2397 21867 2431
rect 22845 2397 22879 2431
rect 23581 2397 23615 2431
rect 24685 2397 24719 2431
rect 25421 2397 25455 2431
rect 26157 2397 26191 2431
rect 27261 2397 27295 2431
rect 27997 2397 28031 2431
rect 28641 2397 28675 2431
rect 29745 2397 29779 2431
rect 30389 2397 30423 2431
rect 31033 2397 31067 2431
rect 32321 2397 32355 2431
rect 32965 2397 32999 2431
rect 33609 2397 33643 2431
rect 34897 2397 34931 2431
rect 35541 2397 35575 2431
rect 36185 2397 36219 2431
rect 37841 2397 37875 2431
rect 6469 2329 6503 2363
rect 9045 2329 9079 2363
rect 11621 2329 11655 2363
rect 16037 2329 16071 2363
rect 31493 2329 31527 2363
rect 34069 2329 34103 2363
rect 36645 2329 36679 2363
rect 3893 2261 3927 2295
rect 5181 2261 5215 2295
rect 7113 2261 7147 2295
rect 7757 2261 7791 2295
rect 8401 2261 8435 2295
rect 10977 2261 11011 2295
rect 12909 2261 12943 2295
rect 13553 2261 13587 2295
rect 17141 2261 17175 2295
rect 17877 2261 17911 2295
rect 18613 2261 18647 2295
rect 19993 2261 20027 2295
rect 20821 2261 20855 2295
rect 22017 2261 22051 2295
rect 23397 2261 23431 2295
rect 24501 2261 24535 2295
rect 27077 2261 27111 2295
rect 29561 2261 29595 2295
rect 30205 2261 30239 2295
rect 32137 2261 32171 2295
rect 32781 2261 32815 2295
rect 33425 2261 33459 2295
rect 34713 2261 34747 2295
rect 36001 2261 36035 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 8386 37448 8392 37460
rect 8347 37420 8392 37448
rect 8386 37408 8392 37420
rect 8444 37408 8450 37460
rect 16114 37448 16120 37460
rect 16075 37420 16120 37448
rect 16114 37408 16120 37420
rect 16172 37448 16178 37460
rect 16172 37420 16574 37448
rect 16172 37408 16178 37420
rect 658 37204 664 37256
rect 716 37244 722 37256
rect 1302 37244 1308 37256
rect 716 37216 1308 37244
rect 716 37204 722 37216
rect 1302 37204 1308 37216
rect 1360 37244 1366 37256
rect 1857 37247 1915 37253
rect 1857 37244 1869 37247
rect 1360 37216 1869 37244
rect 1360 37204 1366 37216
rect 1857 37213 1869 37216
rect 1903 37213 1915 37247
rect 1857 37207 1915 37213
rect 2866 37204 2872 37256
rect 2924 37244 2930 37256
rect 2961 37247 3019 37253
rect 2961 37244 2973 37247
rect 2924 37216 2973 37244
rect 2924 37204 2930 37216
rect 2961 37213 2973 37216
rect 3007 37213 3019 37247
rect 2961 37207 3019 37213
rect 3970 37204 3976 37256
rect 4028 37244 4034 37256
rect 4065 37247 4123 37253
rect 4065 37244 4077 37247
rect 4028 37216 4077 37244
rect 4028 37204 4034 37216
rect 4065 37213 4077 37216
rect 4111 37213 4123 37247
rect 4065 37207 4123 37213
rect 5074 37204 5080 37256
rect 5132 37244 5138 37256
rect 5353 37247 5411 37253
rect 5353 37244 5365 37247
rect 5132 37216 5365 37244
rect 5132 37204 5138 37216
rect 5353 37213 5365 37216
rect 5399 37213 5411 37247
rect 5353 37207 5411 37213
rect 6178 37204 6184 37256
rect 6236 37244 6242 37256
rect 6549 37247 6607 37253
rect 6549 37244 6561 37247
rect 6236 37216 6561 37244
rect 6236 37204 6242 37216
rect 6549 37213 6561 37216
rect 6595 37213 6607 37247
rect 6549 37207 6607 37213
rect 7282 37204 7288 37256
rect 7340 37244 7346 37256
rect 7561 37247 7619 37253
rect 7561 37244 7573 37247
rect 7340 37216 7573 37244
rect 7340 37204 7346 37216
rect 7561 37213 7573 37216
rect 7607 37213 7619 37247
rect 7561 37207 7619 37213
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 9125 37247 9183 37253
rect 9125 37244 9137 37247
rect 8444 37216 9137 37244
rect 8444 37204 8450 37216
rect 9125 37213 9137 37216
rect 9171 37213 9183 37247
rect 9125 37207 9183 37213
rect 9490 37204 9496 37256
rect 9548 37244 9554 37256
rect 9769 37247 9827 37253
rect 9769 37244 9781 37247
rect 9548 37216 9781 37244
rect 9548 37204 9554 37216
rect 9769 37213 9781 37216
rect 9815 37213 9827 37247
rect 9769 37207 9827 37213
rect 10594 37204 10600 37256
rect 10652 37244 10658 37256
rect 10873 37247 10931 37253
rect 10873 37244 10885 37247
rect 10652 37216 10885 37244
rect 10652 37204 10658 37216
rect 10873 37213 10885 37216
rect 10919 37213 10931 37247
rect 10873 37207 10931 37213
rect 11698 37204 11704 37256
rect 11756 37244 11762 37256
rect 11977 37247 12035 37253
rect 11977 37244 11989 37247
rect 11756 37216 11989 37244
rect 11756 37204 11762 37216
rect 11977 37213 11989 37216
rect 12023 37213 12035 37247
rect 11977 37207 12035 37213
rect 12802 37204 12808 37256
rect 12860 37244 12866 37256
rect 13081 37247 13139 37253
rect 13081 37244 13093 37247
rect 12860 37216 13093 37244
rect 12860 37204 12866 37216
rect 13081 37213 13093 37216
rect 13127 37213 13139 37247
rect 13081 37207 13139 37213
rect 13906 37204 13912 37256
rect 13964 37244 13970 37256
rect 14277 37247 14335 37253
rect 14277 37244 14289 37247
rect 13964 37216 14289 37244
rect 13964 37204 13970 37216
rect 14277 37213 14289 37216
rect 14323 37213 14335 37247
rect 14277 37207 14335 37213
rect 15010 37204 15016 37256
rect 15068 37244 15074 37256
rect 15289 37247 15347 37253
rect 15289 37244 15301 37247
rect 15068 37216 15301 37244
rect 15068 37204 15074 37216
rect 15289 37213 15301 37216
rect 15335 37213 15347 37247
rect 16546 37244 16574 37420
rect 31478 37312 31484 37324
rect 31439 37284 31484 37312
rect 31478 37272 31484 37284
rect 31536 37312 31542 37324
rect 31536 37284 32168 37312
rect 31536 37272 31542 37284
rect 16853 37247 16911 37253
rect 16853 37244 16865 37247
rect 16546 37216 16865 37244
rect 15289 37207 15347 37213
rect 16853 37213 16865 37216
rect 16899 37213 16911 37247
rect 16853 37207 16911 37213
rect 17218 37204 17224 37256
rect 17276 37244 17282 37256
rect 17497 37247 17555 37253
rect 17497 37244 17509 37247
rect 17276 37216 17509 37244
rect 17276 37204 17282 37216
rect 17497 37213 17509 37216
rect 17543 37213 17555 37247
rect 17497 37207 17555 37213
rect 18322 37204 18328 37256
rect 18380 37244 18386 37256
rect 18601 37247 18659 37253
rect 18601 37244 18613 37247
rect 18380 37216 18613 37244
rect 18380 37204 18386 37216
rect 18601 37213 18613 37216
rect 18647 37213 18659 37247
rect 18601 37207 18659 37213
rect 19426 37204 19432 37256
rect 19484 37244 19490 37256
rect 19705 37247 19763 37253
rect 19705 37244 19717 37247
rect 19484 37216 19717 37244
rect 19484 37204 19490 37216
rect 19705 37213 19717 37216
rect 19751 37213 19763 37247
rect 19705 37207 19763 37213
rect 20530 37204 20536 37256
rect 20588 37244 20594 37256
rect 20809 37247 20867 37253
rect 20809 37244 20821 37247
rect 20588 37216 20821 37244
rect 20588 37204 20594 37216
rect 20809 37213 20821 37216
rect 20855 37213 20867 37247
rect 21818 37244 21824 37256
rect 21779 37216 21824 37244
rect 20809 37207 20867 37213
rect 21818 37204 21824 37216
rect 21876 37204 21882 37256
rect 23014 37204 23020 37256
rect 23072 37244 23078 37256
rect 23109 37247 23167 37253
rect 23109 37244 23121 37247
rect 23072 37216 23121 37244
rect 23072 37204 23078 37216
rect 23109 37213 23121 37216
rect 23155 37213 23167 37247
rect 23109 37207 23167 37213
rect 23845 37247 23903 37253
rect 23845 37213 23857 37247
rect 23891 37244 23903 37247
rect 24394 37244 24400 37256
rect 23891 37216 24400 37244
rect 23891 37213 23903 37216
rect 23845 37207 23903 37213
rect 24394 37204 24400 37216
rect 24452 37204 24458 37256
rect 25130 37244 25136 37256
rect 25091 37216 25136 37244
rect 25130 37204 25136 37216
rect 25188 37204 25194 37256
rect 26145 37247 26203 37253
rect 26145 37213 26157 37247
rect 26191 37213 26203 37247
rect 27246 37244 27252 37256
rect 27207 37216 27252 37244
rect 26145 37207 26203 37213
rect 4614 37136 4620 37188
rect 4672 37176 4678 37188
rect 4672 37148 5212 37176
rect 4672 37136 4678 37148
rect 1946 37108 1952 37120
rect 1907 37080 1952 37108
rect 1946 37068 1952 37080
rect 2004 37068 2010 37120
rect 3142 37108 3148 37120
rect 3103 37080 3148 37108
rect 3142 37068 3148 37080
rect 3200 37068 3206 37120
rect 4249 37111 4307 37117
rect 4249 37077 4261 37111
rect 4295 37108 4307 37111
rect 4706 37108 4712 37120
rect 4295 37080 4712 37108
rect 4295 37077 4307 37080
rect 4249 37071 4307 37077
rect 4706 37068 4712 37080
rect 4764 37068 4770 37120
rect 5184 37117 5212 37148
rect 10318 37136 10324 37188
rect 10376 37176 10382 37188
rect 10376 37148 12940 37176
rect 10376 37136 10382 37148
rect 5169 37111 5227 37117
rect 5169 37077 5181 37111
rect 5215 37077 5227 37111
rect 6362 37108 6368 37120
rect 6323 37080 6368 37108
rect 5169 37071 5227 37077
rect 6362 37068 6368 37080
rect 6420 37068 6426 37120
rect 7374 37108 7380 37120
rect 7335 37080 7380 37108
rect 7374 37068 7380 37080
rect 7432 37068 7438 37120
rect 8938 37108 8944 37120
rect 8899 37080 8944 37108
rect 8938 37068 8944 37080
rect 8996 37068 9002 37120
rect 9582 37108 9588 37120
rect 9543 37080 9588 37108
rect 9582 37068 9588 37080
rect 9640 37068 9646 37120
rect 10686 37108 10692 37120
rect 10647 37080 10692 37108
rect 10686 37068 10692 37080
rect 10744 37068 10750 37120
rect 11514 37068 11520 37120
rect 11572 37108 11578 37120
rect 12912 37117 12940 37148
rect 15838 37136 15844 37188
rect 15896 37176 15902 37188
rect 15896 37148 17356 37176
rect 15896 37136 15902 37148
rect 11793 37111 11851 37117
rect 11793 37108 11805 37111
rect 11572 37080 11805 37108
rect 11572 37068 11578 37080
rect 11793 37077 11805 37080
rect 11839 37077 11851 37111
rect 11793 37071 11851 37077
rect 12897 37111 12955 37117
rect 12897 37077 12909 37111
rect 12943 37077 12955 37111
rect 14090 37108 14096 37120
rect 14051 37080 14096 37108
rect 12897 37071 12955 37077
rect 14090 37068 14096 37080
rect 14148 37068 14154 37120
rect 15102 37108 15108 37120
rect 15063 37080 15108 37108
rect 15102 37068 15108 37080
rect 15160 37068 15166 37120
rect 16669 37111 16727 37117
rect 16669 37077 16681 37111
rect 16715 37108 16727 37111
rect 16758 37108 16764 37120
rect 16715 37080 16764 37108
rect 16715 37077 16727 37080
rect 16669 37071 16727 37077
rect 16758 37068 16764 37080
rect 16816 37068 16822 37120
rect 17328 37117 17356 37148
rect 26160 37120 26188 37207
rect 27246 37204 27252 37216
rect 27304 37204 27310 37256
rect 28166 37204 28172 37256
rect 28224 37244 28230 37256
rect 28353 37247 28411 37253
rect 28353 37244 28365 37247
rect 28224 37216 28365 37244
rect 28224 37204 28230 37216
rect 28353 37213 28365 37216
rect 28399 37213 28411 37247
rect 28353 37207 28411 37213
rect 29362 37204 29368 37256
rect 29420 37244 29426 37256
rect 29549 37247 29607 37253
rect 29549 37244 29561 37247
rect 29420 37216 29561 37244
rect 29420 37204 29426 37216
rect 29549 37213 29561 37216
rect 29595 37213 29607 37247
rect 29549 37207 29607 37213
rect 30374 37204 30380 37256
rect 30432 37244 30438 37256
rect 32140 37253 32168 37284
rect 30561 37247 30619 37253
rect 30561 37244 30573 37247
rect 30432 37216 30573 37244
rect 30432 37204 30438 37216
rect 30561 37213 30573 37216
rect 30607 37213 30619 37247
rect 30561 37207 30619 37213
rect 32125 37247 32183 37253
rect 32125 37213 32137 37247
rect 32171 37213 32183 37247
rect 32858 37244 32864 37256
rect 32819 37216 32864 37244
rect 32125 37207 32183 37213
rect 32858 37204 32864 37216
rect 32916 37204 32922 37256
rect 33870 37244 33876 37256
rect 33831 37216 33876 37244
rect 33870 37204 33876 37216
rect 33928 37204 33934 37256
rect 34790 37204 34796 37256
rect 34848 37244 34854 37256
rect 34977 37247 35035 37253
rect 34977 37244 34989 37247
rect 34848 37216 34989 37244
rect 34848 37204 34854 37216
rect 34977 37213 34989 37216
rect 35023 37213 35035 37247
rect 34977 37207 35035 37213
rect 35894 37204 35900 37256
rect 35952 37244 35958 37256
rect 36081 37247 36139 37253
rect 36081 37244 36093 37247
rect 35952 37216 36093 37244
rect 35952 37204 35958 37216
rect 36081 37213 36093 37216
rect 36127 37213 36139 37247
rect 36081 37207 36139 37213
rect 37277 37247 37335 37253
rect 37277 37213 37289 37247
rect 37323 37244 37335 37247
rect 37366 37244 37372 37256
rect 37323 37216 37372 37244
rect 37323 37213 37335 37216
rect 37277 37207 37335 37213
rect 37366 37204 37372 37216
rect 37424 37204 37430 37256
rect 17313 37111 17371 37117
rect 17313 37077 17325 37111
rect 17359 37077 17371 37111
rect 18414 37108 18420 37120
rect 18375 37080 18420 37108
rect 17313 37071 17371 37077
rect 18414 37068 18420 37080
rect 18472 37068 18478 37120
rect 19426 37068 19432 37120
rect 19484 37108 19490 37120
rect 19521 37111 19579 37117
rect 19521 37108 19533 37111
rect 19484 37080 19533 37108
rect 19484 37068 19490 37080
rect 19521 37077 19533 37080
rect 19567 37077 19579 37111
rect 20622 37108 20628 37120
rect 20583 37080 20628 37108
rect 19521 37071 19579 37077
rect 20622 37068 20628 37080
rect 20680 37068 20686 37120
rect 21634 37068 21640 37120
rect 21692 37108 21698 37120
rect 22005 37111 22063 37117
rect 22005 37108 22017 37111
rect 21692 37080 22017 37108
rect 21692 37068 21698 37080
rect 22005 37077 22017 37080
rect 22051 37077 22063 37111
rect 22005 37071 22063 37077
rect 22738 37068 22744 37120
rect 22796 37108 22802 37120
rect 22925 37111 22983 37117
rect 22925 37108 22937 37111
rect 22796 37080 22937 37108
rect 22796 37068 22802 37080
rect 22925 37077 22937 37080
rect 22971 37077 22983 37111
rect 22925 37071 22983 37077
rect 23842 37068 23848 37120
rect 23900 37108 23906 37120
rect 24581 37111 24639 37117
rect 24581 37108 24593 37111
rect 23900 37080 24593 37108
rect 23900 37068 23906 37080
rect 24581 37077 24593 37080
rect 24627 37077 24639 37111
rect 24581 37071 24639 37077
rect 24946 37068 24952 37120
rect 25004 37108 25010 37120
rect 25317 37111 25375 37117
rect 25317 37108 25329 37111
rect 25004 37080 25329 37108
rect 25004 37068 25010 37080
rect 25317 37077 25329 37080
rect 25363 37077 25375 37111
rect 25317 37071 25375 37077
rect 26142 37068 26148 37120
rect 26200 37068 26206 37120
rect 26234 37068 26240 37120
rect 26292 37108 26298 37120
rect 26329 37111 26387 37117
rect 26329 37108 26341 37111
rect 26292 37080 26341 37108
rect 26292 37068 26298 37080
rect 26329 37077 26341 37080
rect 26375 37077 26387 37111
rect 26329 37071 26387 37077
rect 27154 37068 27160 37120
rect 27212 37108 27218 37120
rect 27433 37111 27491 37117
rect 27433 37108 27445 37111
rect 27212 37080 27445 37108
rect 27212 37068 27218 37080
rect 27433 37077 27445 37080
rect 27479 37077 27491 37111
rect 27433 37071 27491 37077
rect 28258 37068 28264 37120
rect 28316 37108 28322 37120
rect 28537 37111 28595 37117
rect 28537 37108 28549 37111
rect 28316 37080 28549 37108
rect 28316 37068 28322 37080
rect 28537 37077 28549 37080
rect 28583 37077 28595 37111
rect 28537 37071 28595 37077
rect 29454 37068 29460 37120
rect 29512 37108 29518 37120
rect 29733 37111 29791 37117
rect 29733 37108 29745 37111
rect 29512 37080 29745 37108
rect 29512 37068 29518 37080
rect 29733 37077 29745 37080
rect 29779 37077 29791 37111
rect 29733 37071 29791 37077
rect 30466 37068 30472 37120
rect 30524 37108 30530 37120
rect 30745 37111 30803 37117
rect 30745 37108 30757 37111
rect 30524 37080 30757 37108
rect 30524 37068 30530 37080
rect 30745 37077 30757 37080
rect 30791 37077 30803 37111
rect 30745 37071 30803 37077
rect 31754 37068 31760 37120
rect 31812 37108 31818 37120
rect 32309 37111 32367 37117
rect 32309 37108 32321 37111
rect 31812 37080 32321 37108
rect 31812 37068 31818 37080
rect 32309 37077 32321 37080
rect 32355 37077 32367 37111
rect 32309 37071 32367 37077
rect 32674 37068 32680 37120
rect 32732 37108 32738 37120
rect 33045 37111 33103 37117
rect 33045 37108 33057 37111
rect 32732 37080 33057 37108
rect 32732 37068 32738 37080
rect 33045 37077 33057 37080
rect 33091 37077 33103 37111
rect 33045 37071 33103 37077
rect 33778 37068 33784 37120
rect 33836 37108 33842 37120
rect 34057 37111 34115 37117
rect 34057 37108 34069 37111
rect 33836 37080 34069 37108
rect 33836 37068 33842 37080
rect 34057 37077 34069 37080
rect 34103 37077 34115 37111
rect 34057 37071 34115 37077
rect 34882 37068 34888 37120
rect 34940 37108 34946 37120
rect 35161 37111 35219 37117
rect 35161 37108 35173 37111
rect 34940 37080 35173 37108
rect 34940 37068 34946 37080
rect 35161 37077 35173 37080
rect 35207 37077 35219 37111
rect 35161 37071 35219 37077
rect 35986 37068 35992 37120
rect 36044 37108 36050 37120
rect 36265 37111 36323 37117
rect 36265 37108 36277 37111
rect 36044 37080 36277 37108
rect 36044 37068 36050 37080
rect 36265 37077 36277 37080
rect 36311 37077 36323 37111
rect 36265 37071 36323 37077
rect 37090 37068 37096 37120
rect 37148 37108 37154 37120
rect 37461 37111 37519 37117
rect 37461 37108 37473 37111
rect 37148 37080 37473 37108
rect 37148 37068 37154 37080
rect 37461 37077 37473 37080
rect 37507 37077 37519 37111
rect 38010 37108 38016 37120
rect 37971 37080 38016 37108
rect 37461 37071 37519 37077
rect 38010 37068 38016 37080
rect 38068 37068 38074 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1762 36864 1768 36916
rect 1820 36904 1826 36916
rect 1949 36907 2007 36913
rect 1949 36904 1961 36907
rect 1820 36876 1961 36904
rect 1820 36864 1826 36876
rect 1949 36873 1961 36876
rect 1995 36873 2007 36907
rect 2866 36904 2872 36916
rect 2827 36876 2872 36904
rect 1949 36867 2007 36873
rect 2866 36864 2872 36876
rect 2924 36864 2930 36916
rect 3970 36904 3976 36916
rect 3931 36876 3976 36904
rect 3970 36864 3976 36876
rect 4028 36864 4034 36916
rect 5074 36904 5080 36916
rect 5035 36876 5080 36904
rect 5074 36864 5080 36876
rect 5132 36864 5138 36916
rect 6178 36864 6184 36916
rect 6236 36904 6242 36916
rect 6365 36907 6423 36913
rect 6365 36904 6377 36907
rect 6236 36876 6377 36904
rect 6236 36864 6242 36876
rect 6365 36873 6377 36876
rect 6411 36873 6423 36907
rect 7282 36904 7288 36916
rect 7243 36876 7288 36904
rect 6365 36867 6423 36873
rect 7282 36864 7288 36876
rect 7340 36864 7346 36916
rect 9490 36904 9496 36916
rect 9451 36876 9496 36904
rect 9490 36864 9496 36876
rect 9548 36864 9554 36916
rect 10594 36904 10600 36916
rect 10555 36876 10600 36904
rect 10594 36864 10600 36876
rect 10652 36864 10658 36916
rect 11698 36904 11704 36916
rect 11659 36876 11704 36904
rect 11698 36864 11704 36876
rect 11756 36864 11762 36916
rect 12802 36904 12808 36916
rect 12763 36876 12808 36904
rect 12802 36864 12808 36876
rect 12860 36864 12866 36916
rect 13906 36904 13912 36916
rect 13867 36876 13912 36904
rect 13906 36864 13912 36876
rect 13964 36864 13970 36916
rect 15010 36904 15016 36916
rect 14971 36876 15016 36904
rect 15010 36864 15016 36876
rect 15068 36864 15074 36916
rect 17218 36904 17224 36916
rect 17179 36876 17224 36904
rect 17218 36864 17224 36876
rect 17276 36864 17282 36916
rect 18322 36904 18328 36916
rect 18283 36876 18328 36904
rect 18322 36864 18328 36876
rect 18380 36864 18386 36916
rect 19334 36904 19340 36916
rect 19295 36876 19340 36904
rect 19334 36864 19340 36876
rect 19392 36864 19398 36916
rect 20530 36904 20536 36916
rect 20491 36876 20536 36904
rect 20530 36864 20536 36876
rect 20588 36864 20594 36916
rect 38013 36907 38071 36913
rect 38013 36873 38025 36907
rect 38059 36904 38071 36907
rect 38194 36904 38200 36916
rect 38059 36876 38200 36904
rect 38059 36873 38071 36876
rect 38013 36867 38071 36873
rect 38194 36864 38200 36876
rect 38252 36864 38258 36916
rect 2133 36771 2191 36777
rect 2133 36737 2145 36771
rect 2179 36768 2191 36771
rect 2406 36768 2412 36780
rect 2179 36740 2412 36768
rect 2179 36737 2191 36740
rect 2133 36731 2191 36737
rect 2406 36728 2412 36740
rect 2464 36728 2470 36780
rect 37826 36768 37832 36780
rect 37739 36740 37832 36768
rect 37826 36728 37832 36740
rect 37884 36768 37890 36780
rect 38010 36768 38016 36780
rect 37884 36740 38016 36768
rect 37884 36728 37890 36740
rect 38010 36728 38016 36740
rect 38068 36728 38074 36780
rect 19978 36524 19984 36576
rect 20036 36564 20042 36576
rect 21818 36564 21824 36576
rect 20036 36536 21824 36564
rect 20036 36524 20042 36536
rect 21818 36524 21824 36536
rect 21876 36524 21882 36576
rect 22741 36567 22799 36573
rect 22741 36533 22753 36567
rect 22787 36564 22799 36567
rect 23014 36564 23020 36576
rect 22787 36536 23020 36564
rect 22787 36533 22799 36536
rect 22741 36527 22799 36533
rect 23014 36524 23020 36536
rect 23072 36524 23078 36576
rect 25041 36567 25099 36573
rect 25041 36533 25053 36567
rect 25087 36564 25099 36567
rect 25130 36564 25136 36576
rect 25087 36536 25136 36564
rect 25087 36533 25099 36536
rect 25041 36527 25099 36533
rect 25130 36524 25136 36536
rect 25188 36524 25194 36576
rect 26053 36567 26111 36573
rect 26053 36533 26065 36567
rect 26099 36564 26111 36567
rect 26142 36564 26148 36576
rect 26099 36536 26148 36564
rect 26099 36533 26111 36536
rect 26053 36527 26111 36533
rect 26142 36524 26148 36536
rect 26200 36524 26206 36576
rect 27157 36567 27215 36573
rect 27157 36533 27169 36567
rect 27203 36564 27215 36567
rect 27246 36564 27252 36576
rect 27203 36536 27252 36564
rect 27203 36533 27215 36536
rect 27157 36527 27215 36533
rect 27246 36524 27252 36536
rect 27304 36524 27310 36576
rect 28166 36564 28172 36576
rect 28127 36536 28172 36564
rect 28166 36524 28172 36536
rect 28224 36524 28230 36576
rect 29362 36564 29368 36576
rect 29323 36536 29368 36564
rect 29362 36524 29368 36536
rect 29420 36524 29426 36576
rect 30374 36564 30380 36576
rect 30335 36536 30380 36564
rect 30374 36524 30380 36536
rect 30432 36524 30438 36576
rect 32769 36567 32827 36573
rect 32769 36533 32781 36567
rect 32815 36564 32827 36567
rect 32858 36564 32864 36576
rect 32815 36536 32864 36564
rect 32815 36533 32827 36536
rect 32769 36527 32827 36533
rect 32858 36524 32864 36536
rect 32916 36524 32922 36576
rect 33781 36567 33839 36573
rect 33781 36533 33793 36567
rect 33827 36564 33839 36567
rect 33870 36564 33876 36576
rect 33827 36536 33876 36564
rect 33827 36533 33839 36536
rect 33781 36527 33839 36533
rect 33870 36524 33876 36536
rect 33928 36524 33934 36576
rect 34790 36564 34796 36576
rect 34751 36536 34796 36564
rect 34790 36524 34796 36536
rect 34848 36524 34854 36576
rect 35894 36524 35900 36576
rect 35952 36564 35958 36576
rect 37366 36564 37372 36576
rect 35952 36536 35997 36564
rect 37327 36536 37372 36564
rect 35952 36524 35958 36536
rect 37366 36524 37372 36536
rect 37424 36524 37430 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1302 36320 1308 36372
rect 1360 36360 1366 36372
rect 1581 36363 1639 36369
rect 1581 36360 1593 36363
rect 1360 36332 1593 36360
rect 1360 36320 1366 36332
rect 1581 36329 1593 36332
rect 1627 36329 1639 36363
rect 1581 36323 1639 36329
rect 38013 36363 38071 36369
rect 38013 36329 38025 36363
rect 38059 36360 38071 36363
rect 39298 36360 39304 36372
rect 38059 36332 39304 36360
rect 38059 36329 38071 36332
rect 38013 36323 38071 36329
rect 39298 36320 39304 36332
rect 39356 36320 39362 36372
rect 37829 36159 37887 36165
rect 37829 36156 37841 36159
rect 37292 36128 37841 36156
rect 37292 36032 37320 36128
rect 37829 36125 37841 36128
rect 37875 36125 37887 36159
rect 37829 36119 37887 36125
rect 2317 36023 2375 36029
rect 2317 35989 2329 36023
rect 2363 36020 2375 36023
rect 2406 36020 2412 36032
rect 2363 35992 2412 36020
rect 2363 35989 2375 35992
rect 2317 35983 2375 35989
rect 2406 35980 2412 35992
rect 2464 35980 2470 36032
rect 37274 36020 37280 36032
rect 37235 35992 37280 36020
rect 37274 35980 37280 35992
rect 37332 35980 37338 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 1578 30200 1584 30252
rect 1636 30240 1642 30252
rect 1857 30243 1915 30249
rect 1857 30240 1869 30243
rect 1636 30212 1869 30240
rect 1636 30200 1642 30212
rect 1857 30209 1869 30212
rect 1903 30209 1915 30243
rect 1857 30203 1915 30209
rect 2038 30104 2044 30116
rect 1999 30076 2044 30104
rect 2038 30064 2044 30076
rect 2096 30064 2102 30116
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 7558 22080 7564 22092
rect 3200 22052 7564 22080
rect 3200 22040 3206 22052
rect 7558 22040 7564 22052
rect 7616 22040 7622 22092
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 10505 20859 10563 20865
rect 10505 20825 10517 20859
rect 10551 20856 10563 20859
rect 11422 20856 11428 20868
rect 10551 20828 11428 20856
rect 10551 20825 10563 20828
rect 10505 20819 10563 20825
rect 11422 20816 11428 20828
rect 11480 20816 11486 20868
rect 11057 20791 11115 20797
rect 11057 20757 11069 20791
rect 11103 20788 11115 20791
rect 11793 20791 11851 20797
rect 11793 20788 11805 20791
rect 11103 20760 11805 20788
rect 11103 20757 11115 20760
rect 11057 20751 11115 20757
rect 11793 20757 11805 20760
rect 11839 20788 11851 20791
rect 12250 20788 12256 20800
rect 11839 20760 12256 20788
rect 11839 20757 11851 20760
rect 11793 20751 11851 20757
rect 12250 20748 12256 20760
rect 12308 20788 12314 20800
rect 12713 20791 12771 20797
rect 12713 20788 12725 20791
rect 12308 20760 12725 20788
rect 12308 20748 12314 20760
rect 12713 20757 12725 20760
rect 12759 20757 12771 20791
rect 13354 20788 13360 20800
rect 13315 20760 13360 20788
rect 12713 20751 12771 20757
rect 13354 20748 13360 20760
rect 13412 20748 13418 20800
rect 16574 20788 16580 20800
rect 16535 20760 16580 20788
rect 16574 20748 16580 20760
rect 16632 20748 16638 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 10376 20556 10885 20584
rect 10376 20544 10382 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 10873 20547 10931 20553
rect 13265 20587 13323 20593
rect 13265 20553 13277 20587
rect 13311 20584 13323 20587
rect 14185 20587 14243 20593
rect 14185 20584 14197 20587
rect 13311 20556 14197 20584
rect 13311 20553 13323 20556
rect 13265 20547 13323 20553
rect 14185 20553 14197 20556
rect 14231 20584 14243 20587
rect 16758 20584 16764 20596
rect 14231 20556 16764 20584
rect 14231 20553 14243 20556
rect 14185 20547 14243 20553
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20584 17095 20587
rect 17957 20587 18015 20593
rect 17957 20584 17969 20587
rect 17083 20556 17969 20584
rect 17083 20553 17095 20556
rect 17037 20547 17095 20553
rect 17957 20553 17969 20556
rect 18003 20584 18015 20587
rect 18414 20584 18420 20596
rect 18003 20556 18420 20584
rect 18003 20553 18015 20556
rect 17957 20547 18015 20553
rect 18414 20544 18420 20556
rect 18472 20544 18478 20596
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 10226 20448 10232 20460
rect 10091 20420 10232 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 12250 20448 12256 20460
rect 12211 20420 12256 20448
rect 12250 20408 12256 20420
rect 12308 20448 12314 20460
rect 12308 20420 13492 20448
rect 12308 20408 12314 20420
rect 13354 20380 13360 20392
rect 13315 20352 13360 20380
rect 13354 20340 13360 20352
rect 13412 20340 13418 20392
rect 13464 20389 13492 20420
rect 13449 20383 13507 20389
rect 13449 20349 13461 20383
rect 13495 20380 13507 20383
rect 16025 20383 16083 20389
rect 16025 20380 16037 20383
rect 13495 20352 16037 20380
rect 13495 20349 13507 20352
rect 13449 20343 13507 20349
rect 16025 20349 16037 20352
rect 16071 20349 16083 20383
rect 16025 20343 16083 20349
rect 16040 20312 16068 20343
rect 16298 20340 16304 20392
rect 16356 20380 16362 20392
rect 17129 20383 17187 20389
rect 17129 20380 17141 20383
rect 16356 20352 17141 20380
rect 16356 20340 16362 20352
rect 17129 20349 17141 20352
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 17221 20383 17279 20389
rect 17221 20349 17233 20383
rect 17267 20349 17279 20383
rect 17221 20343 17279 20349
rect 17236 20312 17264 20343
rect 17402 20312 17408 20324
rect 16040 20284 17408 20312
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 9861 20247 9919 20253
rect 9861 20244 9873 20247
rect 9456 20216 9873 20244
rect 9456 20204 9462 20216
rect 9861 20213 9873 20216
rect 9907 20213 9919 20247
rect 9861 20207 9919 20213
rect 10594 20204 10600 20256
rect 10652 20244 10658 20256
rect 11977 20247 12035 20253
rect 11977 20244 11989 20247
rect 10652 20216 11989 20244
rect 10652 20204 10658 20216
rect 11977 20213 11989 20216
rect 12023 20213 12035 20247
rect 12894 20244 12900 20256
rect 12855 20216 12900 20244
rect 11977 20207 12035 20213
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 16666 20244 16672 20256
rect 16627 20216 16672 20244
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 4706 20040 4712 20052
rect 4387 20012 4712 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 4706 20000 4712 20012
rect 4764 20000 4770 20052
rect 7837 20043 7895 20049
rect 7837 20009 7849 20043
rect 7883 20040 7895 20043
rect 8294 20040 8300 20052
rect 7883 20012 8300 20040
rect 7883 20009 7895 20012
rect 7837 20003 7895 20009
rect 8294 20000 8300 20012
rect 8352 20040 8358 20052
rect 9582 20040 9588 20052
rect 8352 20012 9588 20040
rect 8352 20000 8358 20012
rect 9582 20000 9588 20012
rect 9640 20000 9646 20052
rect 14737 20043 14795 20049
rect 14737 20040 14749 20043
rect 11532 20012 14749 20040
rect 10594 19904 10600 19916
rect 10555 19876 10600 19904
rect 10594 19864 10600 19876
rect 10652 19864 10658 19916
rect 10318 19836 10324 19848
rect 10279 19808 10324 19836
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 11532 19845 11560 20012
rect 14737 20009 14749 20012
rect 14783 20040 14795 20043
rect 15838 20040 15844 20052
rect 14783 20012 15844 20040
rect 14783 20009 14795 20012
rect 14737 20003 14795 20009
rect 15838 20000 15844 20012
rect 15896 20000 15902 20052
rect 18141 20043 18199 20049
rect 18141 20040 18153 20043
rect 17236 20012 18153 20040
rect 11698 19904 11704 19916
rect 11659 19876 11704 19904
rect 11698 19864 11704 19876
rect 11756 19904 11762 19916
rect 12250 19904 12256 19916
rect 11756 19876 12256 19904
rect 11756 19864 11762 19876
rect 12250 19864 12256 19876
rect 12308 19904 12314 19916
rect 12989 19907 13047 19913
rect 12989 19904 13001 19907
rect 12308 19876 13001 19904
rect 12308 19864 12314 19876
rect 12989 19873 13001 19876
rect 13035 19904 13047 19907
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13035 19876 14105 19904
rect 13035 19873 13047 19876
rect 12989 19867 13047 19873
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19836 15439 19839
rect 16666 19836 16672 19848
rect 15427 19808 16672 19836
rect 15427 19805 15439 19808
rect 15381 19799 15439 19805
rect 16666 19796 16672 19808
rect 16724 19796 16730 19848
rect 17236 19845 17264 20012
rect 18141 20009 18153 20012
rect 18187 20040 18199 20043
rect 19426 20040 19432 20052
rect 18187 20012 19432 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 17402 19904 17408 19916
rect 17363 19876 17408 19904
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19805 17279 19839
rect 17221 19799 17279 19805
rect 9493 19771 9551 19777
rect 9493 19737 9505 19771
rect 9539 19768 9551 19771
rect 9539 19740 10456 19768
rect 9539 19737 9551 19740
rect 9493 19731 9551 19737
rect 10428 19712 10456 19740
rect 11422 19728 11428 19780
rect 11480 19768 11486 19780
rect 11609 19771 11667 19777
rect 11609 19768 11621 19771
rect 11480 19740 11621 19768
rect 11480 19728 11486 19740
rect 11609 19737 11621 19740
rect 11655 19737 11667 19771
rect 11609 19731 11667 19737
rect 12713 19771 12771 19777
rect 12713 19737 12725 19771
rect 12759 19768 12771 19771
rect 13814 19768 13820 19780
rect 12759 19740 13820 19768
rect 12759 19737 12771 19740
rect 12713 19731 12771 19737
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 16574 19728 16580 19780
rect 16632 19768 16638 19780
rect 17313 19771 17371 19777
rect 17313 19768 17325 19771
rect 16632 19740 17325 19768
rect 16632 19728 16638 19740
rect 17313 19737 17325 19740
rect 17359 19737 17371 19771
rect 17313 19731 17371 19737
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 8297 19703 8355 19709
rect 8297 19700 8309 19703
rect 7708 19672 8309 19700
rect 7708 19660 7714 19672
rect 8297 19669 8309 19672
rect 8343 19669 8355 19703
rect 9950 19700 9956 19712
rect 9911 19672 9956 19700
rect 8297 19663 8355 19669
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 10410 19700 10416 19712
rect 10371 19672 10416 19700
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 11146 19700 11152 19712
rect 11107 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 11848 19672 12357 19700
rect 11848 19660 11854 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 12345 19663 12403 19669
rect 12805 19703 12863 19709
rect 12805 19669 12817 19703
rect 12851 19700 12863 19703
rect 13722 19700 13728 19712
rect 12851 19672 13728 19700
rect 12851 19669 12863 19672
rect 12805 19663 12863 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 15194 19700 15200 19712
rect 15155 19672 15200 19700
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 15654 19660 15660 19712
rect 15712 19700 15718 19712
rect 16298 19700 16304 19712
rect 15712 19672 16304 19700
rect 15712 19660 15718 19672
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 16850 19700 16856 19712
rect 16811 19672 16856 19700
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 2958 19456 2964 19508
rect 3016 19496 3022 19508
rect 3421 19499 3479 19505
rect 3421 19496 3433 19499
rect 3016 19468 3433 19496
rect 3016 19456 3022 19468
rect 3421 19465 3433 19468
rect 3467 19465 3479 19499
rect 3421 19459 3479 19465
rect 3789 19499 3847 19505
rect 3789 19465 3801 19499
rect 3835 19496 3847 19499
rect 4706 19496 4712 19508
rect 3835 19468 4712 19496
rect 3835 19465 3847 19468
rect 3789 19459 3847 19465
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 7653 19499 7711 19505
rect 7653 19465 7665 19499
rect 7699 19496 7711 19499
rect 8294 19496 8300 19508
rect 7699 19468 8300 19496
rect 7699 19465 7711 19468
rect 7653 19459 7711 19465
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 10226 19496 10232 19508
rect 10187 19468 10232 19496
rect 10226 19456 10232 19468
rect 10284 19456 10290 19508
rect 10597 19499 10655 19505
rect 10597 19465 10609 19499
rect 10643 19496 10655 19499
rect 11514 19496 11520 19508
rect 10643 19468 11520 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 9769 19431 9827 19437
rect 9769 19397 9781 19431
rect 9815 19428 9827 19431
rect 10612 19428 10640 19459
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 15749 19499 15807 19505
rect 15749 19496 15761 19499
rect 12860 19468 15761 19496
rect 12860 19456 12866 19468
rect 15749 19465 15761 19468
rect 15795 19465 15807 19499
rect 15749 19459 15807 19465
rect 16945 19499 17003 19505
rect 16945 19465 16957 19499
rect 16991 19465 17003 19499
rect 16945 19459 17003 19465
rect 17313 19499 17371 19505
rect 17313 19465 17325 19499
rect 17359 19496 17371 19499
rect 18233 19499 18291 19505
rect 18233 19496 18245 19499
rect 17359 19468 18245 19496
rect 17359 19465 17371 19468
rect 17313 19459 17371 19465
rect 18233 19465 18245 19468
rect 18279 19496 18291 19499
rect 20622 19496 20628 19508
rect 18279 19468 20628 19496
rect 18279 19465 18291 19468
rect 18233 19459 18291 19465
rect 9815 19400 10640 19428
rect 9815 19397 9827 19400
rect 9769 19391 9827 19397
rect 10686 19388 10692 19440
rect 10744 19388 10750 19440
rect 13265 19431 13323 19437
rect 13265 19397 13277 19431
rect 13311 19428 13323 19431
rect 13814 19428 13820 19440
rect 13311 19400 13820 19428
rect 13311 19397 13323 19400
rect 13265 19391 13323 19397
rect 13814 19388 13820 19400
rect 13872 19428 13878 19440
rect 15102 19428 15108 19440
rect 13872 19400 15108 19428
rect 13872 19388 13878 19400
rect 15102 19388 15108 19400
rect 15160 19388 15166 19440
rect 7650 19320 7656 19372
rect 7708 19360 7714 19372
rect 7745 19363 7803 19369
rect 7745 19360 7757 19363
rect 7708 19332 7757 19360
rect 7708 19320 7714 19332
rect 7745 19329 7757 19332
rect 7791 19329 7803 19363
rect 7745 19323 7803 19329
rect 8849 19363 8907 19369
rect 8849 19329 8861 19363
rect 8895 19360 8907 19363
rect 9674 19360 9680 19372
rect 8895 19332 9680 19360
rect 8895 19329 8907 19332
rect 8849 19323 8907 19329
rect 9674 19320 9680 19332
rect 9732 19360 9738 19372
rect 10704 19360 10732 19388
rect 9732 19332 10732 19360
rect 12253 19363 12311 19369
rect 9732 19320 9738 19332
rect 12253 19329 12265 19363
rect 12299 19360 12311 19363
rect 12710 19360 12716 19372
rect 12299 19332 12716 19360
rect 12299 19329 12311 19332
rect 12253 19323 12311 19329
rect 12710 19320 12716 19332
rect 12768 19360 12774 19372
rect 13906 19360 13912 19372
rect 12768 19332 13912 19360
rect 12768 19320 12774 19332
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19360 15991 19363
rect 16960 19360 16988 19459
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 15979 19332 16988 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 3881 19295 3939 19301
rect 3881 19261 3893 19295
rect 3927 19261 3939 19295
rect 4062 19292 4068 19304
rect 4023 19264 4068 19292
rect 3881 19255 3939 19261
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 3326 19156 3332 19168
rect 3007 19128 3332 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 3326 19116 3332 19128
rect 3384 19156 3390 19168
rect 3896 19156 3924 19255
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5534 19292 5540 19304
rect 5123 19264 5540 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5534 19252 5540 19264
rect 5592 19292 5598 19304
rect 6362 19292 6368 19304
rect 5592 19264 6368 19292
rect 5592 19252 5598 19264
rect 6362 19252 6368 19264
rect 6420 19252 6426 19304
rect 7837 19295 7895 19301
rect 7837 19261 7849 19295
rect 7883 19261 7895 19295
rect 8938 19292 8944 19304
rect 8899 19264 8944 19292
rect 7837 19255 7895 19261
rect 7852 19224 7880 19255
rect 8938 19252 8944 19264
rect 8996 19252 9002 19304
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19261 9183 19295
rect 10686 19292 10692 19304
rect 10647 19264 10692 19292
rect 9125 19255 9183 19261
rect 7926 19224 7932 19236
rect 7839 19196 7932 19224
rect 7926 19184 7932 19196
rect 7984 19224 7990 19236
rect 9140 19224 9168 19255
rect 10686 19252 10692 19264
rect 10744 19252 10750 19304
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19261 10839 19295
rect 10781 19255 10839 19261
rect 10594 19224 10600 19236
rect 7984 19196 10600 19224
rect 7984 19184 7990 19196
rect 10594 19184 10600 19196
rect 10652 19224 10658 19236
rect 10796 19224 10824 19255
rect 11974 19252 11980 19304
rect 12032 19292 12038 19304
rect 12345 19295 12403 19301
rect 12345 19292 12357 19295
rect 12032 19264 12357 19292
rect 12032 19252 12038 19264
rect 12345 19261 12357 19264
rect 12391 19261 12403 19295
rect 12345 19255 12403 19261
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 10652 19196 10824 19224
rect 10652 19184 10658 19196
rect 11698 19184 11704 19236
rect 11756 19224 11762 19236
rect 12452 19224 12480 19255
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 17368 19264 17417 19292
rect 17368 19252 17374 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 17552 19264 17597 19292
rect 17552 19252 17558 19264
rect 11756 19196 12480 19224
rect 11756 19184 11762 19196
rect 7282 19156 7288 19168
rect 3384 19128 3924 19156
rect 7243 19128 7288 19156
rect 3384 19116 3390 19128
rect 7282 19116 7288 19128
rect 7340 19116 7346 19168
rect 8478 19156 8484 19168
rect 8439 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11885 19159 11943 19165
rect 11885 19156 11897 19159
rect 11112 19128 11897 19156
rect 11112 19116 11118 19128
rect 11885 19125 11897 19128
rect 11931 19125 11943 19159
rect 13814 19156 13820 19168
rect 13775 19128 13820 19156
rect 11885 19119 11943 19125
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 6641 18955 6699 18961
rect 6641 18952 6653 18955
rect 6012 18924 6653 18952
rect 4062 18844 4068 18896
rect 4120 18884 4126 18896
rect 4120 18856 5948 18884
rect 4120 18844 4126 18856
rect 4816 18825 4844 18856
rect 5920 18828 5948 18856
rect 4801 18819 4859 18825
rect 4801 18785 4813 18819
rect 4847 18785 4859 18819
rect 5902 18816 5908 18828
rect 5863 18788 5908 18816
rect 4801 18779 4859 18785
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 5534 18748 5540 18760
rect 4571 18720 5540 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 6012 18748 6040 18924
rect 6641 18921 6653 18924
rect 6687 18952 6699 18955
rect 7374 18952 7380 18964
rect 6687 18924 7380 18952
rect 6687 18921 6699 18924
rect 6641 18915 6699 18921
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 9490 18912 9496 18964
rect 9548 18952 9554 18964
rect 11609 18955 11667 18961
rect 11609 18952 11621 18955
rect 9548 18924 11621 18952
rect 9548 18912 9554 18924
rect 11609 18921 11621 18924
rect 11655 18921 11667 18955
rect 12710 18952 12716 18964
rect 12671 18924 12716 18952
rect 11609 18915 11667 18921
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 16761 18955 16819 18961
rect 16761 18921 16773 18955
rect 16807 18952 16819 18955
rect 17221 18955 17279 18961
rect 17221 18952 17233 18955
rect 16807 18924 17233 18952
rect 16807 18921 16819 18924
rect 16761 18915 16819 18921
rect 17221 18921 17233 18924
rect 17267 18952 17279 18955
rect 17402 18952 17408 18964
rect 17267 18924 17408 18952
rect 17267 18921 17279 18924
rect 17221 18915 17279 18921
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 9306 18844 9312 18896
rect 9364 18884 9370 18896
rect 10321 18887 10379 18893
rect 10321 18884 10333 18887
rect 9364 18856 10333 18884
rect 9364 18844 9370 18856
rect 10321 18853 10333 18856
rect 10367 18853 10379 18887
rect 10321 18847 10379 18853
rect 11146 18844 11152 18896
rect 11204 18844 11210 18896
rect 7926 18816 7932 18828
rect 5767 18720 6040 18748
rect 6886 18788 7932 18816
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 3237 18683 3295 18689
rect 3237 18649 3249 18683
rect 3283 18680 3295 18683
rect 3694 18680 3700 18692
rect 3283 18652 3700 18680
rect 3283 18649 3295 18652
rect 3237 18643 3295 18649
rect 3694 18640 3700 18652
rect 3752 18680 3758 18692
rect 4617 18683 4675 18689
rect 4617 18680 4629 18683
rect 3752 18652 4629 18680
rect 3752 18640 3758 18652
rect 4617 18649 4629 18652
rect 4663 18649 4675 18683
rect 4617 18643 4675 18649
rect 5166 18640 5172 18692
rect 5224 18680 5230 18692
rect 5813 18683 5871 18689
rect 5813 18680 5825 18683
rect 5224 18652 5825 18680
rect 5224 18640 5230 18652
rect 5813 18649 5825 18652
rect 5859 18649 5871 18683
rect 5813 18643 5871 18649
rect 5902 18640 5908 18692
rect 5960 18680 5966 18692
rect 6886 18680 6914 18788
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 9217 18819 9275 18825
rect 9217 18785 9229 18819
rect 9263 18816 9275 18819
rect 9674 18816 9680 18828
rect 9263 18788 9680 18816
rect 9263 18785 9275 18788
rect 9217 18779 9275 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11164 18816 11192 18844
rect 12894 18816 12900 18828
rect 9876 18788 11192 18816
rect 11624 18788 12900 18816
rect 7653 18751 7711 18757
rect 7653 18717 7665 18751
rect 7699 18748 7711 18751
rect 8294 18748 8300 18760
rect 7699 18720 8300 18748
rect 7699 18717 7711 18720
rect 7653 18711 7711 18717
rect 8294 18708 8300 18720
rect 8352 18748 8358 18760
rect 8846 18748 8852 18760
rect 8352 18720 8852 18748
rect 8352 18708 8358 18720
rect 8846 18708 8852 18720
rect 8904 18708 8910 18760
rect 9876 18757 9904 18788
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18748 10563 18751
rect 11054 18748 11060 18760
rect 10551 18720 11060 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18748 11207 18751
rect 11624 18748 11652 18788
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 11790 18748 11796 18760
rect 11195 18720 11652 18748
rect 11751 18720 11796 18748
rect 11195 18717 11207 18720
rect 11149 18711 11207 18717
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18748 15899 18751
rect 16850 18748 16856 18760
rect 15887 18720 16856 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 5960 18652 6914 18680
rect 5960 18640 5966 18652
rect 9582 18640 9588 18692
rect 9640 18680 9646 18692
rect 9640 18652 11008 18680
rect 9640 18640 9646 18652
rect 3418 18572 3424 18624
rect 3476 18612 3482 18624
rect 4157 18615 4215 18621
rect 4157 18612 4169 18615
rect 3476 18584 4169 18612
rect 3476 18572 3482 18584
rect 4157 18581 4169 18584
rect 4203 18581 4215 18615
rect 5350 18612 5356 18624
rect 5311 18584 5356 18612
rect 4157 18575 4215 18581
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 7285 18615 7343 18621
rect 7285 18612 7297 18615
rect 7156 18584 7297 18612
rect 7156 18572 7162 18584
rect 7285 18581 7297 18584
rect 7331 18581 7343 18615
rect 7285 18575 7343 18581
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 7800 18584 7845 18612
rect 7800 18572 7806 18584
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 10980 18621 11008 18652
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 9272 18584 9689 18612
rect 9272 18572 9278 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 9677 18575 9735 18581
rect 10965 18615 11023 18621
rect 10965 18581 10977 18615
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 15657 18615 15715 18621
rect 15657 18612 15669 18615
rect 14424 18584 15669 18612
rect 14424 18572 14430 18584
rect 15657 18581 15669 18584
rect 15703 18581 15715 18615
rect 15657 18575 15715 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 3881 18411 3939 18417
rect 3881 18377 3893 18411
rect 3927 18377 3939 18411
rect 3881 18371 3939 18377
rect 4249 18411 4307 18417
rect 4249 18377 4261 18411
rect 4295 18408 4307 18411
rect 4614 18408 4620 18420
rect 4295 18380 4620 18408
rect 4295 18377 4307 18380
rect 4249 18371 4307 18377
rect 3896 18340 3924 18371
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 8386 18408 8392 18420
rect 8299 18380 8392 18408
rect 8386 18368 8392 18380
rect 8444 18408 8450 18420
rect 8938 18408 8944 18420
rect 8444 18380 8944 18408
rect 8444 18368 8450 18380
rect 8938 18368 8944 18380
rect 8996 18368 9002 18420
rect 2792 18312 3924 18340
rect 2792 18281 2820 18312
rect 7742 18300 7748 18352
rect 7800 18340 7806 18352
rect 8202 18340 8208 18352
rect 7800 18312 8208 18340
rect 7800 18300 7806 18312
rect 8202 18300 8208 18312
rect 8260 18340 8266 18352
rect 8849 18343 8907 18349
rect 8849 18340 8861 18343
rect 8260 18312 8861 18340
rect 8260 18300 8266 18312
rect 8849 18309 8861 18312
rect 8895 18309 8907 18343
rect 8849 18303 8907 18309
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18241 2835 18275
rect 3418 18272 3424 18284
rect 3379 18244 3424 18272
rect 2777 18235 2835 18241
rect 3418 18232 3424 18244
rect 3476 18232 3482 18284
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18272 6883 18275
rect 7282 18272 7288 18284
rect 6871 18244 7288 18272
rect 6871 18241 6883 18244
rect 6825 18235 6883 18241
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18272 7527 18275
rect 8478 18272 8484 18284
rect 7515 18244 8484 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 9950 18272 9956 18284
rect 9911 18244 9956 18272
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 4341 18207 4399 18213
rect 4341 18204 4353 18207
rect 3844 18176 4353 18204
rect 3844 18164 3850 18176
rect 4341 18173 4353 18176
rect 4387 18173 4399 18207
rect 4341 18167 4399 18173
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 5902 18204 5908 18216
rect 4571 18176 5908 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 5902 18164 5908 18176
rect 5960 18164 5966 18216
rect 2590 18068 2596 18080
rect 2551 18040 2596 18068
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 3234 18068 3240 18080
rect 3195 18040 3240 18068
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 5166 18068 5172 18080
rect 5127 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 6638 18068 6644 18080
rect 6599 18040 6644 18068
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 6730 18028 6736 18080
rect 6788 18068 6794 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 6788 18040 7297 18068
rect 6788 18028 6794 18040
rect 7285 18037 7297 18040
rect 7331 18037 7343 18071
rect 10134 18068 10140 18080
rect 10095 18040 10140 18068
rect 7285 18031 7343 18037
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10318 18028 10324 18080
rect 10376 18068 10382 18080
rect 10686 18068 10692 18080
rect 10376 18040 10692 18068
rect 10376 18028 10382 18040
rect 10686 18028 10692 18040
rect 10744 18068 10750 18080
rect 10873 18071 10931 18077
rect 10873 18068 10885 18071
rect 10744 18040 10885 18068
rect 10744 18028 10750 18040
rect 10873 18037 10885 18040
rect 10919 18037 10931 18071
rect 10873 18031 10931 18037
rect 11514 18028 11520 18080
rect 11572 18068 11578 18080
rect 11698 18068 11704 18080
rect 11572 18040 11704 18068
rect 11572 18028 11578 18040
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 12253 18071 12311 18077
rect 12253 18068 12265 18071
rect 12032 18040 12265 18068
rect 12032 18028 12038 18040
rect 12253 18037 12265 18040
rect 12299 18037 12311 18071
rect 12253 18031 12311 18037
rect 16761 18071 16819 18077
rect 16761 18037 16773 18071
rect 16807 18068 16819 18071
rect 17310 18068 17316 18080
rect 16807 18040 17316 18068
rect 16807 18037 16819 18040
rect 16761 18031 16819 18037
rect 17310 18028 17316 18040
rect 17368 18068 17374 18080
rect 17862 18068 17868 18080
rect 17368 18040 17868 18068
rect 17368 18028 17374 18040
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 4614 17824 4620 17876
rect 4672 17864 4678 17876
rect 4801 17867 4859 17873
rect 4801 17864 4813 17867
rect 4672 17836 4813 17864
rect 4672 17824 4678 17836
rect 4801 17833 4813 17836
rect 4847 17833 4859 17867
rect 4801 17827 4859 17833
rect 8205 17867 8263 17873
rect 8205 17833 8217 17867
rect 8251 17864 8263 17867
rect 8294 17864 8300 17876
rect 8251 17836 8300 17864
rect 8251 17833 8263 17836
rect 8205 17827 8263 17833
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 2958 17660 2964 17672
rect 2919 17632 2964 17660
rect 2958 17620 2964 17632
rect 3016 17620 3022 17672
rect 4341 17663 4399 17669
rect 4341 17629 4353 17663
rect 4387 17660 4399 17663
rect 5350 17660 5356 17672
rect 4387 17632 5356 17660
rect 4387 17629 4399 17632
rect 4341 17623 4399 17629
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 6733 17663 6791 17669
rect 6733 17629 6745 17663
rect 6779 17660 6791 17663
rect 7098 17660 7104 17672
rect 6779 17632 7104 17660
rect 6779 17629 6791 17632
rect 6733 17623 6791 17629
rect 7098 17620 7104 17632
rect 7156 17620 7162 17672
rect 2777 17527 2835 17533
rect 2777 17493 2789 17527
rect 2823 17524 2835 17527
rect 2866 17524 2872 17536
rect 2823 17496 2872 17524
rect 2823 17493 2835 17496
rect 2777 17487 2835 17493
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 4157 17527 4215 17533
rect 4157 17493 4169 17527
rect 4203 17524 4215 17527
rect 4614 17524 4620 17536
rect 4203 17496 4620 17524
rect 4203 17493 4215 17496
rect 4157 17487 4215 17493
rect 4614 17484 4620 17496
rect 4672 17484 4678 17536
rect 6546 17524 6552 17536
rect 6507 17496 6552 17524
rect 6546 17484 6552 17496
rect 6604 17484 6610 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 3786 17320 3792 17332
rect 3747 17292 3792 17320
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 14544 17187 14602 17193
rect 14544 17153 14556 17187
rect 14590 17184 14602 17187
rect 18046 17184 18052 17196
rect 14590 17156 18052 17184
rect 14590 17153 14602 17156
rect 14544 17147 14602 17153
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 13722 17076 13728 17128
rect 13780 17116 13786 17128
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 13780 17088 14289 17116
rect 13780 17076 13786 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 22278 16980 22284 16992
rect 15703 16952 22284 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 5626 16640 5632 16652
rect 5587 16612 5632 16640
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 5902 16640 5908 16652
rect 5736 16612 5908 16640
rect 5534 16572 5540 16584
rect 5495 16544 5540 16572
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 5736 16581 5764 16612
rect 5902 16600 5908 16612
rect 5960 16600 5966 16652
rect 27246 16640 27252 16652
rect 19904 16612 27252 16640
rect 5721 16575 5779 16581
rect 5721 16541 5733 16575
rect 5767 16574 5779 16575
rect 5767 16546 5801 16574
rect 8938 16572 8944 16584
rect 5767 16541 5779 16546
rect 8899 16544 8944 16572
rect 5721 16535 5779 16541
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12207 16544 12572 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 12544 16516 12572 16544
rect 13722 16532 13728 16584
rect 13780 16572 13786 16584
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 13780 16544 14381 16572
rect 13780 16532 13786 16544
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 15194 16572 15200 16584
rect 14369 16535 14427 16541
rect 14476 16544 15200 16572
rect 9208 16507 9266 16513
rect 9208 16473 9220 16507
rect 9254 16504 9266 16507
rect 9398 16504 9404 16516
rect 9254 16476 9404 16504
rect 9254 16473 9266 16476
rect 9208 16467 9266 16473
rect 9398 16464 9404 16476
rect 9456 16464 9462 16516
rect 12428 16507 12486 16513
rect 12428 16473 12440 16507
rect 12474 16473 12486 16507
rect 12428 16467 12486 16473
rect 10318 16436 10324 16448
rect 10279 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 12452 16436 12480 16467
rect 12526 16464 12532 16516
rect 12584 16464 12590 16516
rect 14476 16504 14504 16544
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 12636 16476 14504 16504
rect 14636 16507 14694 16513
rect 12636 16436 12664 16476
rect 14636 16473 14648 16507
rect 14682 16504 14694 16507
rect 19242 16504 19248 16516
rect 14682 16476 19248 16504
rect 14682 16473 14694 16476
rect 14636 16467 14694 16473
rect 19242 16464 19248 16476
rect 19300 16464 19306 16516
rect 13538 16436 13544 16448
rect 12452 16408 12664 16436
rect 13499 16408 13544 16436
rect 13538 16396 13544 16408
rect 13596 16436 13602 16448
rect 15654 16436 15660 16448
rect 13596 16408 15660 16436
rect 13596 16396 13602 16408
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 19334 16436 19340 16448
rect 15795 16408 19340 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 19334 16396 19340 16408
rect 19392 16396 19398 16448
rect 19426 16396 19432 16448
rect 19484 16436 19490 16448
rect 19904 16445 19932 16612
rect 27246 16600 27252 16612
rect 27304 16600 27310 16652
rect 19889 16439 19947 16445
rect 19889 16436 19901 16439
rect 19484 16408 19901 16436
rect 19484 16396 19490 16408
rect 19889 16405 19901 16408
rect 19935 16405 19947 16439
rect 19889 16399 19947 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 2590 16192 2596 16244
rect 2648 16232 2654 16244
rect 13909 16235 13967 16241
rect 2648 16204 2728 16232
rect 2648 16192 2654 16204
rect 2700 16173 2728 16204
rect 13909 16201 13921 16235
rect 13955 16232 13967 16235
rect 17862 16232 17868 16244
rect 13955 16204 17868 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 19245 16235 19303 16241
rect 19245 16201 19257 16235
rect 19291 16201 19303 16235
rect 19245 16195 19303 16201
rect 20073 16235 20131 16241
rect 20073 16201 20085 16235
rect 20119 16201 20131 16235
rect 20073 16195 20131 16201
rect 6638 16173 6644 16176
rect 2676 16167 2734 16173
rect 2676 16133 2688 16167
rect 2722 16133 2734 16167
rect 6632 16164 6644 16173
rect 6599 16136 6644 16164
rect 2676 16127 2734 16133
rect 6632 16127 6644 16136
rect 6638 16124 6644 16127
rect 6696 16124 6702 16176
rect 9306 16124 9312 16176
rect 9364 16164 9370 16176
rect 12802 16173 12808 16176
rect 9462 16167 9520 16173
rect 9462 16164 9474 16167
rect 9364 16136 9474 16164
rect 9364 16124 9370 16136
rect 9462 16133 9474 16136
rect 9508 16133 9520 16167
rect 12796 16164 12808 16173
rect 12763 16136 12808 16164
rect 9462 16127 9520 16133
rect 12796 16127 12808 16136
rect 12802 16124 12808 16127
rect 12860 16124 12866 16176
rect 14636 16167 14694 16173
rect 14636 16133 14648 16167
rect 14682 16164 14694 16167
rect 19260 16164 19288 16195
rect 14682 16136 19288 16164
rect 14682 16133 14694 16136
rect 14636 16127 14694 16133
rect 8938 16056 8944 16108
rect 8996 16096 9002 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 8996 16068 9229 16096
rect 8996 16056 9002 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16096 19487 16099
rect 20088 16096 20116 16195
rect 20438 16096 20444 16108
rect 19475 16068 20116 16096
rect 20399 16068 20444 16096
rect 19475 16065 19487 16068
rect 19429 16059 19487 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 2409 16031 2467 16037
rect 2409 15997 2421 16031
rect 2455 15997 2467 16031
rect 2409 15991 2467 15997
rect 2424 15892 2452 15991
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 6236 16000 6377 16028
rect 6236 15988 6242 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 12526 16028 12532 16040
rect 12487 16000 12532 16028
rect 6365 15991 6423 15997
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 13722 15988 13728 16040
rect 13780 16028 13786 16040
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 13780 16000 14381 16028
rect 13780 15988 13786 16000
rect 14369 15997 14381 16000
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 16028 20775 16031
rect 21082 16028 21088 16040
rect 20763 16000 21088 16028
rect 20763 15997 20775 16000
rect 20717 15991 20775 15997
rect 15749 15963 15807 15969
rect 15749 15929 15761 15963
rect 15795 15960 15807 15963
rect 19426 15960 19432 15972
rect 15795 15932 19432 15960
rect 15795 15929 15807 15932
rect 15749 15923 15807 15929
rect 19426 15920 19432 15932
rect 19484 15960 19490 15972
rect 20548 15960 20576 15991
rect 21082 15988 21088 16000
rect 21140 15988 21146 16040
rect 19484 15932 20576 15960
rect 19484 15920 19490 15932
rect 2774 15892 2780 15904
rect 2424 15864 2780 15892
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 3789 15895 3847 15901
rect 3789 15861 3801 15895
rect 3835 15892 3847 15895
rect 3970 15892 3976 15904
rect 3835 15864 3976 15892
rect 3835 15861 3847 15864
rect 3789 15855 3847 15861
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 10597 15895 10655 15901
rect 10597 15861 10609 15895
rect 10643 15892 10655 15895
rect 11974 15892 11980 15904
rect 10643 15864 11980 15892
rect 10643 15861 10655 15864
rect 10597 15855 10655 15861
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 10689 15691 10747 15697
rect 10689 15657 10701 15691
rect 10735 15688 10747 15691
rect 13354 15688 13360 15700
rect 10735 15660 13360 15688
rect 10735 15657 10747 15660
rect 10689 15651 10747 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 19334 15580 19340 15632
rect 19392 15620 19398 15632
rect 21729 15623 21787 15629
rect 21729 15620 21741 15623
rect 19392 15592 21741 15620
rect 19392 15580 19398 15592
rect 8938 15512 8944 15564
rect 8996 15552 9002 15564
rect 9306 15552 9312 15564
rect 8996 15524 9312 15552
rect 8996 15512 9002 15524
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 21008 15561 21036 15592
rect 21729 15589 21741 15592
rect 21775 15620 21787 15623
rect 29362 15620 29368 15632
rect 21775 15592 29368 15620
rect 21775 15589 21787 15592
rect 21729 15583 21787 15589
rect 29362 15580 29368 15592
rect 29420 15580 29426 15632
rect 19889 15555 19947 15561
rect 19889 15521 19901 15555
rect 19935 15552 19947 15555
rect 20993 15555 21051 15561
rect 19935 15524 20116 15552
rect 19935 15521 19947 15524
rect 19889 15515 19947 15521
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15484 1915 15487
rect 3786 15484 3792 15496
rect 1903 15456 2820 15484
rect 3747 15456 3792 15484
rect 1903 15453 1915 15456
rect 1857 15447 1915 15453
rect 2792 15428 2820 15456
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 4056 15487 4114 15493
rect 4056 15453 4068 15487
rect 4102 15484 4114 15487
rect 4614 15484 4620 15496
rect 4102 15456 4620 15484
rect 4102 15453 4114 15456
rect 4056 15447 4114 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 6178 15484 6184 15496
rect 6139 15456 6184 15484
rect 6178 15444 6184 15456
rect 6236 15444 6242 15496
rect 6448 15487 6506 15493
rect 6448 15453 6460 15487
rect 6494 15484 6506 15487
rect 6730 15484 6736 15496
rect 6494 15456 6736 15484
rect 6494 15453 6506 15456
rect 6448 15447 6506 15453
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 9324 15484 9352 15512
rect 12161 15487 12219 15493
rect 12161 15484 12173 15487
rect 9324 15456 12173 15484
rect 12161 15453 12173 15456
rect 12207 15484 12219 15487
rect 13722 15484 13728 15496
rect 12207 15456 13728 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 12544 15428 12572 15456
rect 13722 15444 13728 15456
rect 13780 15484 13786 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 13780 15456 14289 15484
rect 13780 15444 13786 15456
rect 14277 15453 14289 15456
rect 14323 15484 14335 15487
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 14323 15456 16129 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 16117 15447 16175 15453
rect 16316 15456 18705 15484
rect 2124 15419 2182 15425
rect 2124 15385 2136 15419
rect 2170 15416 2182 15419
rect 2170 15388 2728 15416
rect 2170 15385 2182 15388
rect 2124 15379 2182 15385
rect 2700 15348 2728 15388
rect 2774 15376 2780 15428
rect 2832 15376 2838 15428
rect 9582 15425 9588 15428
rect 9576 15379 9588 15425
rect 9640 15416 9646 15428
rect 12428 15419 12486 15425
rect 9640 15388 9676 15416
rect 9582 15376 9588 15379
rect 9640 15376 9646 15388
rect 12428 15385 12440 15419
rect 12474 15385 12486 15419
rect 12428 15379 12486 15385
rect 2866 15348 2872 15360
rect 2700 15320 2872 15348
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 3237 15351 3295 15357
rect 3237 15317 3249 15351
rect 3283 15348 3295 15351
rect 3326 15348 3332 15360
rect 3283 15320 3332 15348
rect 3283 15317 3295 15320
rect 3237 15311 3295 15317
rect 3326 15308 3332 15320
rect 3384 15308 3390 15360
rect 5166 15348 5172 15360
rect 5127 15320 5172 15348
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 7561 15351 7619 15357
rect 7561 15317 7573 15351
rect 7607 15348 7619 15351
rect 8110 15348 8116 15360
rect 7607 15320 8116 15348
rect 7607 15317 7619 15320
rect 7561 15311 7619 15317
rect 8110 15308 8116 15320
rect 8168 15348 8174 15360
rect 8386 15348 8392 15360
rect 8168 15320 8392 15348
rect 8168 15308 8174 15320
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 12452 15348 12480 15379
rect 12526 15376 12532 15428
rect 12584 15376 12590 15428
rect 14090 15416 14096 15428
rect 13464 15388 14096 15416
rect 13464 15348 13492 15388
rect 14090 15376 14096 15388
rect 14148 15376 14154 15428
rect 14544 15419 14602 15425
rect 14544 15385 14556 15419
rect 14590 15416 14602 15419
rect 16206 15416 16212 15428
rect 14590 15388 16212 15416
rect 14590 15385 14602 15388
rect 14544 15379 14602 15385
rect 16206 15376 16212 15388
rect 16264 15376 16270 15428
rect 12452 15320 13492 15348
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 15010 15348 15016 15360
rect 13587 15320 15016 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15657 15351 15715 15357
rect 15657 15317 15669 15351
rect 15703 15348 15715 15351
rect 16316 15348 16344 15456
rect 18693 15453 18705 15456
rect 18739 15484 18751 15487
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 18739 15456 19809 15484
rect 18739 15453 18751 15456
rect 18693 15447 18751 15453
rect 19797 15453 19809 15456
rect 19843 15484 19855 15487
rect 19978 15484 19984 15496
rect 19843 15456 19984 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20088 15484 20116 15524
rect 20993 15521 21005 15555
rect 21039 15521 21051 15555
rect 20993 15515 21051 15521
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21140 15524 21185 15552
rect 21140 15512 21146 15524
rect 20714 15484 20720 15496
rect 20088 15456 20720 15484
rect 20714 15444 20720 15456
rect 20772 15484 20778 15496
rect 21100 15484 21128 15512
rect 20772 15456 21128 15484
rect 20772 15444 20778 15456
rect 16384 15419 16442 15425
rect 16384 15385 16396 15419
rect 16430 15416 16442 15419
rect 17678 15416 17684 15428
rect 16430 15388 17684 15416
rect 16430 15385 16442 15388
rect 16384 15379 16442 15385
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 19705 15419 19763 15425
rect 19705 15385 19717 15419
rect 19751 15416 19763 15419
rect 20254 15416 20260 15428
rect 19751 15388 20260 15416
rect 19751 15385 19763 15388
rect 19705 15379 19763 15385
rect 20254 15376 20260 15388
rect 20312 15376 20318 15428
rect 20901 15419 20959 15425
rect 20901 15385 20913 15419
rect 20947 15416 20959 15419
rect 21542 15416 21548 15428
rect 20947 15388 21548 15416
rect 20947 15385 20959 15388
rect 20901 15379 20959 15385
rect 21542 15376 21548 15388
rect 21600 15376 21606 15428
rect 17494 15348 17500 15360
rect 15703 15320 16344 15348
rect 17455 15320 17500 15348
rect 15703 15317 15715 15320
rect 15657 15311 15715 15317
rect 17494 15308 17500 15320
rect 17552 15308 17558 15360
rect 18690 15308 18696 15360
rect 18748 15348 18754 15360
rect 19337 15351 19395 15357
rect 19337 15348 19349 15351
rect 18748 15320 19349 15348
rect 18748 15308 18754 15320
rect 19337 15317 19349 15320
rect 19383 15317 19395 15351
rect 20530 15348 20536 15360
rect 20491 15320 20536 15348
rect 19337 15311 19395 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 22278 15308 22284 15360
rect 22336 15348 22342 15360
rect 22373 15351 22431 15357
rect 22373 15348 22385 15351
rect 22336 15320 22385 15348
rect 22336 15308 22342 15320
rect 22373 15317 22385 15320
rect 22419 15348 22431 15351
rect 31478 15348 31484 15360
rect 22419 15320 31484 15348
rect 22419 15317 22431 15320
rect 22373 15311 22431 15317
rect 31478 15308 31484 15320
rect 31536 15308 31542 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 2774 15104 2780 15156
rect 2832 15104 2838 15156
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 6604 15116 6684 15144
rect 6604 15104 6610 15116
rect 2792 15076 2820 15104
rect 3786 15076 3792 15088
rect 2516 15048 3792 15076
rect 2516 15017 2544 15048
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 6656 15085 6684 15116
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 18046 15144 18052 15156
rect 9548 15116 9628 15144
rect 18007 15116 18052 15144
rect 9548 15104 9554 15116
rect 9600 15085 9628 15116
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 18693 15147 18751 15153
rect 18693 15113 18705 15147
rect 18739 15113 18751 15147
rect 21821 15147 21879 15153
rect 21821 15144 21833 15147
rect 18693 15107 18751 15113
rect 18800 15116 21833 15144
rect 6632 15079 6690 15085
rect 6632 15045 6644 15079
rect 6678 15045 6690 15079
rect 6632 15039 6690 15045
rect 9576 15079 9634 15085
rect 9576 15045 9588 15079
rect 9622 15045 9634 15079
rect 9576 15039 9634 15045
rect 14636 15079 14694 15085
rect 14636 15045 14648 15079
rect 14682 15076 14694 15079
rect 18708 15076 18736 15107
rect 14682 15048 18736 15076
rect 14682 15045 14694 15048
rect 14636 15039 14694 15045
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2768 15011 2826 15017
rect 2768 14977 2780 15011
rect 2814 15008 2826 15011
rect 3234 15008 3240 15020
rect 2814 14980 3240 15008
rect 2814 14977 2826 14980
rect 2768 14971 2826 14977
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 9306 15008 9312 15020
rect 9267 14980 9312 15008
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 12796 15011 12854 15017
rect 12796 14977 12808 15011
rect 12842 15008 12854 15011
rect 15102 15008 15108 15020
rect 12842 14980 15108 15008
rect 12842 14977 12854 14980
rect 12796 14971 12854 14977
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 15008 18291 15011
rect 18800 15008 18828 15116
rect 21821 15113 21833 15116
rect 21867 15113 21879 15147
rect 22278 15144 22284 15156
rect 22239 15116 22284 15144
rect 21821 15107 21879 15113
rect 22278 15104 22284 15116
rect 22336 15104 22342 15156
rect 19797 15079 19855 15085
rect 19797 15076 19809 15079
rect 19260 15048 19809 15076
rect 18279 14980 18828 15008
rect 18877 15011 18935 15017
rect 18279 14977 18291 14980
rect 18233 14971 18291 14977
rect 18877 14977 18889 15011
rect 18923 15008 18935 15011
rect 19150 15008 19156 15020
rect 18923 14980 19156 15008
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 19150 14968 19156 14980
rect 19208 14968 19214 15020
rect 6178 14900 6184 14952
rect 6236 14940 6242 14952
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 6236 14912 6377 14940
rect 6236 14900 6242 14912
rect 6365 14909 6377 14912
rect 6411 14909 6423 14943
rect 12526 14940 12532 14952
rect 12487 14912 12532 14940
rect 6365 14903 6423 14909
rect 3878 14804 3884 14816
rect 3839 14776 3884 14804
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 6380 14804 6408 14903
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 13722 14900 13728 14952
rect 13780 14940 13786 14952
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 13780 14912 14381 14940
rect 13780 14900 13786 14912
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 17494 14900 17500 14952
rect 17552 14940 17558 14952
rect 17589 14943 17647 14949
rect 17589 14940 17601 14943
rect 17552 14912 17601 14940
rect 17552 14900 17558 14912
rect 17589 14909 17601 14912
rect 17635 14940 17647 14943
rect 19260 14940 19288 15048
rect 19797 15045 19809 15048
rect 19843 15076 19855 15079
rect 30374 15076 30380 15088
rect 19843 15048 30380 15076
rect 19843 15045 19855 15048
rect 19797 15039 19855 15045
rect 30374 15036 30380 15048
rect 30432 15036 30438 15088
rect 19705 15011 19763 15017
rect 19705 14977 19717 15011
rect 19751 15008 19763 15011
rect 19978 15008 19984 15020
rect 19751 14980 19984 15008
rect 19751 14977 19763 14980
rect 19705 14971 19763 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 20947 14980 21496 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 17635 14912 19288 14940
rect 19889 14943 19947 14949
rect 17635 14909 17647 14912
rect 17589 14903 17647 14909
rect 19889 14909 19901 14943
rect 19935 14940 19947 14943
rect 20714 14940 20720 14952
rect 19935 14912 20720 14940
rect 19935 14909 19947 14912
rect 19889 14903 19947 14909
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 20806 14900 20812 14952
rect 20864 14940 20870 14952
rect 20993 14943 21051 14949
rect 20993 14940 21005 14943
rect 20864 14912 21005 14940
rect 20864 14900 20870 14912
rect 20993 14909 21005 14912
rect 21039 14909 21051 14943
rect 20993 14903 21051 14909
rect 21082 14900 21088 14952
rect 21140 14940 21146 14952
rect 21468 14940 21496 14980
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 21968 14980 22201 15008
rect 21968 14968 21974 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 21140 14912 21185 14940
rect 21468 14912 22324 14940
rect 21140 14900 21146 14912
rect 22002 14872 22008 14884
rect 15580 14844 22008 14872
rect 6730 14804 6736 14816
rect 6380 14776 6736 14804
rect 6730 14764 6736 14776
rect 6788 14764 6794 14816
rect 7745 14807 7803 14813
rect 7745 14773 7757 14807
rect 7791 14804 7803 14807
rect 8294 14804 8300 14816
rect 7791 14776 8300 14804
rect 7791 14773 7803 14776
rect 7745 14767 7803 14773
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 13630 14804 13636 14816
rect 10735 14776 13636 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 15010 14764 15016 14816
rect 15068 14804 15074 14816
rect 15580 14804 15608 14844
rect 22002 14832 22008 14844
rect 22060 14832 22066 14884
rect 22296 14872 22324 14912
rect 22370 14900 22376 14952
rect 22428 14940 22434 14952
rect 22428 14912 22473 14940
rect 22428 14900 22434 14912
rect 24394 14872 24400 14884
rect 22296 14844 24400 14872
rect 24394 14832 24400 14844
rect 24452 14832 24458 14884
rect 15746 14804 15752 14816
rect 15068 14776 15608 14804
rect 15707 14776 15752 14804
rect 15068 14764 15074 14776
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 19242 14764 19248 14816
rect 19300 14804 19306 14816
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 19300 14776 19349 14804
rect 19300 14764 19306 14776
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 19337 14767 19395 14773
rect 20070 14764 20076 14816
rect 20128 14804 20134 14816
rect 20533 14807 20591 14813
rect 20533 14804 20545 14807
rect 20128 14776 20545 14804
rect 20128 14764 20134 14776
rect 20533 14773 20545 14776
rect 20579 14773 20591 14807
rect 20533 14767 20591 14773
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 23014 14804 23020 14816
rect 20864 14776 23020 14804
rect 20864 14764 20870 14776
rect 23014 14764 23020 14776
rect 23072 14764 23078 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 13998 14600 14004 14612
rect 3936 14572 14004 14600
rect 3936 14560 3942 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14090 14560 14096 14612
rect 14148 14600 14154 14612
rect 14148 14572 15884 14600
rect 14148 14560 14154 14572
rect 15856 14532 15884 14572
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 16264 14572 18521 14600
rect 16264 14560 16270 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 19208 14572 20545 14600
rect 19208 14560 19214 14572
rect 20533 14569 20545 14572
rect 20579 14569 20591 14603
rect 20533 14563 20591 14569
rect 19245 14535 19303 14541
rect 19245 14532 19257 14535
rect 15856 14504 19257 14532
rect 19245 14501 19257 14504
rect 19291 14501 19303 14535
rect 21729 14535 21787 14541
rect 21729 14532 21741 14535
rect 19245 14495 19303 14501
rect 19444 14504 21741 14532
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 3844 14436 5488 14464
rect 3844 14424 3850 14436
rect 5460 14405 5488 14436
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 13722 14464 13728 14476
rect 12584 14436 13728 14464
rect 12584 14424 12590 14436
rect 13722 14424 13728 14436
rect 13780 14464 13786 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 13780 14436 14105 14464
rect 13780 14424 13786 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 6178 14396 6184 14408
rect 5491 14368 6184 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 4632 14328 4660 14359
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 14366 14405 14372 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 9364 14368 10425 14396
rect 9364 14356 9370 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 14360 14396 14372 14405
rect 14327 14368 14372 14396
rect 10413 14359 10471 14365
rect 14360 14359 14372 14368
rect 14366 14356 14372 14359
rect 14424 14356 14430 14408
rect 18690 14396 18696 14408
rect 18651 14368 18696 14396
rect 18690 14356 18696 14368
rect 18748 14356 18754 14408
rect 19444 14405 19472 14504
rect 21729 14501 21741 14504
rect 21775 14501 21787 14535
rect 21729 14495 21787 14501
rect 20990 14464 20996 14476
rect 20951 14436 20996 14464
rect 20990 14424 20996 14436
rect 21048 14424 21054 14476
rect 21082 14424 21088 14476
rect 21140 14464 21146 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 21140 14436 22293 14464
rect 21140 14424 21146 14436
rect 22281 14433 22293 14436
rect 22327 14464 22339 14467
rect 22370 14464 22376 14476
rect 22327 14436 22376 14464
rect 22327 14433 22339 14436
rect 22281 14427 22339 14433
rect 22370 14424 22376 14436
rect 22428 14424 22434 14476
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 20070 14396 20076 14408
rect 20031 14368 20076 14396
rect 19429 14359 19487 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 21008 14396 21036 14424
rect 28166 14396 28172 14408
rect 21008 14368 28172 14396
rect 28166 14356 28172 14368
rect 28224 14356 28230 14408
rect 5534 14328 5540 14340
rect 4632 14300 5540 14328
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 5718 14337 5724 14340
rect 5712 14291 5724 14337
rect 5776 14328 5782 14340
rect 10134 14328 10140 14340
rect 10192 14337 10198 14340
rect 5776 14300 5812 14328
rect 10104 14300 10140 14328
rect 5718 14288 5724 14291
rect 5776 14288 5782 14300
rect 10134 14288 10140 14300
rect 10192 14291 10204 14337
rect 10192 14288 10198 14291
rect 13906 14288 13912 14340
rect 13964 14328 13970 14340
rect 20714 14328 20720 14340
rect 13964 14300 20720 14328
rect 13964 14288 13970 14300
rect 20714 14288 20720 14300
rect 20772 14288 20778 14340
rect 20901 14331 20959 14337
rect 20901 14297 20913 14331
rect 20947 14328 20959 14331
rect 21634 14328 21640 14340
rect 20947 14300 21640 14328
rect 20947 14297 20959 14300
rect 20901 14291 20959 14297
rect 21634 14288 21640 14300
rect 21692 14288 21698 14340
rect 22097 14331 22155 14337
rect 22097 14297 22109 14331
rect 22143 14328 22155 14331
rect 24118 14328 24124 14340
rect 22143 14300 24124 14328
rect 22143 14297 22155 14300
rect 22097 14291 22155 14297
rect 24118 14288 24124 14300
rect 24176 14288 24182 14340
rect 4430 14260 4436 14272
rect 4391 14232 4436 14260
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 6822 14260 6828 14272
rect 6783 14232 6828 14260
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 9033 14263 9091 14269
rect 9033 14229 9045 14263
rect 9079 14260 9091 14263
rect 10410 14260 10416 14272
rect 9079 14232 10416 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 10410 14220 10416 14232
rect 10468 14260 10474 14272
rect 10594 14260 10600 14272
rect 10468 14232 10600 14260
rect 10468 14220 10474 14232
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14260 15531 14263
rect 16482 14260 16488 14272
rect 15519 14232 16488 14260
rect 15519 14229 15531 14232
rect 15473 14223 15531 14229
rect 16482 14220 16488 14232
rect 16540 14220 16546 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19392 14232 19901 14260
rect 19392 14220 19398 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 19889 14223 19947 14229
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22186 14260 22192 14272
rect 22060 14232 22192 14260
rect 22060 14220 22066 14232
rect 22186 14220 22192 14232
rect 22244 14260 22250 14272
rect 24302 14260 24308 14272
rect 22244 14232 24308 14260
rect 22244 14220 22250 14232
rect 24302 14220 24308 14232
rect 24360 14220 24366 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 10502 14056 10508 14068
rect 6880 14028 10508 14056
rect 6880 14016 6886 14028
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 17678 14016 17684 14068
rect 17736 14056 17742 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 17736 14028 19073 14056
rect 17736 14016 17742 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 19426 14016 19432 14068
rect 19484 14056 19490 14068
rect 19705 14059 19763 14065
rect 19705 14056 19717 14059
rect 19484 14028 19717 14056
rect 19484 14016 19490 14028
rect 19705 14025 19717 14028
rect 19751 14025 19763 14059
rect 19705 14019 19763 14025
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 20993 14059 21051 14065
rect 20993 14056 21005 14059
rect 20772 14028 21005 14056
rect 20772 14016 20778 14028
rect 20993 14025 21005 14028
rect 21039 14056 21051 14059
rect 21174 14056 21180 14068
rect 21039 14028 21180 14056
rect 21039 14025 21051 14028
rect 20993 14019 21051 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 21913 14059 21971 14065
rect 21913 14025 21925 14059
rect 21959 14056 21971 14059
rect 22186 14056 22192 14068
rect 21959 14028 22192 14056
rect 21959 14025 21971 14028
rect 21913 14019 21971 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 3544 13991 3602 13997
rect 3544 13957 3556 13991
rect 3590 13988 3602 13991
rect 4430 13988 4436 14000
rect 3590 13960 4436 13988
rect 3590 13957 3602 13960
rect 3544 13951 3602 13957
rect 4430 13948 4436 13960
rect 4488 13948 4494 14000
rect 14636 13991 14694 13997
rect 14636 13957 14648 13991
rect 14682 13988 14694 13991
rect 19334 13988 19340 14000
rect 14682 13960 19340 13988
rect 14682 13957 14694 13960
rect 14636 13951 14694 13957
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 21192 13988 21220 14016
rect 25130 13988 25136 14000
rect 21192 13960 25136 13988
rect 25130 13948 25136 13960
rect 25188 13948 25194 14000
rect 3786 13920 3792 13932
rect 3747 13892 3792 13920
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 8588 13892 9137 13920
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8588 13861 8616 13892
rect 9125 13889 9137 13892
rect 9171 13889 9183 13923
rect 9125 13883 9183 13889
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 13780 13892 14381 13920
rect 13780 13880 13786 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 19242 13920 19248 13932
rect 19203 13892 19248 13920
rect 14369 13883 14427 13889
rect 19242 13880 19248 13892
rect 19300 13880 19306 13932
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20530 13920 20536 13932
rect 19935 13892 20536 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 20901 13923 20959 13929
rect 20901 13889 20913 13923
rect 20947 13920 20959 13923
rect 22370 13920 22376 13932
rect 20947 13892 22376 13920
rect 20947 13889 20959 13892
rect 20901 13883 20959 13889
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8260 13824 8585 13852
rect 8260 13812 8266 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 20806 13852 20812 13864
rect 8573 13815 8631 13821
rect 15764 13824 20812 13852
rect 15764 13793 15792 13824
rect 20806 13812 20812 13824
rect 20864 13812 20870 13864
rect 21082 13852 21088 13864
rect 20995 13824 21088 13852
rect 21082 13812 21088 13824
rect 21140 13812 21146 13864
rect 15749 13787 15807 13793
rect 15749 13753 15761 13787
rect 15795 13753 15807 13787
rect 15749 13747 15807 13753
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 21100 13784 21128 13812
rect 20956 13756 21128 13784
rect 20956 13744 20962 13756
rect 10410 13716 10416 13728
rect 10371 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 19518 13716 19524 13728
rect 13688 13688 19524 13716
rect 13688 13676 13694 13688
rect 19518 13676 19524 13688
rect 19576 13676 19582 13728
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20533 13719 20591 13725
rect 20533 13716 20545 13719
rect 20220 13688 20545 13716
rect 20220 13676 20226 13688
rect 20533 13685 20545 13688
rect 20579 13685 20591 13719
rect 20533 13679 20591 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 15102 13472 15108 13524
rect 15160 13512 15166 13524
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 15160 13484 19993 13512
rect 15160 13472 15166 13484
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 19981 13475 20039 13481
rect 20717 13515 20775 13521
rect 20717 13481 20729 13515
rect 20763 13512 20775 13515
rect 20990 13512 20996 13524
rect 20763 13484 20996 13512
rect 20763 13481 20775 13484
rect 20717 13475 20775 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 21174 13512 21180 13524
rect 21135 13484 21180 13512
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 10318 13404 10324 13456
rect 10376 13444 10382 13456
rect 10376 13416 12940 13444
rect 10376 13404 10382 13416
rect 12161 13379 12219 13385
rect 12161 13345 12173 13379
rect 12207 13376 12219 13379
rect 12526 13376 12532 13388
rect 12207 13348 12532 13376
rect 12207 13345 12219 13348
rect 12161 13339 12219 13345
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 12912 13376 12940 13416
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 19426 13444 19432 13456
rect 14056 13416 19432 13444
rect 14056 13404 14062 13416
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 19518 13404 19524 13456
rect 19576 13444 19582 13456
rect 25130 13444 25136 13456
rect 19576 13416 25136 13444
rect 19576 13404 19582 13416
rect 25130 13404 25136 13416
rect 25188 13404 25194 13456
rect 23474 13376 23480 13388
rect 12912 13348 23480 13376
rect 23474 13336 23480 13348
rect 23532 13336 23538 13388
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 11422 13308 11428 13320
rect 11112 13280 11428 13308
rect 11112 13268 11118 13280
rect 11422 13268 11428 13280
rect 11480 13308 11486 13320
rect 17218 13308 17224 13320
rect 11480 13280 17224 13308
rect 11480 13268 11486 13280
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 20162 13308 20168 13320
rect 20123 13280 20168 13308
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 5258 13240 5264 13252
rect 5219 13212 5264 13240
rect 5258 13200 5264 13212
rect 5316 13240 5322 13252
rect 10410 13240 10416 13252
rect 5316 13212 10416 13240
rect 5316 13200 5322 13212
rect 10410 13200 10416 13212
rect 10468 13200 10474 13252
rect 13538 13200 13544 13252
rect 13596 13240 13602 13252
rect 27614 13240 27620 13252
rect 13596 13212 27620 13240
rect 13596 13200 13602 13212
rect 27614 13200 27620 13212
rect 27672 13200 27678 13252
rect 6730 13172 6736 13184
rect 6691 13144 6736 13172
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 10321 12971 10379 12977
rect 10321 12937 10333 12971
rect 10367 12968 10379 12971
rect 11054 12968 11060 12980
rect 10367 12940 11060 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 17218 12928 17224 12980
rect 17276 12968 17282 12980
rect 25590 12968 25596 12980
rect 17276 12940 25596 12968
rect 17276 12928 17282 12940
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 2866 12900 2872 12912
rect 2424 12872 2872 12900
rect 2424 12841 2452 12872
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 9214 12909 9220 12912
rect 9208 12900 9220 12909
rect 6788 12872 8984 12900
rect 9175 12872 9220 12900
rect 6788 12860 6794 12872
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 2676 12835 2734 12841
rect 2676 12801 2688 12835
rect 2722 12832 2734 12835
rect 2958 12832 2964 12844
rect 2722 12804 2964 12832
rect 2722 12801 2734 12804
rect 2676 12795 2734 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 7368 12835 7426 12841
rect 7368 12801 7380 12835
rect 7414 12832 7426 12835
rect 8846 12832 8852 12844
rect 7414 12804 8852 12832
rect 7414 12801 7426 12804
rect 7368 12795 7426 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 8956 12841 8984 12872
rect 9208 12863 9220 12872
rect 9214 12860 9220 12863
rect 9272 12860 9278 12912
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 14636 12835 14694 12841
rect 14636 12801 14648 12835
rect 14682 12832 14694 12835
rect 15562 12832 15568 12844
rect 14682 12804 15568 12832
rect 14682 12801 14694 12804
rect 14636 12795 14694 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 7098 12764 7104 12776
rect 7059 12736 7104 12764
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14332 12736 14381 12764
rect 14332 12724 14338 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3789 12631 3847 12637
rect 3789 12628 3801 12631
rect 3200 12600 3801 12628
rect 3200 12588 3206 12600
rect 3789 12597 3801 12600
rect 3835 12597 3847 12631
rect 3789 12591 3847 12597
rect 8481 12631 8539 12637
rect 8481 12597 8493 12631
rect 8527 12628 8539 12631
rect 9950 12628 9956 12640
rect 8527 12600 9956 12628
rect 8527 12597 8539 12600
rect 8481 12591 8539 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 15749 12631 15807 12637
rect 15749 12597 15761 12631
rect 15795 12628 15807 12631
rect 19334 12628 19340 12640
rect 15795 12600 19340 12628
rect 15795 12597 15807 12600
rect 15749 12591 15807 12597
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 8110 12384 8116 12436
rect 8168 12424 8174 12436
rect 8168 12396 15516 12424
rect 8168 12384 8174 12396
rect 15488 12356 15516 12396
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 19613 12427 19671 12433
rect 19613 12424 19625 12427
rect 15620 12396 19625 12424
rect 15620 12384 15626 12396
rect 19613 12393 19625 12396
rect 19659 12393 19671 12427
rect 19613 12387 19671 12393
rect 20625 12427 20683 12433
rect 20625 12393 20637 12427
rect 20671 12424 20683 12427
rect 20898 12424 20904 12436
rect 20671 12396 20904 12424
rect 20671 12393 20683 12396
rect 20625 12387 20683 12393
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 16298 12356 16304 12368
rect 15488 12328 16304 12356
rect 16298 12316 16304 12328
rect 16356 12316 16362 12368
rect 20070 12248 20076 12300
rect 20128 12288 20134 12300
rect 20128 12260 20760 12288
rect 20128 12248 20134 12260
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 2866 12220 2872 12232
rect 1903 12192 2872 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 6273 12223 6331 12229
rect 6273 12189 6285 12223
rect 6319 12220 6331 12223
rect 7098 12220 7104 12232
rect 6319 12192 7104 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 10042 12220 10048 12232
rect 10003 12192 10048 12220
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 14274 12220 14280 12232
rect 14235 12192 14280 12220
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12220 19855 12223
rect 20346 12220 20352 12232
rect 19843 12192 20352 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 20346 12180 20352 12192
rect 20404 12180 20410 12232
rect 20732 12229 20760 12260
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12189 20775 12223
rect 20717 12183 20775 12189
rect 2124 12155 2182 12161
rect 2124 12121 2136 12155
rect 2170 12152 2182 12155
rect 2406 12152 2412 12164
rect 2170 12124 2412 12152
rect 2170 12121 2182 12124
rect 2124 12115 2182 12121
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 6540 12155 6598 12161
rect 6540 12121 6552 12155
rect 6586 12152 6598 12155
rect 7282 12152 7288 12164
rect 6586 12124 7288 12152
rect 6586 12121 6598 12124
rect 6540 12115 6598 12121
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 10312 12155 10370 12161
rect 10312 12121 10324 12155
rect 10358 12152 10370 12155
rect 11330 12152 11336 12164
rect 10358 12124 11336 12152
rect 10358 12121 10370 12124
rect 10312 12115 10370 12121
rect 11330 12112 11336 12124
rect 11388 12112 11394 12164
rect 14544 12155 14602 12161
rect 14544 12121 14556 12155
rect 14590 12152 14602 12155
rect 18782 12152 18788 12164
rect 14590 12124 18788 12152
rect 14590 12121 14602 12124
rect 14544 12115 14602 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 19978 12112 19984 12164
rect 20036 12152 20042 12164
rect 20622 12152 20628 12164
rect 20036 12124 20628 12152
rect 20036 12112 20042 12124
rect 20622 12112 20628 12124
rect 20680 12112 20686 12164
rect 3234 12084 3240 12096
rect 3195 12056 3240 12084
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 7653 12087 7711 12093
rect 7653 12053 7665 12087
rect 7699 12084 7711 12087
rect 10226 12084 10232 12096
rect 7699 12056 10232 12084
rect 7699 12053 7711 12056
rect 7653 12047 7711 12053
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 11425 12087 11483 12093
rect 11425 12053 11437 12087
rect 11471 12084 11483 12087
rect 12066 12084 12072 12096
rect 11471 12056 12072 12084
rect 11471 12053 11483 12056
rect 11425 12047 11483 12053
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 15657 12087 15715 12093
rect 15657 12053 15669 12087
rect 15703 12084 15715 12087
rect 20162 12084 20168 12096
rect 15703 12056 20168 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 20162 12044 20168 12056
rect 20220 12044 20226 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 16206 11880 16212 11892
rect 5224 11852 16212 11880
rect 5224 11840 5230 11852
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17862 11840 17868 11892
rect 17920 11840 17926 11892
rect 18782 11880 18788 11892
rect 18743 11852 18788 11880
rect 18782 11840 18788 11852
rect 18840 11840 18846 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19794 11880 19800 11892
rect 19392 11852 19800 11880
rect 19392 11840 19398 11852
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 20346 11880 20352 11892
rect 20307 11852 20352 11880
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 28994 11880 29000 11892
rect 20456 11852 29000 11880
rect 7098 11812 7104 11824
rect 2884 11784 7104 11812
rect 2884 11756 2912 11784
rect 2866 11744 2872 11756
rect 2779 11716 2872 11744
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 3136 11747 3194 11753
rect 3136 11713 3148 11747
rect 3182 11744 3194 11747
rect 4706 11744 4712 11756
rect 3182 11716 4712 11744
rect 3182 11713 3194 11716
rect 3136 11707 3194 11713
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 6380 11753 6408 11784
rect 7098 11772 7104 11784
rect 7156 11772 7162 11824
rect 9760 11815 9818 11821
rect 9760 11781 9772 11815
rect 9806 11812 9818 11815
rect 13998 11812 14004 11824
rect 9806 11784 14004 11812
rect 9806 11781 9818 11784
rect 9760 11775 9818 11781
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 17880 11812 17908 11840
rect 20456 11812 20484 11852
rect 28994 11840 29000 11852
rect 29052 11840 29058 11892
rect 37366 11812 37372 11824
rect 17880 11784 20484 11812
rect 31726 11784 37372 11812
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6632 11747 6690 11753
rect 6632 11713 6644 11747
rect 6678 11744 6690 11747
rect 7834 11744 7840 11756
rect 6678 11716 7840 11744
rect 6678 11713 6690 11716
rect 6632 11707 6690 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 10042 11744 10048 11756
rect 9508 11716 10048 11744
rect 9508 11685 9536 11716
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 14544 11747 14602 11753
rect 14544 11713 14556 11747
rect 14590 11744 14602 11747
rect 17862 11744 17868 11756
rect 14590 11716 17868 11744
rect 14590 11713 14602 11716
rect 14544 11707 14602 11713
rect 17862 11704 17868 11716
rect 17920 11704 17926 11756
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11744 19027 11747
rect 19978 11744 19984 11756
rect 19015 11716 19984 11744
rect 19015 11713 19027 11716
rect 18969 11707 19027 11713
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 20990 11744 20996 11756
rect 20763 11716 20996 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11645 9551 11679
rect 14274 11676 14280 11688
rect 14235 11648 14280 11676
rect 9493 11639 9551 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 19794 11636 19800 11688
rect 19852 11676 19858 11688
rect 20809 11679 20867 11685
rect 20809 11676 20821 11679
rect 19852 11648 20821 11676
rect 19852 11636 19858 11648
rect 20809 11645 20821 11648
rect 20855 11645 20867 11679
rect 20809 11639 20867 11645
rect 15657 11611 15715 11617
rect 15657 11577 15669 11611
rect 15703 11608 15715 11611
rect 20714 11608 20720 11620
rect 15703 11580 20720 11608
rect 15703 11577 15715 11580
rect 15657 11571 15715 11577
rect 20714 11568 20720 11580
rect 20772 11568 20778 11620
rect 20824 11608 20852 11639
rect 20898 11636 20904 11688
rect 20956 11676 20962 11688
rect 20956 11648 21001 11676
rect 20956 11636 20962 11648
rect 26142 11608 26148 11620
rect 20824 11580 26148 11608
rect 26142 11568 26148 11580
rect 26200 11568 26206 11620
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 4798 11540 4804 11552
rect 4295 11512 4804 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 7742 11540 7748 11552
rect 7703 11512 7748 11540
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 10873 11543 10931 11549
rect 10873 11509 10885 11543
rect 10919 11540 10931 11543
rect 11698 11540 11704 11552
rect 10919 11512 11704 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 18230 11540 18236 11552
rect 18191 11512 18236 11540
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 18322 11500 18328 11552
rect 18380 11540 18386 11552
rect 19150 11540 19156 11552
rect 18380 11512 19156 11540
rect 18380 11500 18386 11512
rect 19150 11500 19156 11512
rect 19208 11540 19214 11552
rect 31726 11540 31754 11784
rect 37366 11772 37372 11784
rect 37424 11772 37430 11824
rect 19208 11512 31754 11540
rect 19208 11500 19214 11512
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11336 5227 11339
rect 7374 11336 7380 11348
rect 5215 11308 7380 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 8389 11339 8447 11345
rect 8389 11305 8401 11339
rect 8435 11336 8447 11339
rect 10318 11336 10324 11348
rect 8435 11308 10324 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 19242 11336 19248 11348
rect 15703 11308 19248 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 19242 11296 19248 11308
rect 19300 11296 19306 11348
rect 20162 11296 20168 11348
rect 20220 11336 20226 11348
rect 20441 11339 20499 11345
rect 20441 11336 20453 11339
rect 20220 11308 20453 11336
rect 20220 11296 20226 11308
rect 20441 11305 20453 11308
rect 20487 11305 20499 11339
rect 20441 11299 20499 11305
rect 3237 11271 3295 11277
rect 3237 11237 3249 11271
rect 3283 11268 3295 11271
rect 3602 11268 3608 11280
rect 3283 11240 3608 11268
rect 3283 11237 3295 11240
rect 3237 11231 3295 11237
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 13722 11268 13728 11280
rect 11471 11240 13728 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 17589 11271 17647 11277
rect 17589 11237 17601 11271
rect 17635 11268 17647 11271
rect 18322 11268 18328 11280
rect 17635 11240 18328 11268
rect 17635 11237 17647 11240
rect 17589 11231 17647 11237
rect 18322 11228 18328 11240
rect 18380 11228 18386 11280
rect 18509 11271 18567 11277
rect 18509 11237 18521 11271
rect 18555 11237 18567 11271
rect 18509 11231 18567 11237
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 1857 11135 1915 11141
rect 1857 11101 1869 11135
rect 1903 11132 1915 11135
rect 2866 11132 2872 11144
rect 1903 11104 2872 11132
rect 1903 11101 1915 11104
rect 1857 11095 1915 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 6549 11135 6607 11141
rect 6549 11101 6561 11135
rect 6595 11132 6607 11135
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6595 11104 7021 11132
rect 6595 11101 6607 11104
rect 6549 11095 6607 11101
rect 7009 11101 7021 11104
rect 7055 11132 7067 11135
rect 7098 11132 7104 11144
rect 7055 11104 7104 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11132 14338 11144
rect 16209 11135 16267 11141
rect 16209 11132 16221 11135
rect 14332 11104 16221 11132
rect 14332 11092 14338 11104
rect 16209 11101 16221 11104
rect 16255 11101 16267 11135
rect 18524 11132 18552 11231
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11200 19947 11203
rect 20070 11200 20076 11212
rect 19935 11172 20076 11200
rect 19935 11169 19947 11172
rect 19889 11163 19947 11169
rect 20070 11160 20076 11172
rect 20128 11160 20134 11212
rect 18690 11132 18696 11144
rect 16209 11095 16267 11101
rect 16408 11104 18552 11132
rect 18651 11104 18696 11132
rect 2124 11067 2182 11073
rect 2124 11033 2136 11067
rect 2170 11064 2182 11067
rect 2682 11064 2688 11076
rect 2170 11036 2688 11064
rect 2170 11033 2182 11036
rect 2124 11027 2182 11033
rect 2682 11024 2688 11036
rect 2740 11024 2746 11076
rect 6270 11064 6276 11076
rect 6328 11073 6334 11076
rect 6240 11036 6276 11064
rect 6270 11024 6276 11036
rect 6328 11027 6340 11073
rect 7276 11067 7334 11073
rect 7276 11033 7288 11067
rect 7322 11064 7334 11067
rect 8754 11064 8760 11076
rect 7322 11036 8760 11064
rect 7322 11033 7334 11036
rect 7276 11027 7334 11033
rect 6328 11024 6334 11027
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 10312 11067 10370 11073
rect 10312 11033 10324 11067
rect 10358 11064 10370 11067
rect 10778 11064 10784 11076
rect 10358 11036 10784 11064
rect 10358 11033 10370 11036
rect 10312 11027 10370 11033
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 14544 11067 14602 11073
rect 14544 11033 14556 11067
rect 14590 11064 14602 11067
rect 16408 11064 16436 11104
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 18840 11104 19625 11132
rect 18840 11092 18846 11104
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 34790 11132 34796 11144
rect 19613 11095 19671 11101
rect 19720 11104 34796 11132
rect 14590 11036 16436 11064
rect 16476 11067 16534 11073
rect 14590 11033 14602 11036
rect 14544 11027 14602 11033
rect 16476 11033 16488 11067
rect 16522 11064 16534 11067
rect 18138 11064 18144 11076
rect 16522 11036 18144 11064
rect 16522 11033 16534 11036
rect 16476 11027 16534 11033
rect 18138 11024 18144 11036
rect 18196 11024 18202 11076
rect 18230 11024 18236 11076
rect 18288 11064 18294 11076
rect 19720 11073 19748 11104
rect 34790 11092 34796 11104
rect 34848 11092 34854 11144
rect 19705 11067 19763 11073
rect 19705 11064 19717 11067
rect 18288 11036 19717 11064
rect 18288 11024 18294 11036
rect 19705 11033 19717 11036
rect 19751 11033 19763 11067
rect 19705 11027 19763 11033
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 37826 11064 37832 11076
rect 20220 11036 37832 11064
rect 20220 11024 20226 11036
rect 37826 11024 37832 11036
rect 37884 11024 37890 11076
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 19245 10999 19303 11005
rect 19245 10996 19257 10999
rect 18012 10968 19257 10996
rect 18012 10956 18018 10968
rect 19245 10965 19257 10968
rect 19291 10965 19303 10999
rect 19245 10959 19303 10965
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 2866 10792 2872 10804
rect 2827 10764 2872 10792
rect 2866 10752 2872 10764
rect 2924 10752 2930 10804
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 8202 10792 8208 10804
rect 3476 10764 8208 10792
rect 3476 10752 3482 10764
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 17497 10795 17555 10801
rect 8352 10764 12434 10792
rect 8352 10752 8358 10764
rect 4341 10727 4399 10733
rect 4341 10693 4353 10727
rect 4387 10724 4399 10727
rect 5258 10724 5264 10736
rect 4387 10696 5264 10724
rect 4387 10693 4399 10696
rect 4341 10687 4399 10693
rect 5258 10684 5264 10696
rect 5316 10684 5322 10736
rect 10042 10684 10048 10736
rect 10100 10724 10106 10736
rect 10100 10696 10732 10724
rect 10100 10684 10106 10696
rect 3970 10616 3976 10668
rect 4028 10656 4034 10668
rect 10134 10656 10140 10668
rect 4028 10628 10140 10656
rect 4028 10616 4034 10628
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10704 10665 10732 10696
rect 10433 10659 10491 10665
rect 10433 10625 10445 10659
rect 10479 10656 10491 10659
rect 10689 10659 10747 10665
rect 10479 10628 10640 10656
rect 10479 10625 10491 10628
rect 10433 10619 10491 10625
rect 10612 10588 10640 10628
rect 10689 10625 10701 10659
rect 10735 10656 10747 10659
rect 10962 10656 10968 10668
rect 10735 10628 10968 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 12406 10656 12434 10764
rect 17497 10761 17509 10795
rect 17543 10761 17555 10795
rect 17497 10755 17555 10761
rect 14544 10727 14602 10733
rect 14544 10693 14556 10727
rect 14590 10724 14602 10727
rect 17512 10724 17540 10755
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 18785 10795 18843 10801
rect 18785 10792 18797 10795
rect 18748 10764 18797 10792
rect 18748 10752 18754 10764
rect 18785 10761 18797 10764
rect 18831 10761 18843 10795
rect 19242 10792 19248 10804
rect 19203 10764 19248 10792
rect 18785 10755 18843 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 19978 10792 19984 10804
rect 19939 10764 19984 10792
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20162 10752 20168 10804
rect 20220 10792 20226 10804
rect 20441 10795 20499 10801
rect 20441 10792 20453 10795
rect 20220 10764 20453 10792
rect 20220 10752 20226 10764
rect 20441 10761 20453 10764
rect 20487 10761 20499 10795
rect 20441 10755 20499 10761
rect 14590 10696 17540 10724
rect 14590 10693 14602 10696
rect 14544 10687 14602 10693
rect 18046 10684 18052 10736
rect 18104 10724 18110 10736
rect 19153 10727 19211 10733
rect 19153 10724 19165 10727
rect 18104 10696 19165 10724
rect 18104 10684 18110 10696
rect 19153 10693 19165 10696
rect 19199 10693 19211 10727
rect 19260 10724 19288 10752
rect 19260 10696 22094 10724
rect 19153 10687 19211 10693
rect 17681 10659 17739 10665
rect 12406 10628 15332 10656
rect 10870 10588 10876 10600
rect 10612 10560 10876 10588
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 14274 10588 14280 10600
rect 14235 10560 14280 10588
rect 14274 10548 14280 10560
rect 14332 10548 14338 10600
rect 15304 10588 15332 10628
rect 17681 10625 17693 10659
rect 17727 10656 17739 10659
rect 17954 10656 17960 10668
rect 17727 10628 17960 10656
rect 17727 10625 17739 10628
rect 17681 10619 17739 10625
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18874 10656 18880 10668
rect 18371 10628 18880 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 20346 10656 20352 10668
rect 20307 10628 20352 10656
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 19429 10591 19487 10597
rect 15304 10560 18368 10588
rect 15657 10523 15715 10529
rect 15657 10489 15669 10523
rect 15703 10520 15715 10523
rect 18230 10520 18236 10532
rect 15703 10492 18236 10520
rect 15703 10489 15715 10492
rect 15657 10483 15715 10489
rect 18230 10480 18236 10492
rect 18288 10480 18294 10532
rect 18340 10520 18368 10560
rect 19429 10557 19441 10591
rect 19475 10588 19487 10591
rect 19978 10588 19984 10600
rect 19475 10560 19984 10588
rect 19475 10557 19487 10560
rect 19429 10551 19487 10557
rect 19978 10548 19984 10560
rect 20036 10588 20042 10600
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 20036 10560 20545 10588
rect 20036 10548 20042 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 22066 10588 22094 10696
rect 35894 10588 35900 10600
rect 22066 10560 35900 10588
rect 20533 10551 20591 10557
rect 35894 10548 35900 10560
rect 35952 10548 35958 10600
rect 20070 10520 20076 10532
rect 18340 10492 20076 10520
rect 20070 10480 20076 10492
rect 20128 10480 20134 10532
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 11054 10452 11060 10464
rect 9355 10424 11060 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 18141 10455 18199 10461
rect 18141 10452 18153 10455
rect 15804 10424 18153 10452
rect 15804 10412 15810 10424
rect 18141 10421 18153 10424
rect 18187 10421 18199 10455
rect 18141 10415 18199 10421
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 20530 10452 20536 10464
rect 19484 10424 20536 10452
rect 19484 10412 19490 10424
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11020 10220 11713 10248
rect 11020 10208 11026 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 17862 10248 17868 10260
rect 17823 10220 17868 10248
rect 11701 10211 11759 10217
rect 11716 10112 11744 10211
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 18432 10220 18521 10248
rect 18138 10140 18144 10192
rect 18196 10180 18202 10192
rect 18432 10180 18460 10220
rect 18509 10217 18521 10220
rect 18555 10217 18567 10251
rect 18509 10211 18567 10217
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 19521 10251 19579 10257
rect 19521 10248 19533 10251
rect 18932 10220 19533 10248
rect 18932 10208 18938 10220
rect 19521 10217 19533 10220
rect 19567 10217 19579 10251
rect 19521 10211 19579 10217
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20036 10220 21220 10248
rect 20036 10208 20042 10220
rect 18196 10152 18460 10180
rect 18196 10140 18202 10152
rect 18598 10140 18604 10192
rect 18656 10180 18662 10192
rect 20717 10183 20775 10189
rect 20717 10180 20729 10183
rect 18656 10152 20729 10180
rect 18656 10140 18662 10152
rect 20717 10149 20729 10152
rect 20763 10149 20775 10183
rect 20717 10143 20775 10149
rect 14274 10112 14280 10124
rect 11716 10084 14280 10112
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 20073 10115 20131 10121
rect 20073 10112 20085 10115
rect 20036 10084 20085 10112
rect 20036 10072 20042 10084
rect 20073 10081 20085 10084
rect 20119 10081 20131 10115
rect 21192 10112 21220 10220
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 21192 10084 21281 10112
rect 20073 10075 20131 10081
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 2866 10044 2872 10056
rect 1903 10016 2872 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 10410 10044 10416 10056
rect 10371 10016 10416 10044
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 14544 10047 14602 10053
rect 14544 10013 14556 10047
rect 14590 10044 14602 10047
rect 15746 10044 15752 10056
rect 14590 10016 15752 10044
rect 14590 10013 14602 10016
rect 14544 10007 14602 10013
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 17954 10044 17960 10056
rect 17696 10016 17960 10044
rect 2124 9979 2182 9985
rect 2124 9945 2136 9979
rect 2170 9976 2182 9979
rect 3786 9976 3792 9988
rect 2170 9948 3792 9976
rect 2170 9945 2182 9948
rect 2124 9939 2182 9945
rect 3786 9936 3792 9948
rect 3844 9936 3850 9988
rect 17696 9976 17724 10016
rect 17954 10004 17960 10016
rect 18012 10004 18018 10056
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10044 18107 10047
rect 18414 10044 18420 10056
rect 18095 10016 18420 10044
rect 18095 10013 18107 10016
rect 18049 10007 18107 10013
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 18690 10044 18696 10056
rect 18651 10016 18696 10044
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 18874 10004 18880 10056
rect 18932 10044 18938 10056
rect 21085 10047 21143 10053
rect 21085 10044 21097 10047
rect 18932 10016 21097 10044
rect 18932 10004 18938 10016
rect 21085 10013 21097 10016
rect 21131 10013 21143 10047
rect 32858 10044 32864 10056
rect 21085 10007 21143 10013
rect 22066 10016 32864 10044
rect 12406 9948 17724 9976
rect 19889 9979 19947 9985
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 4614 9908 4620 9920
rect 3283 9880 4620 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 12406 9908 12434 9948
rect 19889 9945 19901 9979
rect 19935 9976 19947 9979
rect 20162 9976 20168 9988
rect 19935 9948 20168 9976
rect 19935 9945 19947 9948
rect 19889 9939 19947 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 22066 9976 22094 10016
rect 32858 10004 32864 10016
rect 32916 10004 32922 10056
rect 20640 9948 22094 9976
rect 10192 9880 12434 9908
rect 15657 9911 15715 9917
rect 10192 9868 10198 9880
rect 15657 9877 15669 9911
rect 15703 9908 15715 9911
rect 18414 9908 18420 9920
rect 15703 9880 18420 9908
rect 15703 9877 15715 9880
rect 15657 9871 15715 9877
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 18506 9868 18512 9920
rect 18564 9908 18570 9920
rect 19426 9908 19432 9920
rect 18564 9880 19432 9908
rect 18564 9868 18570 9880
rect 19426 9868 19432 9880
rect 19484 9908 19490 9920
rect 19981 9911 20039 9917
rect 19981 9908 19993 9911
rect 19484 9880 19993 9908
rect 19484 9868 19490 9880
rect 19981 9877 19993 9880
rect 20027 9908 20039 9911
rect 20640 9908 20668 9948
rect 20027 9880 20668 9908
rect 20027 9877 20039 9880
rect 19981 9871 20039 9877
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 21177 9911 21235 9917
rect 21177 9908 21189 9911
rect 20772 9880 21189 9908
rect 20772 9868 20778 9880
rect 21177 9877 21189 9880
rect 21223 9908 21235 9911
rect 33870 9908 33876 9920
rect 21223 9880 33876 9908
rect 21223 9877 21235 9880
rect 21177 9871 21235 9877
rect 33870 9868 33876 9880
rect 33928 9868 33934 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18230 9704 18236 9716
rect 18012 9676 18236 9704
rect 18012 9664 18018 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 18690 9664 18696 9716
rect 18748 9704 18754 9716
rect 19153 9707 19211 9713
rect 19153 9704 19165 9707
rect 18748 9676 19165 9704
rect 18748 9664 18754 9676
rect 19153 9673 19165 9676
rect 19199 9673 19211 9707
rect 19153 9667 19211 9673
rect 20625 9639 20683 9645
rect 20625 9605 20637 9639
rect 20671 9636 20683 9639
rect 20714 9636 20720 9648
rect 20671 9608 20720 9636
rect 20671 9605 20683 9608
rect 20625 9599 20683 9605
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3050 9568 3056 9580
rect 3007 9540 3056 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 8938 9568 8944 9580
rect 8899 9540 8944 9568
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 10962 9568 10968 9580
rect 10923 9540 10968 9568
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 14274 9568 14280 9580
rect 14235 9540 14280 9568
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 14544 9571 14602 9577
rect 14544 9537 14556 9571
rect 14590 9568 14602 9571
rect 15562 9568 15568 9580
rect 14590 9540 15568 9568
rect 14590 9537 14602 9540
rect 14544 9531 14602 9537
rect 15562 9528 15568 9540
rect 15620 9528 15626 9580
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 19242 9568 19248 9580
rect 18739 9540 19248 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19521 9571 19579 9577
rect 19521 9568 19533 9571
rect 19392 9540 19533 9568
rect 19392 9528 19398 9540
rect 19521 9537 19533 9540
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 18141 9503 18199 9509
rect 18141 9469 18153 9503
rect 18187 9500 18199 9503
rect 19150 9500 19156 9512
rect 18187 9472 19156 9500
rect 18187 9469 18199 9472
rect 18141 9463 18199 9469
rect 19150 9460 19156 9472
rect 19208 9500 19214 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19208 9472 19625 9500
rect 19208 9460 19214 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9500 19855 9503
rect 19978 9500 19984 9512
rect 19843 9472 19984 9500
rect 19843 9469 19855 9472
rect 19797 9463 19855 9469
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 2777 9435 2835 9441
rect 2777 9401 2789 9435
rect 2823 9432 2835 9435
rect 2958 9432 2964 9444
rect 2823 9404 2964 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 2958 9392 2964 9404
rect 3016 9392 3022 9444
rect 8754 9432 8760 9444
rect 8715 9404 8760 9432
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 10778 9432 10784 9444
rect 10739 9404 10784 9432
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9432 15715 9435
rect 17310 9432 17316 9444
rect 15703 9404 17316 9432
rect 15703 9401 15715 9404
rect 15657 9395 15715 9401
rect 17310 9392 17316 9404
rect 17368 9432 17374 9444
rect 37274 9432 37280 9444
rect 17368 9404 37280 9432
rect 17368 9392 17374 9404
rect 37274 9392 37280 9404
rect 37332 9392 37338 9444
rect 11974 9324 11980 9376
rect 12032 9364 12038 9376
rect 15470 9364 15476 9376
rect 12032 9336 15476 9364
rect 12032 9324 12038 9336
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 3786 9160 3792 9172
rect 3747 9132 3792 9160
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 5629 9163 5687 9169
rect 5629 9160 5641 9163
rect 5592 9132 5641 9160
rect 5592 9120 5598 9132
rect 5629 9129 5641 9132
rect 5675 9129 5687 9163
rect 5629 9123 5687 9129
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 8904 9132 9873 9160
rect 8904 9120 8910 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 9861 9123 9919 9129
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 11425 9163 11483 9169
rect 11425 9160 11437 9163
rect 11388 9132 11437 9160
rect 11388 9120 11394 9132
rect 11425 9129 11437 9132
rect 11471 9129 11483 9163
rect 11425 9123 11483 9129
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 26510 9160 26516 9172
rect 15528 9132 26516 9160
rect 15528 9120 15534 9132
rect 26510 9120 26516 9132
rect 26568 9120 26574 9172
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 5077 9095 5135 9101
rect 5077 9092 5089 9095
rect 2556 9064 5089 9092
rect 2556 9052 2562 9064
rect 5077 9061 5089 9064
rect 5123 9061 5135 9095
rect 14090 9092 14096 9104
rect 5077 9055 5135 9061
rect 6886 9064 14096 9092
rect 3142 9024 3148 9036
rect 3068 8996 3148 9024
rect 2590 8956 2596 8968
rect 2551 8928 2596 8956
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 3068 8965 3096 8996
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4614 9024 4620 9036
rect 4295 8996 4620 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 5092 9024 5120 9055
rect 6089 9027 6147 9033
rect 6089 9024 6101 9027
rect 5092 8996 6101 9024
rect 6089 8993 6101 8996
rect 6135 8993 6147 9027
rect 6089 8987 6147 8993
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 9024 6331 9027
rect 6886 9024 6914 9064
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 19426 9092 19432 9104
rect 19387 9064 19432 9092
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 6319 8996 6914 9024
rect 6319 8993 6331 8996
rect 6273 8987 6331 8993
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 2832 8928 3065 8956
rect 2832 8916 2838 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3053 8919 3111 8925
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 4154 8956 4160 8968
rect 4115 8928 4160 8956
rect 3973 8919 4031 8925
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 3988 8888 4016 8919
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 6104 8956 6132 8987
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10008 8996 10180 9024
rect 10008 8984 10014 8996
rect 6638 8956 6644 8968
rect 6104 8928 6644 8956
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 10152 8965 10180 8996
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 26234 9024 26240 9036
rect 13412 8996 26240 9024
rect 13412 8984 13418 8996
rect 26234 8984 26240 8996
rect 26292 8984 26298 9036
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 10137 8919 10195 8925
rect 5166 8888 5172 8900
rect 2924 8860 5172 8888
rect 2924 8848 2930 8860
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 10060 8888 10088 8919
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 10502 8956 10508 8968
rect 10459 8928 10508 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 12342 8956 12348 8968
rect 11655 8928 12348 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 27062 8956 27068 8968
rect 16540 8928 27068 8956
rect 16540 8916 16546 8928
rect 27062 8916 27068 8928
rect 27120 8916 27126 8968
rect 11790 8888 11796 8900
rect 10060 8860 11796 8888
rect 11790 8848 11796 8860
rect 11848 8848 11854 8900
rect 3234 8820 3240 8832
rect 3195 8792 3240 8820
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 5994 8820 6000 8832
rect 5955 8792 6000 8820
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 2593 8619 2651 8625
rect 2593 8585 2605 8619
rect 2639 8616 2651 8619
rect 2866 8616 2872 8628
rect 2639 8588 2872 8616
rect 2639 8585 2651 8588
rect 2593 8579 2651 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3050 8616 3056 8628
rect 3011 8588 3056 8616
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8585 4215 8619
rect 4706 8616 4712 8628
rect 4667 8588 4712 8616
rect 4157 8579 4215 8585
rect 2774 8548 2780 8560
rect 2516 8520 2780 8548
rect 2516 8421 2544 8520
rect 2774 8508 2780 8520
rect 2832 8508 2838 8560
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 4172 8548 4200 8579
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 5626 8616 5632 8628
rect 4816 8588 5632 8616
rect 4816 8548 4844 8588
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6052 8588 6561 8616
rect 6052 8576 6058 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 7834 8616 7840 8628
rect 7795 8588 7840 8616
rect 6549 8579 6607 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8938 8616 8944 8628
rect 8899 8588 8944 8616
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 10962 8616 10968 8628
rect 10923 8588 10968 8616
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8585 11575 8619
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 11517 8579 11575 8585
rect 3292 8520 4108 8548
rect 4172 8520 4844 8548
rect 3292 8508 3298 8520
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 2685 8443 2743 8449
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2700 8344 2728 8443
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 3786 8480 3792 8492
rect 3660 8452 3705 8480
rect 3747 8452 3792 8480
rect 3660 8440 3666 8452
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 3978 8483 4036 8489
rect 3978 8449 3990 8483
rect 4024 8480 4036 8483
rect 4080 8480 4108 8520
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 9122 8548 9128 8560
rect 5040 8520 5396 8548
rect 5040 8508 5046 8520
rect 4024 8452 4108 8480
rect 4024 8449 4036 8452
rect 3978 8443 4036 8449
rect 3234 8372 3240 8424
rect 3292 8412 3298 8424
rect 3896 8412 3924 8443
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4212 8452 4905 8480
rect 4212 8440 4218 8452
rect 4893 8449 4905 8452
rect 4939 8480 4951 8483
rect 5074 8480 5080 8492
rect 4939 8452 5080 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5368 8489 5396 8520
rect 8036 8520 9128 8548
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7466 8480 7472 8492
rect 6871 8452 7472 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 3292 8384 3924 8412
rect 5184 8412 5212 8443
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8036 8489 8064 8520
rect 9122 8508 9128 8520
rect 9180 8548 9186 8560
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 9180 8520 9413 8548
rect 9180 8508 9186 8520
rect 9401 8517 9413 8520
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 10781 8551 10839 8557
rect 10781 8517 10793 8551
rect 10827 8548 10839 8551
rect 11422 8548 11428 8560
rect 10827 8520 11428 8548
rect 10827 8517 10839 8520
rect 10781 8511 10839 8517
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 11532 8480 11560 8579
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 15562 8616 15568 8628
rect 15523 8588 15568 8616
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 12066 8480 12072 8492
rect 8527 8452 11560 8480
rect 12027 8452 12072 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 6086 8412 6092 8424
rect 5184 8384 6092 8412
rect 3292 8372 3298 8384
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 6730 8412 6736 8424
rect 6691 8384 6736 8412
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7834 8412 7840 8424
rect 7055 8384 7840 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 5902 8344 5908 8356
rect 2700 8316 5908 8344
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 6932 8288 6960 8375
rect 7834 8372 7840 8384
rect 7892 8412 7898 8424
rect 8312 8412 8340 8443
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 15746 8480 15752 8492
rect 15707 8452 15752 8480
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8449 17463 8483
rect 18046 8480 18052 8492
rect 18007 8452 18052 8480
rect 17405 8443 17463 8449
rect 7892 8384 8340 8412
rect 7892 8372 7898 8384
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 17420 8412 17448 8443
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 14976 8384 17448 8412
rect 18141 8415 18199 8421
rect 14976 8372 14982 8384
rect 18141 8381 18153 8415
rect 18187 8412 18199 8415
rect 19978 8412 19984 8424
rect 18187 8384 19984 8412
rect 18187 8381 18199 8384
rect 18141 8375 18199 8381
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 9033 8347 9091 8353
rect 9033 8344 9045 8347
rect 8996 8316 9045 8344
rect 8996 8304 9002 8316
rect 9033 8313 9045 8316
rect 9079 8313 9091 8347
rect 9033 8307 9091 8313
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 10318 8344 10324 8356
rect 9180 8316 10324 8344
rect 9180 8304 9186 8316
rect 10318 8304 10324 8316
rect 10376 8344 10382 8356
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 10376 8316 10425 8344
rect 10376 8304 10382 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 10413 8307 10471 8313
rect 6914 8236 6920 8288
rect 6972 8236 6978 8288
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10781 8279 10839 8285
rect 10781 8276 10793 8279
rect 10008 8248 10793 8276
rect 10008 8236 10014 8248
rect 10781 8245 10793 8248
rect 10827 8245 10839 8279
rect 10781 8239 10839 8245
rect 11701 8279 11759 8285
rect 11701 8245 11713 8279
rect 11747 8276 11759 8279
rect 11974 8276 11980 8288
rect 11747 8248 11980 8276
rect 11747 8245 11759 8248
rect 11701 8239 11759 8245
rect 11974 8236 11980 8248
rect 12032 8276 12038 8288
rect 12529 8279 12587 8285
rect 12529 8276 12541 8279
rect 12032 8248 12541 8276
rect 12032 8236 12038 8248
rect 12529 8245 12541 8248
rect 12575 8245 12587 8279
rect 12529 8239 12587 8245
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 18693 8279 18751 8285
rect 18693 8276 18705 8279
rect 18196 8248 18705 8276
rect 18196 8236 18202 8248
rect 18693 8245 18705 8248
rect 18739 8245 18751 8279
rect 18693 8239 18751 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3568 8044 3801 8072
rect 3568 8032 3574 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 5074 8072 5080 8084
rect 5035 8044 5080 8072
rect 3789 8035 3847 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5902 8072 5908 8084
rect 5863 8044 5908 8072
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 6825 8075 6883 8081
rect 6825 8041 6837 8075
rect 6871 8072 6883 8075
rect 6914 8072 6920 8084
rect 6871 8044 6920 8072
rect 6871 8041 6883 8044
rect 6825 8035 6883 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 9950 8072 9956 8084
rect 9911 8044 9956 8072
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10502 8072 10508 8084
rect 10152 8044 10508 8072
rect 3234 8004 3240 8016
rect 3195 7976 3240 8004
rect 3234 7964 3240 7976
rect 3292 7964 3298 8016
rect 8202 8004 8208 8016
rect 3988 7976 8208 8004
rect 2038 7896 2044 7948
rect 2096 7936 2102 7948
rect 3988 7936 4016 7976
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 4614 7936 4620 7948
rect 2096 7908 4016 7936
rect 4264 7908 4620 7936
rect 2096 7896 2102 7908
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 2869 7871 2927 7877
rect 2869 7868 2881 7871
rect 2832 7840 2881 7868
rect 2832 7828 2838 7840
rect 2869 7837 2881 7840
rect 2915 7837 2927 7871
rect 2869 7831 2927 7837
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3142 7868 3148 7880
rect 3099 7840 3148 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 4264 7877 4292 7908
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 10152 7945 10180 8044
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 11790 8072 11796 8084
rect 11751 8044 11796 8072
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 14090 8072 14096 8084
rect 14051 8044 14096 8072
rect 14090 8032 14096 8044
rect 14148 8032 14154 8084
rect 14645 8075 14703 8081
rect 14645 8041 14657 8075
rect 14691 8072 14703 8075
rect 16114 8072 16120 8084
rect 14691 8044 16120 8072
rect 14691 8041 14703 8044
rect 14645 8035 14703 8041
rect 10413 8007 10471 8013
rect 10413 7973 10425 8007
rect 10459 8004 10471 8007
rect 14918 8004 14924 8016
rect 10459 7976 14924 8004
rect 10459 7973 10471 7976
rect 10413 7967 10471 7973
rect 14918 7964 14924 7976
rect 14976 7964 14982 8016
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7905 10195 7939
rect 11054 7936 11060 7948
rect 10137 7899 10195 7905
rect 10244 7908 11060 7936
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3660 7840 3985 7868
rect 3660 7828 3666 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 4798 7868 4804 7880
rect 4488 7840 4804 7868
rect 4488 7828 4494 7840
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6236 7840 6281 7868
rect 6236 7828 6242 7840
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6696 7840 6745 7868
rect 6696 7828 6702 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 10244 7877 10272 7908
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 11164 7908 13768 7936
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 6880 7840 7573 7868
rect 6880 7828 6886 7840
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10502 7828 10508 7880
rect 10560 7868 10566 7880
rect 10560 7840 11100 7868
rect 10560 7828 10566 7840
rect 4816 7800 4844 7828
rect 5445 7803 5503 7809
rect 5445 7800 5457 7803
rect 4816 7772 5457 7800
rect 5445 7769 5457 7772
rect 5491 7769 5503 7803
rect 5445 7763 5503 7769
rect 9953 7803 10011 7809
rect 9953 7769 9965 7803
rect 9999 7800 10011 7803
rect 10134 7800 10140 7812
rect 9999 7772 10140 7800
rect 9999 7769 10011 7772
rect 9953 7763 10011 7769
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 10410 7760 10416 7812
rect 10468 7800 10474 7812
rect 10686 7800 10692 7812
rect 10468 7772 10692 7800
rect 10468 7760 10474 7772
rect 10686 7760 10692 7772
rect 10744 7800 10750 7812
rect 11072 7809 11100 7840
rect 10873 7803 10931 7809
rect 10873 7800 10885 7803
rect 10744 7772 10885 7800
rect 10744 7760 10750 7772
rect 10873 7769 10885 7772
rect 10919 7769 10931 7803
rect 10873 7763 10931 7769
rect 11057 7803 11115 7809
rect 11057 7769 11069 7803
rect 11103 7769 11115 7803
rect 11057 7763 11115 7769
rect 5245 7735 5303 7741
rect 5245 7701 5257 7735
rect 5291 7732 5303 7735
rect 5718 7732 5724 7744
rect 5291 7704 5724 7732
rect 5291 7701 5303 7704
rect 5245 7695 5303 7701
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9674 7732 9680 7744
rect 9539 7704 9680 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10888 7732 10916 7763
rect 11164 7732 11192 7908
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11480 7840 11897 7868
rect 11480 7828 11486 7840
rect 11885 7837 11897 7840
rect 11931 7868 11943 7871
rect 13170 7868 13176 7880
rect 11931 7840 13176 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 13740 7800 13768 7908
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 14369 7939 14427 7945
rect 14369 7936 14381 7939
rect 13872 7908 14381 7936
rect 13872 7896 13878 7908
rect 14369 7905 14381 7908
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 13964 7840 14289 7868
rect 13964 7828 13970 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 15028 7868 15056 8044
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 18046 8004 18052 8016
rect 17052 7976 18052 8004
rect 17052 7945 17080 7976
rect 18046 7964 18052 7976
rect 18104 7964 18110 8016
rect 17037 7939 17095 7945
rect 17037 7905 17049 7939
rect 17083 7905 17095 7939
rect 17037 7899 17095 7905
rect 17129 7939 17187 7945
rect 17129 7905 17141 7939
rect 17175 7936 17187 7939
rect 17957 7939 18015 7945
rect 17957 7936 17969 7939
rect 17175 7908 17969 7936
rect 17175 7905 17187 7908
rect 17129 7899 17187 7905
rect 17957 7905 17969 7908
rect 18003 7905 18015 7939
rect 17957 7899 18015 7905
rect 17052 7868 17080 7899
rect 17218 7868 17224 7880
rect 14277 7831 14335 7837
rect 14384 7840 15056 7868
rect 15396 7840 17080 7868
rect 17179 7840 17224 7868
rect 14384 7800 14412 7840
rect 13740 7772 14412 7800
rect 14737 7803 14795 7809
rect 14737 7769 14749 7803
rect 14783 7800 14795 7803
rect 14918 7800 14924 7812
rect 14783 7772 14924 7800
rect 14783 7769 14795 7772
rect 14737 7763 14795 7769
rect 14918 7760 14924 7772
rect 14976 7800 14982 7812
rect 15396 7800 15424 7840
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 18046 7868 18052 7880
rect 17368 7840 17413 7868
rect 18007 7840 18052 7868
rect 17368 7828 17374 7840
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 14976 7772 15424 7800
rect 16393 7803 16451 7809
rect 14976 7760 14982 7772
rect 16393 7769 16405 7803
rect 16439 7800 16451 7803
rect 17328 7800 17356 7828
rect 16439 7772 17356 7800
rect 16439 7769 16451 7772
rect 16393 7763 16451 7769
rect 10888 7704 11192 7732
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 16850 7732 16856 7744
rect 11296 7704 11341 7732
rect 16811 7704 16856 7732
rect 11296 7692 11302 7704
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2590 7528 2596 7540
rect 2455 7500 2596 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 3786 7528 3792 7540
rect 3747 7500 3792 7528
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7834 7528 7840 7540
rect 7795 7500 7840 7528
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 9122 7528 9128 7540
rect 9083 7500 9128 7528
rect 9122 7488 9128 7500
rect 9180 7528 9186 7540
rect 9398 7528 9404 7540
rect 9180 7500 9404 7528
rect 9180 7488 9186 7500
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 11514 7528 11520 7540
rect 10735 7500 11520 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 14918 7528 14924 7540
rect 14879 7500 14924 7528
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15804 7500 16037 7528
rect 15804 7488 15810 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16025 7491 16083 7497
rect 16945 7531 17003 7537
rect 16945 7497 16957 7531
rect 16991 7528 17003 7531
rect 17218 7528 17224 7540
rect 16991 7500 17224 7528
rect 16991 7497 17003 7500
rect 16945 7491 17003 7497
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 20254 7528 20260 7540
rect 20215 7500 20260 7528
rect 20254 7488 20260 7500
rect 20312 7488 20318 7540
rect 2777 7463 2835 7469
rect 2777 7429 2789 7463
rect 2823 7460 2835 7463
rect 2866 7460 2872 7472
rect 2823 7432 2872 7460
rect 2823 7429 2835 7432
rect 2777 7423 2835 7429
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 3712 7432 4568 7460
rect 3142 7392 3148 7404
rect 2884 7364 3148 7392
rect 2884 7333 2912 7364
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3712 7401 3740 7432
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 4430 7392 4436 7404
rect 3927 7364 4436 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4540 7401 4568 7432
rect 6886 7432 8156 7460
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7392 4583 7395
rect 4614 7392 4620 7404
rect 4571 7364 4620 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7392 4767 7395
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 4755 7364 5641 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 5629 7361 5641 7364
rect 5675 7392 5687 7395
rect 6178 7392 6184 7404
rect 5675 7364 6184 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 6886 7392 6914 7432
rect 6288 7364 6914 7392
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7293 2927 7327
rect 3050 7324 3056 7336
rect 3011 7296 3056 7324
rect 2869 7287 2927 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 5258 7324 5264 7336
rect 5171 7296 5264 7324
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7324 5411 7327
rect 5718 7324 5724 7336
rect 5399 7296 5724 7324
rect 5399 7293 5411 7296
rect 5353 7287 5411 7293
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 5276 7256 5304 7284
rect 6288 7256 6316 7364
rect 7742 7352 7748 7404
rect 7800 7392 7806 7404
rect 8018 7392 8024 7404
rect 7800 7364 8024 7392
rect 7800 7352 7806 7364
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8128 7392 8156 7432
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 9033 7463 9091 7469
rect 9033 7460 9045 7463
rect 8260 7432 9045 7460
rect 8260 7420 8266 7432
rect 9033 7429 9045 7432
rect 9079 7460 9091 7463
rect 9674 7460 9680 7472
rect 9079 7432 9680 7460
rect 9079 7429 9091 7432
rect 9033 7423 9091 7429
rect 9674 7420 9680 7432
rect 9732 7460 9738 7472
rect 9950 7460 9956 7472
rect 9732 7432 9956 7460
rect 9732 7420 9738 7432
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 14936 7460 14964 7488
rect 15838 7460 15844 7472
rect 10336 7432 14964 7460
rect 15799 7432 15844 7460
rect 10336 7392 10364 7432
rect 15838 7420 15844 7432
rect 15896 7420 15902 7472
rect 19518 7420 19524 7472
rect 19576 7460 19582 7472
rect 20073 7463 20131 7469
rect 20073 7460 20085 7463
rect 19576 7432 20085 7460
rect 19576 7420 19582 7432
rect 20073 7429 20085 7432
rect 20119 7460 20131 7463
rect 20119 7432 20760 7460
rect 20119 7429 20131 7432
rect 20073 7423 20131 7429
rect 10502 7392 10508 7404
rect 8128 7364 10364 7392
rect 10463 7364 10508 7392
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 13722 7392 13728 7404
rect 13683 7364 13728 7392
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13832 7364 13921 7392
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 6880 7296 8217 7324
rect 6880 7284 6886 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7324 8355 7327
rect 9490 7324 9496 7336
rect 8343 7296 9496 7324
rect 8343 7293 8355 7296
rect 8297 7287 8355 7293
rect 9490 7284 9496 7296
rect 9548 7284 9554 7336
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 13832 7324 13860 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 14550 7392 14556 7404
rect 14511 7364 14556 7392
rect 13909 7355 13967 7361
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 15194 7392 15200 7404
rect 14783 7364 15200 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 15194 7352 15200 7364
rect 15252 7392 15258 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 15252 7364 16865 7392
rect 15252 7352 15258 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7392 19947 7395
rect 19978 7392 19984 7404
rect 19935 7364 19984 7392
rect 19935 7361 19947 7364
rect 19889 7355 19947 7361
rect 19978 7352 19984 7364
rect 20036 7352 20042 7404
rect 20732 7401 20760 7432
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 11940 7296 13860 7324
rect 11940 7284 11946 7296
rect 5276 7228 6316 7256
rect 13832 7256 13860 7296
rect 14090 7284 14096 7336
rect 14148 7324 14154 7336
rect 19337 7327 19395 7333
rect 19337 7324 19349 7327
rect 14148 7296 19349 7324
rect 14148 7284 14154 7296
rect 19337 7293 19349 7296
rect 19383 7324 19395 7327
rect 19794 7324 19800 7336
rect 19383 7296 19800 7324
rect 19383 7293 19395 7296
rect 19337 7287 19395 7293
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 15010 7256 15016 7268
rect 13832 7228 15016 7256
rect 15010 7216 15016 7228
rect 15068 7216 15074 7268
rect 15473 7259 15531 7265
rect 15473 7225 15485 7259
rect 15519 7225 15531 7259
rect 15473 7219 15531 7225
rect 5534 7188 5540 7200
rect 5495 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 13262 7188 13268 7200
rect 13223 7160 13268 7188
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14093 7191 14151 7197
rect 14093 7188 14105 7191
rect 13872 7160 14105 7188
rect 13872 7148 13878 7160
rect 14093 7157 14105 7160
rect 14139 7157 14151 7191
rect 14093 7151 14151 7157
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 14553 7191 14611 7197
rect 14553 7188 14565 7191
rect 14240 7160 14565 7188
rect 14240 7148 14246 7160
rect 14553 7157 14565 7160
rect 14599 7157 14611 7191
rect 14553 7151 14611 7157
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 15488 7188 15516 7219
rect 14700 7160 15516 7188
rect 15841 7191 15899 7197
rect 14700 7148 14706 7160
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 16850 7188 16856 7200
rect 15887 7160 16856 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 20901 7191 20959 7197
rect 20901 7157 20913 7191
rect 20947 7188 20959 7191
rect 21450 7188 21456 7200
rect 20947 7160 21456 7188
rect 20947 7157 20959 7160
rect 20901 7151 20959 7157
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 3053 6987 3111 6993
rect 3053 6953 3065 6987
rect 3099 6984 3111 6987
rect 3602 6984 3608 6996
rect 3099 6956 3608 6984
rect 3099 6953 3111 6956
rect 3053 6947 3111 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5997 6987 6055 6993
rect 5997 6984 6009 6987
rect 5592 6956 6009 6984
rect 5592 6944 5598 6956
rect 5997 6953 6009 6956
rect 6043 6953 6055 6987
rect 11790 6984 11796 6996
rect 5997 6947 6055 6953
rect 6104 6956 11796 6984
rect 4338 6876 4344 6928
rect 4396 6916 4402 6928
rect 6104 6916 6132 6956
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12216 6956 13124 6984
rect 12216 6944 12222 6956
rect 4396 6888 6132 6916
rect 4396 6876 4402 6888
rect 6178 6876 6184 6928
rect 6236 6916 6242 6928
rect 6549 6919 6607 6925
rect 6549 6916 6561 6919
rect 6236 6888 6561 6916
rect 6236 6876 6242 6888
rect 6549 6885 6561 6888
rect 6595 6885 6607 6919
rect 6549 6879 6607 6885
rect 12802 6876 12808 6928
rect 12860 6916 12866 6928
rect 12860 6888 13032 6916
rect 12860 6876 12866 6888
rect 6822 6848 6828 6860
rect 5920 6820 6828 6848
rect 2774 6780 2780 6792
rect 2735 6752 2780 6780
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 3050 6780 3056 6792
rect 2832 6752 3056 6780
rect 2832 6740 2838 6752
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 5920 6789 5948 6820
rect 6822 6808 6828 6820
rect 6880 6848 6886 6860
rect 8938 6848 8944 6860
rect 6880 6820 8064 6848
rect 8899 6820 8944 6848
rect 6880 6808 6886 6820
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5684 6752 5917 6780
rect 5684 6740 5690 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6780 6791 6783
rect 7834 6780 7840 6792
rect 6779 6752 7840 6780
rect 6779 6749 6791 6752
rect 6733 6743 6791 6749
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 2924 6684 3832 6712
rect 2924 6672 2930 6684
rect 3804 6656 3832 6684
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3237 6647 3295 6653
rect 3237 6644 3249 6647
rect 3200 6616 3249 6644
rect 3200 6604 3206 6616
rect 3237 6613 3249 6616
rect 3283 6613 3295 6647
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3237 6607 3295 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 6104 6644 6132 6743
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8036 6780 8064 6820
rect 8938 6808 8944 6820
rect 8996 6808 9002 6860
rect 9306 6848 9312 6860
rect 9267 6820 9312 6848
rect 9306 6808 9312 6820
rect 9364 6848 9370 6860
rect 11054 6848 11060 6860
rect 9364 6820 11060 6848
rect 9364 6808 9370 6820
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 11974 6848 11980 6860
rect 11848 6820 11980 6848
rect 11848 6808 11854 6820
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 13004 6857 13032 6888
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 13096 6848 13124 6956
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13780 6956 14105 6984
rect 13780 6944 13786 6956
rect 14093 6953 14105 6956
rect 14139 6984 14151 6987
rect 14274 6984 14280 6996
rect 14139 6956 14280 6984
rect 14139 6953 14151 6956
rect 14093 6947 14151 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 14461 6987 14519 6993
rect 14461 6953 14473 6987
rect 14507 6984 14519 6987
rect 14550 6984 14556 6996
rect 14507 6956 14556 6984
rect 14507 6953 14519 6956
rect 14461 6947 14519 6953
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 15010 6984 15016 6996
rect 14971 6956 15016 6984
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 15565 6987 15623 6993
rect 15565 6953 15577 6987
rect 15611 6984 15623 6987
rect 15838 6984 15844 6996
rect 15611 6956 15844 6984
rect 15611 6953 15623 6956
rect 15565 6947 15623 6953
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 16117 6987 16175 6993
rect 16117 6953 16129 6987
rect 16163 6953 16175 6987
rect 19794 6984 19800 6996
rect 19755 6956 19800 6984
rect 16117 6947 16175 6953
rect 15028 6916 15056 6944
rect 16132 6916 16160 6947
rect 19794 6944 19800 6956
rect 19852 6944 19858 6996
rect 18046 6916 18052 6928
rect 13740 6888 14320 6916
rect 15028 6888 18052 6916
rect 13740 6848 13768 6888
rect 13096 6820 13768 6848
rect 12989 6811 13047 6817
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8036 6752 9137 6780
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9401 6783 9459 6789
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 10134 6780 10140 6792
rect 9447 6752 10140 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 7101 6715 7159 6721
rect 6972 6684 7017 6712
rect 6972 6672 6978 6684
rect 7101 6681 7113 6715
rect 7147 6712 7159 6715
rect 8018 6712 8024 6724
rect 7147 6684 8024 6712
rect 7147 6681 7159 6684
rect 7101 6675 7159 6681
rect 8018 6672 8024 6684
rect 8076 6672 8082 6724
rect 9232 6712 9260 6743
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 14090 6780 14096 6792
rect 14051 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 14292 6789 14320 6888
rect 14366 6808 14372 6860
rect 14424 6848 14430 6860
rect 15197 6851 15255 6857
rect 15197 6848 15209 6851
rect 14424 6820 15209 6848
rect 14424 6808 14430 6820
rect 15197 6817 15209 6820
rect 15243 6817 15255 6851
rect 16209 6851 16267 6857
rect 16209 6848 16221 6851
rect 15197 6811 15255 6817
rect 15396 6820 16221 6848
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14550 6740 14556 6792
rect 14608 6780 14614 6792
rect 14921 6783 14979 6789
rect 14921 6780 14933 6783
rect 14608 6752 14933 6780
rect 14608 6740 14614 6752
rect 14921 6749 14933 6752
rect 14967 6749 14979 6783
rect 14921 6743 14979 6749
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 15396 6789 15424 6820
rect 16209 6817 16221 6820
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15344 6752 15393 6780
rect 15344 6740 15350 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 16114 6780 16120 6792
rect 16075 6752 16120 6780
rect 15381 6743 15439 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 16224 6752 16957 6780
rect 9582 6712 9588 6724
rect 9232 6684 9588 6712
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 11698 6672 11704 6724
rect 11756 6712 11762 6724
rect 12066 6712 12072 6724
rect 11756 6684 12072 6712
rect 11756 6672 11762 6684
rect 12066 6672 12072 6684
rect 12124 6712 12130 6724
rect 12805 6715 12863 6721
rect 12805 6712 12817 6715
rect 12124 6684 12817 6712
rect 12124 6672 12130 6684
rect 12805 6681 12817 6684
rect 12851 6681 12863 6715
rect 12805 6675 12863 6681
rect 6730 6644 6736 6656
rect 6104 6616 6736 6644
rect 6730 6604 6736 6616
rect 6788 6644 6794 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6788 6616 6837 6644
rect 6788 6604 6794 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 8036 6644 8064 6672
rect 11974 6644 11980 6656
rect 8036 6616 11980 6644
rect 6825 6607 6883 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12342 6644 12348 6656
rect 12303 6616 12348 6644
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12710 6644 12716 6656
rect 12671 6616 12716 6644
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 13262 6604 13268 6656
rect 13320 6644 13326 6656
rect 14182 6644 14188 6656
rect 13320 6616 14188 6644
rect 13320 6604 13326 6616
rect 14182 6604 14188 6616
rect 14240 6604 14246 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 16224 6644 16252 6752
rect 16945 6749 16957 6752
rect 16991 6749 17003 6783
rect 17678 6780 17684 6792
rect 16945 6743 17003 6749
rect 17144 6752 17684 6780
rect 16482 6644 16488 6656
rect 14332 6616 16252 6644
rect 16443 6616 16488 6644
rect 14332 6604 14338 6616
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 17144 6653 17172 6752
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 17880 6789 17908 6888
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6848 19487 6851
rect 20441 6851 20499 6857
rect 20441 6848 20453 6851
rect 19475 6820 20453 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 20441 6817 20453 6820
rect 20487 6817 20499 6851
rect 20990 6848 20996 6860
rect 20951 6820 20996 6848
rect 20441 6811 20499 6817
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 17218 6672 17224 6724
rect 17276 6712 17282 6724
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 17276 6684 17785 6712
rect 17276 6672 17282 6684
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17773 6675 17831 6681
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 18601 6647 18659 6653
rect 18601 6644 18613 6647
rect 17644 6616 18613 6644
rect 17644 6604 17650 6616
rect 18601 6613 18613 6616
rect 18647 6644 18659 6647
rect 19444 6644 19472 6811
rect 20456 6780 20484 6811
rect 20990 6808 20996 6820
rect 21048 6808 21054 6860
rect 21100 6820 21404 6848
rect 21100 6780 21128 6820
rect 21376 6789 21404 6820
rect 20456 6752 21128 6780
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 19518 6672 19524 6724
rect 19576 6712 19582 6724
rect 19797 6715 19855 6721
rect 19797 6712 19809 6715
rect 19576 6684 19809 6712
rect 19576 6672 19582 6684
rect 19797 6681 19809 6684
rect 19843 6681 19855 6715
rect 21082 6712 21088 6724
rect 19797 6675 19855 6681
rect 19996 6684 21088 6712
rect 19996 6653 20024 6684
rect 21082 6672 21088 6684
rect 21140 6672 21146 6724
rect 21192 6712 21220 6743
rect 21450 6740 21456 6792
rect 21508 6780 21514 6792
rect 22002 6780 22008 6792
rect 21508 6752 22008 6780
rect 21508 6740 21514 6752
rect 22002 6740 22008 6752
rect 22060 6740 22066 6792
rect 21726 6712 21732 6724
rect 21192 6684 21732 6712
rect 21726 6672 21732 6684
rect 21784 6672 21790 6724
rect 18647 6616 19472 6644
rect 19981 6647 20039 6653
rect 18647 6613 18659 6616
rect 18601 6607 18659 6613
rect 19981 6613 19993 6647
rect 20027 6613 20039 6647
rect 19981 6607 20039 6613
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2682 6440 2688 6452
rect 2643 6412 2688 6440
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 8202 6440 8208 6452
rect 8163 6412 8208 6440
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 10502 6440 10508 6452
rect 9815 6412 10508 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10836 6412 10977 6440
rect 10836 6400 10842 6412
rect 10965 6409 10977 6412
rect 11011 6440 11023 6443
rect 11790 6440 11796 6452
rect 11011 6412 11796 6440
rect 11011 6409 11023 6412
rect 10965 6403 11023 6409
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 11974 6400 11980 6452
rect 12032 6440 12038 6452
rect 12032 6412 14780 6440
rect 12032 6400 12038 6412
rect 2866 6304 2872 6316
rect 2827 6276 2872 6304
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 3142 6304 3148 6316
rect 3103 6276 3148 6304
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 8220 6304 8248 6400
rect 9950 6372 9956 6384
rect 9600 6344 9956 6372
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8220 6276 8677 6304
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3007 6208 4292 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 2774 6128 2780 6180
rect 2832 6168 2838 6180
rect 4264 6177 4292 6208
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 7892 6208 8769 6236
rect 7892 6196 7898 6208
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 8864 6236 8892 6267
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9600 6313 9628 6344
rect 9950 6332 9956 6344
rect 10008 6372 10014 6384
rect 10229 6375 10287 6381
rect 10229 6372 10241 6375
rect 10008 6344 10241 6372
rect 10008 6332 10014 6344
rect 10229 6341 10241 6344
rect 10275 6341 10287 6375
rect 11882 6372 11888 6384
rect 11843 6344 11888 6372
rect 10229 6335 10287 6341
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 14366 6372 14372 6384
rect 12308 6344 14372 6372
rect 12308 6332 12314 6344
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 9088 6276 9413 6304
rect 9088 6264 9094 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6273 9643 6307
rect 11238 6304 11244 6316
rect 9585 6267 9643 6273
rect 10980 6276 11244 6304
rect 10980 6236 11008 6276
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 11848 6276 11893 6304
rect 11848 6264 11854 6276
rect 11974 6264 11980 6316
rect 12032 6313 12038 6316
rect 12032 6307 12061 6313
rect 12049 6273 12061 6307
rect 12032 6267 12061 6273
rect 12032 6264 12038 6267
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 13357 6307 13415 6313
rect 13357 6304 13369 6307
rect 12676 6276 13369 6304
rect 12676 6264 12682 6276
rect 13357 6273 13369 6276
rect 13403 6273 13415 6307
rect 13357 6267 13415 6273
rect 13725 6307 13783 6313
rect 13725 6273 13737 6307
rect 13771 6304 13783 6307
rect 13906 6304 13912 6316
rect 13771 6276 13912 6304
rect 13771 6273 13783 6276
rect 13725 6267 13783 6273
rect 13906 6264 13912 6276
rect 13964 6264 13970 6316
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 14056 6276 14565 6304
rect 14056 6264 14062 6276
rect 14553 6273 14565 6276
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 8864 6208 11008 6236
rect 8757 6199 8815 6205
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 12158 6236 12164 6248
rect 11112 6208 12164 6236
rect 11112 6196 11118 6208
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 13262 6236 13268 6248
rect 13223 6208 13268 6236
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 13924 6236 13952 6264
rect 14642 6236 14648 6248
rect 13924 6208 14648 6236
rect 14642 6196 14648 6208
rect 14700 6196 14706 6248
rect 3053 6171 3111 6177
rect 3053 6168 3065 6171
rect 2832 6140 3065 6168
rect 2832 6128 2838 6140
rect 3053 6137 3065 6140
rect 3099 6168 3111 6171
rect 4249 6171 4307 6177
rect 3099 6140 4016 6168
rect 3099 6137 3111 6140
rect 3053 6131 3111 6137
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3988 6100 4016 6140
rect 4249 6137 4261 6171
rect 4295 6168 4307 6171
rect 4338 6168 4344 6180
rect 4295 6140 4344 6168
rect 4295 6137 4307 6140
rect 4249 6131 4307 6137
rect 4338 6128 4344 6140
rect 4396 6168 4402 6180
rect 4706 6168 4712 6180
rect 4396 6140 4712 6168
rect 4396 6128 4402 6140
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 12802 6168 12808 6180
rect 6886 6140 12808 6168
rect 6886 6100 6914 6140
rect 12802 6128 12808 6140
rect 12860 6168 12866 6180
rect 13909 6171 13967 6177
rect 13909 6168 13921 6171
rect 12860 6140 13921 6168
rect 12860 6128 12866 6140
rect 13909 6137 13921 6140
rect 13955 6137 13967 6171
rect 13909 6131 13967 6137
rect 3988 6072 6914 6100
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9585 6103 9643 6109
rect 9585 6100 9597 6103
rect 9548 6072 9597 6100
rect 9548 6060 9554 6072
rect 9585 6069 9597 6072
rect 9631 6100 9643 6103
rect 10594 6100 10600 6112
rect 9631 6072 10600 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11480 6072 11529 6100
rect 11480 6060 11486 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 13630 6100 13636 6112
rect 11848 6072 13636 6100
rect 11848 6060 11854 6072
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13725 6103 13783 6109
rect 13725 6069 13737 6103
rect 13771 6100 13783 6103
rect 13814 6100 13820 6112
rect 13771 6072 13820 6100
rect 13771 6069 13783 6072
rect 13725 6063 13783 6069
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14752 6109 14780 6412
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 17586 6440 17592 6452
rect 16448 6412 17592 6440
rect 16448 6400 16454 6412
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18969 6443 19027 6449
rect 18969 6440 18981 6443
rect 18012 6412 18981 6440
rect 18012 6400 18018 6412
rect 18969 6409 18981 6412
rect 19015 6409 19027 6443
rect 19334 6440 19340 6452
rect 19295 6412 19340 6440
rect 18969 6403 19027 6409
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 20438 6440 20444 6452
rect 20399 6412 20444 6440
rect 20438 6400 20444 6412
rect 20496 6400 20502 6452
rect 22370 6440 22376 6452
rect 22331 6412 22376 6440
rect 22370 6400 22376 6412
rect 22428 6400 22434 6452
rect 28810 6440 28816 6452
rect 22572 6412 28816 6440
rect 15010 6372 15016 6384
rect 14971 6344 15016 6372
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 16482 6332 16488 6384
rect 16540 6372 16546 6384
rect 17221 6375 17279 6381
rect 17221 6372 17233 6375
rect 16540 6344 17233 6372
rect 16540 6332 16546 6344
rect 17221 6341 17233 6344
rect 17267 6341 17279 6375
rect 17221 6335 17279 6341
rect 17678 6332 17684 6384
rect 17736 6372 17742 6384
rect 18325 6375 18383 6381
rect 17736 6344 18282 6372
rect 17736 6332 17742 6344
rect 18254 6313 18282 6344
rect 18325 6341 18337 6375
rect 18371 6372 18383 6375
rect 20714 6372 20720 6384
rect 18371 6344 19334 6372
rect 18371 6341 18383 6344
rect 18325 6335 18383 6341
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18414 6304 18420 6316
rect 18375 6276 18420 6304
rect 18233 6267 18291 6273
rect 14936 6236 14964 6267
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 18892 6313 18920 6344
rect 19306 6316 19334 6344
rect 19996 6344 20720 6372
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6273 18935 6307
rect 19150 6304 19156 6316
rect 19111 6276 19156 6304
rect 18877 6267 18935 6273
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19306 6276 19340 6316
rect 19334 6264 19340 6276
rect 19392 6264 19398 6316
rect 19996 6313 20024 6344
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 20809 6375 20867 6381
rect 20809 6341 20821 6375
rect 20855 6372 20867 6375
rect 22572 6372 22600 6412
rect 28810 6400 28816 6412
rect 28868 6400 28874 6452
rect 22738 6372 22744 6384
rect 20855 6344 22600 6372
rect 22651 6344 22744 6372
rect 20855 6341 20867 6344
rect 20809 6335 20867 6341
rect 22738 6332 22744 6344
rect 22796 6372 22802 6384
rect 22796 6344 23428 6372
rect 22796 6332 22802 6344
rect 19981 6307 20039 6313
rect 19981 6273 19993 6307
rect 20027 6273 20039 6307
rect 20579 6307 20637 6313
rect 20579 6304 20591 6307
rect 19981 6267 20039 6273
rect 20272 6276 20591 6304
rect 19889 6239 19947 6245
rect 19889 6236 19901 6239
rect 14936 6208 19901 6236
rect 19889 6205 19901 6208
rect 19935 6205 19947 6239
rect 19889 6199 19947 6205
rect 15102 6128 15108 6180
rect 15160 6168 15166 6180
rect 20272 6168 20300 6276
rect 20579 6273 20591 6276
rect 20625 6273 20637 6307
rect 20579 6267 20637 6273
rect 20898 6264 20904 6316
rect 20956 6313 20962 6316
rect 20956 6307 20995 6313
rect 20983 6273 20995 6307
rect 20956 6267 20995 6273
rect 20956 6264 20962 6267
rect 21082 6264 21088 6316
rect 21140 6304 21146 6316
rect 22554 6304 22560 6316
rect 21140 6276 21185 6304
rect 22515 6276 22560 6304
rect 21140 6264 21146 6276
rect 22554 6264 22560 6276
rect 22612 6264 22618 6316
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6273 22891 6307
rect 22833 6267 22891 6273
rect 22002 6196 22008 6248
rect 22060 6236 22066 6248
rect 22848 6236 22876 6267
rect 22060 6208 22876 6236
rect 22060 6196 22066 6208
rect 15160 6140 20300 6168
rect 15160 6128 15166 6140
rect 14737 6103 14795 6109
rect 14737 6069 14749 6103
rect 14783 6100 14795 6103
rect 17218 6100 17224 6112
rect 14783 6072 17224 6100
rect 14783 6069 14795 6072
rect 14737 6063 14795 6069
rect 17218 6060 17224 6072
rect 17276 6060 17282 6112
rect 17313 6103 17371 6109
rect 17313 6069 17325 6103
rect 17359 6100 17371 6103
rect 17770 6100 17776 6112
rect 17359 6072 17776 6100
rect 17359 6069 17371 6072
rect 17313 6063 17371 6069
rect 17770 6060 17776 6072
rect 17828 6100 17834 6112
rect 18414 6100 18420 6112
rect 17828 6072 18420 6100
rect 17828 6060 17834 6072
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 23400 6109 23428 6344
rect 23385 6103 23443 6109
rect 23385 6069 23397 6103
rect 23431 6100 23443 6103
rect 37826 6100 37832 6112
rect 23431 6072 37832 6100
rect 23431 6069 23443 6072
rect 23385 6063 23443 6069
rect 37826 6060 37832 6072
rect 37884 6060 37890 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 5776 5868 7389 5896
rect 5776 5856 5782 5868
rect 7377 5865 7389 5868
rect 7423 5865 7435 5899
rect 9030 5896 9036 5908
rect 8991 5868 9036 5896
rect 7377 5859 7435 5865
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 12434 5896 12440 5908
rect 9140 5868 12440 5896
rect 7926 5760 7932 5772
rect 7760 5732 7932 5760
rect 7760 5701 7788 5732
rect 7926 5720 7932 5732
rect 7984 5760 7990 5772
rect 9048 5760 9076 5856
rect 7984 5732 9076 5760
rect 7984 5720 7990 5732
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 7668 5624 7696 5655
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 7892 5664 7937 5692
rect 7892 5652 7898 5664
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8076 5664 8121 5692
rect 8076 5652 8082 5664
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8260 5664 9045 5692
rect 8260 5652 8266 5664
rect 9033 5661 9045 5664
rect 9079 5692 9091 5695
rect 9140 5692 9168 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12618 5896 12624 5908
rect 12544 5868 12624 5896
rect 10413 5831 10471 5837
rect 10413 5797 10425 5831
rect 10459 5828 10471 5831
rect 12544 5828 12572 5868
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 13630 5856 13636 5908
rect 13688 5896 13694 5908
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 13688 5868 14381 5896
rect 13688 5856 13694 5868
rect 14369 5865 14381 5868
rect 14415 5896 14427 5899
rect 15010 5896 15016 5908
rect 14415 5868 15016 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 19705 5899 19763 5905
rect 19705 5865 19717 5899
rect 19751 5896 19763 5899
rect 20346 5896 20352 5908
rect 19751 5868 20352 5896
rect 19751 5865 19763 5868
rect 19705 5859 19763 5865
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 20441 5899 20499 5905
rect 20441 5865 20453 5899
rect 20487 5896 20499 5899
rect 20714 5896 20720 5908
rect 20487 5868 20720 5896
rect 20487 5865 20499 5868
rect 20441 5859 20499 5865
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 10459 5800 12572 5828
rect 10459 5797 10471 5800
rect 10413 5791 10471 5797
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 9456 5732 10517 5760
rect 9456 5720 9462 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 9079 5664 9168 5692
rect 9217 5695 9275 5701
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9306 5692 9312 5704
rect 9263 5664 9312 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 10226 5692 10232 5704
rect 10187 5664 10232 5692
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10520 5692 10548 5723
rect 10594 5720 10600 5772
rect 10652 5760 10658 5772
rect 11974 5760 11980 5772
rect 10652 5732 11980 5760
rect 10652 5720 10658 5732
rect 11974 5720 11980 5732
rect 12032 5720 12038 5772
rect 12158 5720 12164 5772
rect 12216 5760 12222 5772
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 12216 5732 12357 5760
rect 12216 5720 12222 5732
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12492 5732 12541 5760
rect 12492 5720 12498 5732
rect 12529 5729 12541 5732
rect 12575 5760 12587 5763
rect 15194 5760 15200 5772
rect 12575 5732 15200 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 11149 5695 11207 5701
rect 11149 5692 11161 5695
rect 10520 5664 11161 5692
rect 11149 5661 11161 5664
rect 11195 5661 11207 5695
rect 11422 5692 11428 5704
rect 11383 5664 11428 5692
rect 11149 5655 11207 5661
rect 9582 5624 9588 5636
rect 7668 5596 9588 5624
rect 9582 5584 9588 5596
rect 9640 5584 9646 5636
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 10965 5627 11023 5633
rect 10965 5624 10977 5627
rect 10928 5596 10977 5624
rect 10928 5584 10934 5596
rect 10965 5593 10977 5596
rect 11011 5593 11023 5627
rect 10965 5587 11023 5593
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 10045 5559 10103 5565
rect 10045 5556 10057 5559
rect 8352 5528 10057 5556
rect 8352 5516 8358 5528
rect 10045 5525 10057 5528
rect 10091 5525 10103 5559
rect 11164 5556 11192 5655
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11609 5695 11667 5701
rect 11609 5661 11621 5695
rect 11655 5692 11667 5695
rect 12250 5692 12256 5704
rect 11655 5664 12256 5692
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5692 12679 5695
rect 14090 5692 14096 5704
rect 12667 5664 14096 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 11238 5584 11244 5636
rect 11296 5624 11302 5636
rect 12636 5624 12664 5655
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 19334 5692 19340 5704
rect 19291 5664 19340 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5661 19579 5695
rect 20254 5692 20260 5704
rect 20215 5664 20260 5692
rect 19521 5655 19579 5661
rect 11296 5596 12664 5624
rect 11296 5584 11302 5596
rect 19058 5584 19064 5636
rect 19116 5624 19122 5636
rect 19536 5624 19564 5655
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 19116 5596 19564 5624
rect 19116 5584 19122 5596
rect 13906 5556 13912 5568
rect 11164 5528 13912 5556
rect 10045 5519 10103 5525
rect 13906 5516 13912 5528
rect 13964 5516 13970 5568
rect 19337 5559 19395 5565
rect 19337 5525 19349 5559
rect 19383 5556 19395 5559
rect 19426 5556 19432 5568
rect 19383 5528 19432 5556
rect 19383 5525 19395 5528
rect 19337 5519 19395 5525
rect 19426 5516 19432 5528
rect 19484 5516 19490 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 6362 5352 6368 5364
rect 6323 5324 6368 5352
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 7282 5352 7288 5364
rect 7243 5324 7288 5352
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 7708 5324 8309 5352
rect 7708 5312 7714 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 18230 5352 18236 5364
rect 18191 5324 18236 5352
rect 8297 5315 8355 5321
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 20622 5312 20628 5364
rect 20680 5352 20686 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 20680 5324 21833 5352
rect 20680 5312 20686 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 22002 5312 22008 5364
rect 22060 5312 22066 5364
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 17310 5284 17316 5296
rect 3384 5256 17316 5284
rect 3384 5244 3390 5256
rect 17310 5244 17316 5256
rect 17368 5284 17374 5296
rect 17497 5287 17555 5293
rect 17497 5284 17509 5287
rect 17368 5256 17509 5284
rect 17368 5244 17374 5256
rect 17497 5253 17509 5256
rect 17543 5253 17555 5287
rect 17497 5247 17555 5253
rect 21358 5244 21364 5296
rect 21416 5284 21422 5296
rect 22020 5284 22048 5312
rect 21416 5256 22324 5284
rect 21416 5244 21422 5256
rect 6546 5216 6552 5228
rect 6507 5188 6552 5216
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 6886 5188 7573 5216
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6886 5148 6914 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 8294 5216 8300 5228
rect 7791 5188 8300 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19889 5219 19947 5225
rect 19889 5216 19901 5219
rect 19392 5188 19901 5216
rect 19392 5176 19398 5188
rect 19889 5185 19901 5188
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 22005 5219 22063 5225
rect 22005 5185 22017 5219
rect 22051 5216 22063 5219
rect 22094 5216 22100 5228
rect 22051 5188 22100 5216
rect 22051 5185 22063 5188
rect 22005 5179 22063 5185
rect 22094 5176 22100 5188
rect 22152 5176 22158 5228
rect 22296 5225 22324 5256
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5185 22247 5219
rect 22189 5179 22247 5185
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 24762 5216 24768 5228
rect 22327 5188 24768 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 6788 5120 6914 5148
rect 7469 5151 7527 5157
rect 6788 5108 6794 5120
rect 7469 5117 7481 5151
rect 7515 5117 7527 5151
rect 7650 5148 7656 5160
rect 7611 5120 7656 5148
rect 7469 5111 7527 5117
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7484 5080 7512 5111
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 22204 5148 22232 5179
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 15436 5120 22232 5148
rect 15436 5108 15442 5120
rect 7834 5080 7840 5092
rect 7156 5052 7840 5080
rect 7156 5040 7162 5052
rect 7834 5040 7840 5052
rect 7892 5040 7898 5092
rect 20073 5083 20131 5089
rect 20073 5049 20085 5083
rect 20119 5080 20131 5083
rect 20530 5080 20536 5092
rect 20119 5052 20536 5080
rect 20119 5049 20131 5052
rect 20073 5043 20131 5049
rect 20530 5040 20536 5052
rect 20588 5080 20594 5092
rect 20898 5080 20904 5092
rect 20588 5052 20904 5080
rect 20588 5040 20594 5052
rect 20898 5040 20904 5052
rect 20956 5040 20962 5092
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 10226 5012 10232 5024
rect 9999 4984 10232 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 10226 4972 10232 4984
rect 10284 5012 10290 5024
rect 16761 5015 16819 5021
rect 16761 5012 16773 5015
rect 10284 4984 16773 5012
rect 10284 4972 10290 4984
rect 16761 4981 16773 4984
rect 16807 5012 16819 5015
rect 17034 5012 17040 5024
rect 16807 4984 17040 5012
rect 16807 4981 16819 4984
rect 16761 4975 16819 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1946 4768 1952 4820
rect 2004 4808 2010 4820
rect 6089 4811 6147 4817
rect 6089 4808 6101 4811
rect 2004 4780 6101 4808
rect 2004 4768 2010 4780
rect 6089 4777 6101 4780
rect 6135 4777 6147 4811
rect 6089 4771 6147 4777
rect 6104 4604 6132 4771
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 7708 4780 9597 4808
rect 7708 4768 7714 4780
rect 9585 4777 9597 4780
rect 9631 4808 9643 4811
rect 9674 4808 9680 4820
rect 9631 4780 9680 4808
rect 9631 4777 9643 4780
rect 9585 4771 9643 4777
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 10134 4808 10140 4820
rect 10095 4780 10140 4808
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 18782 4808 18788 4820
rect 17819 4780 18788 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 20162 4808 20168 4820
rect 20123 4780 20168 4808
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 21821 4811 21879 4817
rect 21821 4777 21833 4811
rect 21867 4808 21879 4811
rect 21910 4808 21916 4820
rect 21867 4780 21916 4808
rect 21867 4777 21879 4780
rect 21821 4771 21879 4777
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 23474 4808 23480 4820
rect 23435 4780 23480 4808
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 24394 4808 24400 4820
rect 24355 4780 24400 4808
rect 24394 4768 24400 4780
rect 24452 4768 24458 4820
rect 6914 4740 6920 4752
rect 6656 4712 6920 4740
rect 6656 4613 6684 4712
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 15102 4740 15108 4752
rect 7340 4712 15108 4740
rect 7340 4700 7346 4712
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 18693 4743 18751 4749
rect 15212 4712 18460 4740
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 6788 4644 7941 4672
rect 6788 4632 6794 4644
rect 6840 4613 6868 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 10686 4672 10692 4684
rect 7929 4635 7987 4641
rect 10336 4644 10692 4672
rect 6641 4607 6699 4613
rect 6641 4604 6653 4607
rect 6104 4576 6653 4604
rect 6641 4573 6653 4576
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 7009 4607 7067 4613
rect 6871 4576 6905 4604
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 7834 4604 7840 4616
rect 7055 4576 7840 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 9490 4604 9496 4616
rect 8067 4576 9496 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 10336 4613 10364 4644
rect 10686 4632 10692 4644
rect 10744 4632 10750 4684
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4573 10379 4607
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10321 4567 10379 4573
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 6917 4539 6975 4545
rect 6917 4505 6929 4539
rect 6963 4536 6975 4539
rect 7374 4536 7380 4548
rect 6963 4508 7380 4536
rect 6963 4505 6975 4508
rect 6917 4499 6975 4505
rect 7024 4480 7052 4508
rect 7374 4496 7380 4508
rect 7432 4536 7438 4548
rect 10612 4536 10640 4567
rect 15102 4564 15108 4616
rect 15160 4604 15166 4616
rect 15212 4604 15240 4712
rect 15838 4632 15844 4684
rect 15896 4672 15902 4684
rect 18432 4672 18460 4712
rect 18693 4709 18705 4743
rect 18739 4740 18751 4743
rect 18874 4740 18880 4752
rect 18739 4712 18880 4740
rect 18739 4709 18751 4712
rect 18693 4703 18751 4709
rect 18874 4700 18880 4712
rect 18932 4700 18938 4752
rect 15896 4644 18368 4672
rect 18432 4644 19840 4672
rect 15896 4632 15902 4644
rect 15160 4576 15240 4604
rect 15381 4607 15439 4613
rect 15160 4564 15166 4576
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 16574 4604 16580 4616
rect 15427 4576 16580 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 16574 4564 16580 4576
rect 16632 4564 16638 4616
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 17276 4576 17325 4604
rect 17276 4564 17282 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 18340 4613 18368 4644
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 17460 4576 17601 4604
rect 17460 4564 17466 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 18233 4607 18291 4613
rect 18233 4573 18245 4607
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4573 18383 4607
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18325 4567 18383 4573
rect 11054 4536 11060 4548
rect 7432 4508 11060 4536
rect 7432 4496 7438 4508
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 11149 4539 11207 4545
rect 11149 4505 11161 4539
rect 11195 4536 11207 4539
rect 11882 4536 11888 4548
rect 11195 4508 11888 4536
rect 11195 4505 11207 4508
rect 11149 4499 11207 4505
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 16482 4496 16488 4548
rect 16540 4536 16546 4548
rect 16540 4508 17448 4536
rect 16540 4496 16546 4508
rect 7006 4428 7012 4480
rect 7064 4428 7070 4480
rect 7190 4468 7196 4480
rect 7151 4440 7196 4468
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 11698 4468 11704 4480
rect 11659 4440 11704 4468
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 15654 4428 15660 4480
rect 15712 4468 15718 4480
rect 15841 4471 15899 4477
rect 15841 4468 15853 4471
rect 15712 4440 15853 4468
rect 15712 4428 15718 4440
rect 15841 4437 15853 4440
rect 15887 4437 15899 4471
rect 15841 4431 15899 4437
rect 16666 4428 16672 4480
rect 16724 4468 16730 4480
rect 17420 4477 17448 4508
rect 17494 4496 17500 4548
rect 17552 4536 17558 4548
rect 18248 4536 18276 4567
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 19812 4613 19840 4644
rect 20162 4632 20168 4684
rect 20220 4672 20226 4684
rect 20346 4672 20352 4684
rect 20220 4644 20352 4672
rect 20220 4632 20226 4644
rect 20346 4632 20352 4644
rect 20404 4632 20410 4684
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4573 19855 4607
rect 19978 4604 19984 4616
rect 19939 4576 19984 4604
rect 19797 4567 19855 4573
rect 19720 4536 19748 4567
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 21358 4604 21364 4616
rect 21271 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 21637 4607 21695 4613
rect 21637 4573 21649 4607
rect 21683 4604 21695 4607
rect 22094 4604 22100 4616
rect 21683 4576 22100 4604
rect 21683 4573 21695 4576
rect 21637 4567 21695 4573
rect 22094 4564 22100 4576
rect 22152 4564 22158 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24581 4567 24639 4573
rect 21376 4536 21404 4564
rect 17552 4508 21404 4536
rect 24596 4536 24624 4567
rect 24762 4564 24768 4616
rect 24820 4604 24826 4616
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 24820 4576 24869 4604
rect 24820 4564 24826 4576
rect 24857 4573 24869 4576
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 24946 4536 24952 4548
rect 24596 4508 24952 4536
rect 17552 4496 17558 4508
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 16761 4471 16819 4477
rect 16761 4468 16773 4471
rect 16724 4440 16773 4468
rect 16724 4428 16730 4440
rect 16761 4437 16773 4440
rect 16807 4437 16819 4471
rect 16761 4431 16819 4437
rect 17405 4471 17463 4477
rect 17405 4437 17417 4471
rect 17451 4437 17463 4471
rect 21450 4468 21456 4480
rect 21411 4440 21456 4468
rect 17405 4431 17463 4437
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 21910 4428 21916 4480
rect 21968 4468 21974 4480
rect 22925 4471 22983 4477
rect 22925 4468 22937 4471
rect 21968 4440 22937 4468
rect 21968 4428 21974 4440
rect 22925 4437 22937 4440
rect 22971 4468 22983 4471
rect 23198 4468 23204 4480
rect 22971 4440 23204 4468
rect 22971 4437 22983 4440
rect 22925 4431 22983 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4468 24823 4471
rect 34422 4468 34428 4480
rect 24811 4440 34428 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 34422 4428 34428 4440
rect 34480 4428 34486 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 6546 4224 6552 4276
rect 6604 4264 6610 4276
rect 6733 4267 6791 4273
rect 6733 4264 6745 4267
rect 6604 4236 6745 4264
rect 6604 4224 6610 4236
rect 6733 4233 6745 4236
rect 6779 4233 6791 4267
rect 6733 4227 6791 4233
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 12161 4267 12219 4273
rect 6972 4236 9352 4264
rect 6972 4224 6978 4236
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7190 4128 7196 4140
rect 6963 4100 7196 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 9324 4137 9352 4236
rect 12161 4233 12173 4267
rect 12207 4264 12219 4267
rect 12250 4264 12256 4276
rect 12207 4236 12256 4264
rect 12207 4233 12219 4236
rect 12161 4227 12219 4233
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 17494 4264 17500 4276
rect 17276 4236 17500 4264
rect 17276 4224 17282 4236
rect 17494 4224 17500 4236
rect 17552 4224 17558 4276
rect 17678 4224 17684 4276
rect 17736 4224 17742 4276
rect 22094 4224 22100 4276
rect 22152 4264 22158 4276
rect 22152 4236 22197 4264
rect 22152 4224 22158 4236
rect 23566 4224 23572 4276
rect 23624 4224 23630 4276
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 17589 4199 17647 4205
rect 9732 4168 10180 4196
rect 9732 4156 9738 4168
rect 10152 4137 10180 4168
rect 17589 4165 17601 4199
rect 17635 4196 17647 4199
rect 17696 4196 17724 4224
rect 18046 4196 18052 4208
rect 17635 4168 18052 4196
rect 17635 4165 17647 4168
rect 17589 4159 17647 4165
rect 18046 4156 18052 4168
rect 18104 4196 18110 4208
rect 18785 4199 18843 4205
rect 18785 4196 18797 4199
rect 18104 4168 18797 4196
rect 18104 4156 18110 4168
rect 18785 4165 18797 4168
rect 18831 4165 18843 4199
rect 18785 4159 18843 4165
rect 18966 4156 18972 4208
rect 19024 4196 19030 4208
rect 22002 4196 22008 4208
rect 19024 4168 22008 4196
rect 19024 4156 19030 4168
rect 22002 4156 22008 4168
rect 22060 4156 22066 4208
rect 23106 4156 23112 4208
rect 23164 4196 23170 4208
rect 23477 4199 23535 4205
rect 23164 4168 23428 4196
rect 23164 4156 23170 4168
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9355 4100 10057 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4128 10287 4131
rect 10413 4131 10471 4137
rect 10275 4100 10364 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 7098 4060 7104 4072
rect 7059 4032 7104 4060
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9640 4032 9781 4060
rect 9640 4020 9646 4032
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 10060 4060 10088 4091
rect 10060 4032 10180 4060
rect 9769 4023 9827 4029
rect 8757 3995 8815 4001
rect 8757 3961 8769 3995
rect 8803 3992 8815 3995
rect 9490 3992 9496 4004
rect 8803 3964 9496 3992
rect 8803 3961 8815 3964
rect 8757 3955 8815 3961
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 5442 3924 5448 3936
rect 5399 3896 5448 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 8202 3924 8208 3936
rect 8163 3896 8208 3924
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 10152 3924 10180 4032
rect 10336 3992 10364 4100
rect 10413 4097 10425 4131
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10428 4060 10456 4091
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 12002 4131 12060 4137
rect 12002 4128 12014 4131
rect 10744 4100 12014 4128
rect 10744 4088 10750 4100
rect 12002 4097 12014 4100
rect 12048 4097 12060 4131
rect 12002 4091 12060 4097
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 13320 4100 15117 4128
rect 13320 4088 13326 4100
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 15289 4131 15347 4137
rect 15289 4128 15301 4131
rect 15252 4100 15301 4128
rect 15252 4088 15258 4100
rect 15289 4097 15301 4100
rect 15335 4097 15347 4131
rect 15289 4091 15347 4097
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4128 15623 4131
rect 15654 4128 15660 4140
rect 15611 4100 15660 4128
rect 15611 4097 15623 4100
rect 15565 4091 15623 4097
rect 10428 4032 11008 4060
rect 10594 3992 10600 4004
rect 10336 3964 10600 3992
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10778 3924 10784 3936
rect 10152 3896 10784 3924
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 10980 3933 11008 4032
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 11517 4063 11575 4069
rect 11517 4060 11529 4063
rect 11112 4032 11529 4060
rect 11112 4020 11118 4032
rect 11517 4029 11529 4032
rect 11563 4029 11575 4063
rect 11790 4060 11796 4072
rect 11751 4032 11796 4060
rect 11517 4023 11575 4029
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12713 4063 12771 4069
rect 12713 4060 12725 4063
rect 11940 4032 12725 4060
rect 11940 4020 11946 4032
rect 12713 4029 12725 4032
rect 12759 4060 12771 4063
rect 15580 4060 15608 4091
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 15746 4088 15752 4140
rect 15804 4128 15810 4140
rect 15804 4100 15849 4128
rect 15804 4088 15810 4100
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 16816 4100 17509 4128
rect 16816 4088 16822 4100
rect 17497 4097 17509 4100
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 17681 4131 17739 4137
rect 17681 4097 17693 4131
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 12759 4032 15608 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 17126 4020 17132 4072
rect 17184 4060 17190 4072
rect 17696 4060 17724 4091
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 17828 4100 17877 4128
rect 17828 4088 17834 4100
rect 17865 4097 17877 4100
rect 17911 4128 17923 4131
rect 18509 4131 18567 4137
rect 18509 4128 18521 4131
rect 17911 4100 18521 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18509 4097 18521 4100
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 17184 4032 17724 4060
rect 17184 4020 17190 4032
rect 12250 3952 12256 4004
rect 12308 3992 12314 4004
rect 13173 3995 13231 4001
rect 13173 3992 13185 3995
rect 12308 3964 13185 3992
rect 12308 3952 12314 3964
rect 13173 3961 13185 3964
rect 13219 3961 13231 3995
rect 13173 3955 13231 3961
rect 14645 3995 14703 4001
rect 14645 3961 14657 3995
rect 14691 3992 14703 3995
rect 15286 3992 15292 4004
rect 14691 3964 15292 3992
rect 14691 3961 14703 3964
rect 14645 3955 14703 3961
rect 15286 3952 15292 3964
rect 15344 3952 15350 4004
rect 15381 3995 15439 4001
rect 15381 3961 15393 3995
rect 15427 3961 15439 3995
rect 15381 3955 15439 3961
rect 15473 3995 15531 4001
rect 15473 3961 15485 3995
rect 15519 3992 15531 3995
rect 15562 3992 15568 4004
rect 15519 3964 15568 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11238 3924 11244 3936
rect 11011 3896 11244 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11238 3884 11244 3896
rect 11296 3924 11302 3936
rect 11882 3924 11888 3936
rect 11296 3896 11888 3924
rect 11296 3884 11302 3896
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 15396 3924 15424 3955
rect 15562 3952 15568 3964
rect 15620 3952 15626 4004
rect 16853 3995 16911 4001
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 16942 3992 16948 4004
rect 16899 3964 16948 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 16942 3952 16948 3964
rect 17000 3952 17006 4004
rect 17313 3995 17371 4001
rect 17313 3961 17325 3995
rect 17359 3992 17371 3995
rect 17586 3992 17592 4004
rect 17359 3964 17592 3992
rect 17359 3961 17371 3964
rect 17313 3955 17371 3961
rect 17586 3952 17592 3964
rect 17644 3952 17650 4004
rect 18708 3992 18736 4091
rect 18874 4088 18880 4140
rect 18932 4128 18938 4140
rect 19613 4131 19671 4137
rect 18932 4100 18977 4128
rect 18932 4088 18938 4100
rect 19613 4097 19625 4131
rect 19659 4128 19671 4131
rect 22094 4128 22100 4140
rect 19659 4100 22100 4128
rect 19659 4097 19671 4100
rect 19613 4091 19671 4097
rect 19628 4060 19656 4091
rect 22094 4088 22100 4100
rect 22152 4088 22158 4140
rect 22278 4128 22284 4140
rect 22239 4100 22284 4128
rect 22278 4088 22284 4100
rect 22336 4088 22342 4140
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4097 22431 4131
rect 22373 4091 22431 4097
rect 18892 4032 19656 4060
rect 18892 3992 18920 4032
rect 21818 4020 21824 4072
rect 21876 4060 21882 4072
rect 22388 4060 22416 4091
rect 22462 4088 22468 4140
rect 22520 4128 22526 4140
rect 22649 4131 22707 4137
rect 22520 4100 22565 4128
rect 22520 4088 22526 4100
rect 22649 4097 22661 4131
rect 22695 4128 22707 4131
rect 22922 4128 22928 4140
rect 22695 4100 22928 4128
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 22922 4088 22928 4100
rect 22980 4088 22986 4140
rect 23198 4088 23204 4140
rect 23256 4137 23262 4140
rect 23400 4137 23428 4168
rect 23477 4165 23489 4199
rect 23523 4196 23535 4199
rect 23584 4196 23612 4224
rect 23523 4168 23612 4196
rect 23523 4165 23535 4168
rect 23477 4159 23535 4165
rect 23750 4156 23756 4208
rect 23808 4196 23814 4208
rect 33318 4196 33324 4208
rect 23808 4168 33324 4196
rect 23808 4156 23814 4168
rect 33318 4156 33324 4168
rect 33376 4156 33382 4208
rect 23256 4131 23305 4137
rect 23256 4097 23259 4131
rect 23293 4097 23305 4131
rect 23256 4091 23305 4097
rect 23361 4131 23428 4137
rect 23361 4097 23373 4131
rect 23407 4100 23428 4131
rect 23661 4131 23719 4137
rect 23407 4097 23419 4100
rect 23361 4091 23419 4097
rect 23661 4097 23673 4131
rect 23707 4097 23719 4131
rect 24118 4128 24124 4140
rect 24079 4100 24124 4128
rect 23661 4091 23719 4097
rect 23256 4088 23262 4091
rect 22738 4060 22744 4072
rect 21876 4032 22416 4060
rect 22480 4032 22744 4060
rect 21876 4020 21882 4032
rect 19058 3992 19064 4004
rect 18708 3964 18920 3992
rect 19019 3964 19064 3992
rect 19058 3952 19064 3964
rect 19116 3952 19122 4004
rect 22480 3992 22508 4032
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 22940 4060 22968 4088
rect 23676 4060 23704 4091
rect 24118 4088 24124 4100
rect 24176 4088 24182 4140
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4128 24363 4131
rect 24394 4128 24400 4140
rect 24351 4100 24400 4128
rect 24351 4097 24363 4100
rect 24305 4091 24363 4097
rect 24394 4088 24400 4100
rect 24452 4088 24458 4140
rect 24489 4131 24547 4137
rect 24489 4097 24501 4131
rect 24535 4097 24547 4131
rect 24489 4091 24547 4097
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4128 24639 4131
rect 24762 4128 24768 4140
rect 24627 4100 24768 4128
rect 24627 4097 24639 4100
rect 24581 4091 24639 4097
rect 22940 4032 23704 4060
rect 24504 4060 24532 4091
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 25590 4128 25596 4140
rect 25551 4100 25596 4128
rect 25590 4088 25596 4100
rect 25648 4088 25654 4140
rect 26234 4128 26240 4140
rect 26195 4100 26240 4128
rect 26234 4088 26240 4100
rect 26292 4088 26298 4140
rect 36630 4128 36636 4140
rect 31726 4100 36636 4128
rect 31726 4060 31754 4100
rect 36630 4088 36636 4100
rect 36688 4088 36694 4140
rect 24504 4032 31754 4060
rect 19168 3964 22508 3992
rect 16114 3924 16120 3936
rect 15396 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 19168 3924 19196 3964
rect 22554 3952 22560 4004
rect 22612 3992 22618 4004
rect 23109 3995 23167 4001
rect 23109 3992 23121 3995
rect 22612 3964 23121 3992
rect 22612 3952 22618 3964
rect 23109 3961 23121 3964
rect 23155 3961 23167 3995
rect 23109 3955 23167 3961
rect 16356 3896 19196 3924
rect 16356 3884 16362 3896
rect 19794 3884 19800 3936
rect 19852 3924 19858 3936
rect 20073 3927 20131 3933
rect 20073 3924 20085 3927
rect 19852 3896 20085 3924
rect 19852 3884 19858 3896
rect 20073 3893 20085 3896
rect 20119 3924 20131 3927
rect 20622 3924 20628 3936
rect 20119 3896 20628 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 20622 3884 20628 3896
rect 20680 3884 20686 3936
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 22646 3924 22652 3936
rect 22152 3896 22652 3924
rect 22152 3884 22158 3896
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 24762 3884 24768 3936
rect 24820 3924 24826 3936
rect 25041 3927 25099 3933
rect 25041 3924 25053 3927
rect 24820 3896 25053 3924
rect 24820 3884 24826 3896
rect 25041 3893 25053 3896
rect 25087 3893 25099 3927
rect 25041 3887 25099 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9674 3720 9680 3732
rect 9539 3692 9680 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 11977 3723 12035 3729
rect 11977 3720 11989 3723
rect 11940 3692 11989 3720
rect 11940 3680 11946 3692
rect 11977 3689 11989 3692
rect 12023 3689 12035 3723
rect 15378 3720 15384 3732
rect 15339 3692 15384 3720
rect 11977 3683 12035 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15562 3720 15568 3732
rect 15523 3692 15568 3720
rect 15562 3680 15568 3692
rect 15620 3680 15626 3732
rect 16114 3720 16120 3732
rect 16075 3692 16120 3720
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16482 3720 16488 3732
rect 16264 3692 16488 3720
rect 16264 3680 16270 3692
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 17129 3723 17187 3729
rect 17129 3689 17141 3723
rect 17175 3720 17187 3723
rect 17402 3720 17408 3732
rect 17175 3692 17408 3720
rect 17175 3689 17187 3692
rect 17129 3683 17187 3689
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 19150 3720 19156 3732
rect 18739 3692 19156 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 19150 3680 19156 3692
rect 19208 3680 19214 3732
rect 19426 3720 19432 3732
rect 19260 3692 19432 3720
rect 15746 3652 15752 3664
rect 10980 3624 11836 3652
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3584 7895 3587
rect 8386 3584 8392 3596
rect 7883 3556 8392 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 10594 3544 10600 3596
rect 10652 3584 10658 3596
rect 10980 3593 11008 3624
rect 11808 3596 11836 3624
rect 12406 3624 15752 3652
rect 10965 3587 11023 3593
rect 10965 3584 10977 3587
rect 10652 3556 10977 3584
rect 10652 3544 10658 3556
rect 10965 3553 10977 3556
rect 11011 3553 11023 3587
rect 10965 3547 11023 3553
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 6181 3519 6239 3525
rect 6181 3485 6193 3519
rect 6227 3516 6239 3519
rect 6730 3516 6736 3528
rect 6227 3488 6736 3516
rect 6227 3485 6239 3488
rect 6181 3479 6239 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 9674 3476 9680 3528
rect 9732 3516 9738 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9732 3488 10425 3516
rect 9732 3476 9738 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3516 10747 3519
rect 10778 3516 10784 3528
rect 10735 3488 10784 3516
rect 10735 3485 10747 3488
rect 10689 3479 10747 3485
rect 7285 3451 7343 3457
rect 7285 3417 7297 3451
rect 7331 3448 7343 3451
rect 7834 3448 7840 3460
rect 7331 3420 7840 3448
rect 7331 3417 7343 3420
rect 7285 3411 7343 3417
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 8389 3451 8447 3457
rect 8389 3417 8401 3451
rect 8435 3448 8447 3451
rect 10704 3448 10732 3479
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 11238 3516 11244 3528
rect 11199 3488 11244 3516
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11532 3516 11560 3547
rect 11790 3544 11796 3596
rect 11848 3584 11854 3596
rect 12406 3584 12434 3624
rect 15746 3612 15752 3624
rect 15804 3612 15810 3664
rect 16942 3652 16948 3664
rect 16500 3624 16948 3652
rect 11848 3556 12434 3584
rect 15289 3587 15347 3593
rect 11848 3544 11854 3556
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15838 3584 15844 3596
rect 15335 3556 15844 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16500 3593 16528 3624
rect 16942 3612 16948 3624
rect 17000 3652 17006 3664
rect 19260 3652 19288 3692
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 19978 3720 19984 3732
rect 19939 3692 19984 3720
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20993 3723 21051 3729
rect 20993 3720 21005 3723
rect 20864 3692 21005 3720
rect 20864 3680 20870 3692
rect 20993 3689 21005 3692
rect 21039 3689 21051 3723
rect 21542 3720 21548 3732
rect 21503 3692 21548 3720
rect 20993 3683 21051 3689
rect 21542 3680 21548 3692
rect 21600 3680 21606 3732
rect 22094 3720 22100 3732
rect 21652 3692 22100 3720
rect 17000 3624 19288 3652
rect 19337 3655 19395 3661
rect 17000 3612 17006 3624
rect 19337 3621 19349 3655
rect 19383 3652 19395 3655
rect 21652 3652 21680 3692
rect 22094 3680 22100 3692
rect 22152 3680 22158 3732
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 23569 3723 23627 3729
rect 23569 3720 23581 3723
rect 22796 3692 23581 3720
rect 22796 3680 22802 3692
rect 23569 3689 23581 3692
rect 23615 3689 23627 3723
rect 24946 3720 24952 3732
rect 24907 3692 24952 3720
rect 23569 3683 23627 3689
rect 24946 3680 24952 3692
rect 25004 3680 25010 3732
rect 26510 3720 26516 3732
rect 26471 3692 26516 3720
rect 26510 3680 26516 3692
rect 26568 3680 26574 3732
rect 27062 3720 27068 3732
rect 27023 3692 27068 3720
rect 27062 3680 27068 3692
rect 27120 3680 27126 3732
rect 27614 3720 27620 3732
rect 27575 3692 27620 3720
rect 27614 3680 27620 3692
rect 27672 3680 27678 3732
rect 36630 3720 36636 3732
rect 36591 3692 36636 3720
rect 36630 3680 36636 3692
rect 36688 3680 36694 3732
rect 19383 3624 21680 3652
rect 19383 3621 19395 3624
rect 19337 3615 19395 3621
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3553 16543 3587
rect 17954 3584 17960 3596
rect 16485 3547 16543 3553
rect 16592 3556 17960 3584
rect 11974 3516 11980 3528
rect 11532 3488 11980 3516
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 15102 3516 15108 3528
rect 15063 3488 15108 3516
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 16114 3516 16120 3528
rect 15427 3488 16120 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 8435 3420 10732 3448
rect 8435 3417 8447 3420
rect 8389 3411 8447 3417
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 15396 3448 15424 3479
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 16298 3516 16304 3528
rect 16259 3488 16304 3516
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16390 3476 16396 3528
rect 16448 3516 16454 3528
rect 16592 3525 16620 3556
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 19352 3584 19380 3615
rect 21726 3612 21732 3664
rect 21784 3652 21790 3664
rect 22557 3655 22615 3661
rect 22557 3652 22569 3655
rect 21784 3624 22569 3652
rect 21784 3612 21790 3624
rect 22557 3621 22569 3624
rect 22603 3621 22615 3655
rect 22557 3615 22615 3621
rect 18340 3556 19380 3584
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 16448 3488 16589 3516
rect 16448 3476 16454 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 16850 3476 16856 3528
rect 16908 3516 16914 3528
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 16908 3488 17325 3516
rect 16908 3476 16914 3488
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 17313 3479 17371 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 17770 3516 17776 3528
rect 17727 3488 17776 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 17770 3476 17776 3488
rect 17828 3516 17834 3528
rect 18340 3525 18368 3556
rect 21542 3544 21548 3596
rect 21600 3584 21606 3596
rect 22370 3584 22376 3596
rect 21600 3556 21956 3584
rect 21600 3544 21606 3556
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17828 3488 18153 3516
rect 17828 3476 17834 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 13688 3420 15424 3448
rect 17405 3451 17463 3457
rect 13688 3408 13694 3420
rect 17405 3417 17417 3451
rect 17451 3448 17463 3451
rect 18046 3448 18052 3460
rect 17451 3420 18052 3448
rect 17451 3417 17463 3420
rect 17405 3411 17463 3417
rect 18046 3408 18052 3420
rect 18104 3448 18110 3460
rect 18417 3451 18475 3457
rect 18417 3448 18429 3451
rect 18104 3420 18429 3448
rect 18104 3408 18110 3420
rect 18417 3417 18429 3420
rect 18463 3417 18475 3451
rect 18417 3411 18475 3417
rect 3970 3380 3976 3392
rect 3931 3352 3976 3380
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 4525 3383 4583 3389
rect 4525 3349 4537 3383
rect 4571 3380 4583 3383
rect 4614 3380 4620 3392
rect 4571 3352 4620 3380
rect 4571 3349 4583 3352
rect 4525 3343 4583 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5074 3380 5080 3392
rect 5035 3352 5080 3380
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5626 3380 5632 3392
rect 5587 3352 5632 3380
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 6733 3383 6791 3389
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 6914 3380 6920 3392
rect 6779 3352 6920 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 12805 3383 12863 3389
rect 12805 3349 12817 3383
rect 12851 3380 12863 3383
rect 12894 3380 12900 3392
rect 12851 3352 12900 3380
rect 12851 3349 12863 3352
rect 12805 3343 12863 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 13446 3380 13452 3392
rect 13403 3352 13452 3380
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 13446 3340 13452 3352
rect 13504 3340 13510 3392
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 15930 3380 15936 3392
rect 14691 3352 15936 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16022 3340 16028 3392
rect 16080 3380 16086 3392
rect 18524 3380 18552 3479
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20165 3519 20223 3525
rect 20165 3516 20177 3519
rect 19484 3488 20177 3516
rect 19484 3476 19490 3488
rect 20165 3485 20177 3488
rect 20211 3485 20223 3519
rect 20530 3516 20536 3528
rect 20491 3488 20536 3516
rect 20165 3479 20223 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 21726 3516 21732 3528
rect 21687 3488 21732 3516
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 20254 3448 20260 3460
rect 20215 3420 20260 3448
rect 20254 3408 20260 3420
rect 20312 3408 20318 3460
rect 20346 3408 20352 3460
rect 20404 3448 20410 3460
rect 20404 3420 20449 3448
rect 20404 3408 20410 3420
rect 16080 3352 18552 3380
rect 20548 3380 20576 3476
rect 21818 3448 21824 3460
rect 21779 3420 21824 3448
rect 21818 3408 21824 3420
rect 21876 3408 21882 3460
rect 21928 3457 21956 3556
rect 22112 3556 22376 3584
rect 22112 3525 22140 3556
rect 22370 3544 22376 3556
rect 22428 3584 22434 3596
rect 22922 3584 22928 3596
rect 22428 3556 22928 3584
rect 22428 3544 22434 3556
rect 22922 3544 22928 3556
rect 22980 3584 22986 3596
rect 22980 3556 23152 3584
rect 22980 3544 22986 3556
rect 22077 3519 22140 3525
rect 22077 3485 22089 3519
rect 22123 3488 22140 3519
rect 22738 3516 22744 3528
rect 22699 3488 22744 3516
rect 22123 3485 22135 3488
rect 22077 3479 22135 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 23124 3525 23152 3556
rect 24210 3544 24216 3596
rect 24268 3584 24274 3596
rect 25409 3587 25467 3593
rect 25409 3584 25421 3587
rect 24268 3556 25421 3584
rect 24268 3544 24274 3556
rect 25409 3553 25421 3556
rect 25455 3553 25467 3587
rect 25409 3547 25467 3553
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23109 3519 23167 3525
rect 23109 3485 23121 3519
rect 23155 3516 23167 3519
rect 23290 3516 23296 3528
rect 23155 3488 23296 3516
rect 23155 3485 23167 3488
rect 23109 3479 23167 3485
rect 21913 3451 21971 3457
rect 21913 3417 21925 3451
rect 21959 3417 21971 3451
rect 21913 3411 21971 3417
rect 22554 3408 22560 3460
rect 22612 3448 22618 3460
rect 22848 3448 22876 3479
rect 23290 3476 23296 3488
rect 23348 3516 23354 3528
rect 24397 3519 24455 3525
rect 24397 3516 24409 3519
rect 23348 3488 24409 3516
rect 23348 3476 23354 3488
rect 24397 3485 24409 3488
rect 24443 3485 24455 3519
rect 24762 3516 24768 3528
rect 24723 3488 24768 3516
rect 24397 3479 24455 3485
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 36538 3476 36544 3528
rect 36596 3516 36602 3528
rect 36817 3519 36875 3525
rect 36817 3516 36829 3519
rect 36596 3488 36829 3516
rect 36596 3476 36602 3488
rect 36817 3485 36829 3488
rect 36863 3516 36875 3519
rect 37277 3519 37335 3525
rect 37277 3516 37289 3519
rect 36863 3488 37289 3516
rect 36863 3485 36875 3488
rect 36817 3479 36875 3485
rect 37277 3485 37289 3488
rect 37323 3485 37335 3519
rect 37277 3479 37335 3485
rect 22612 3420 22876 3448
rect 22612 3408 22618 3420
rect 22370 3380 22376 3392
rect 20548 3352 22376 3380
rect 16080 3340 16086 3352
rect 22370 3340 22376 3352
rect 22428 3340 22434 3392
rect 22848 3380 22876 3420
rect 22925 3451 22983 3457
rect 22925 3417 22937 3451
rect 22971 3448 22983 3451
rect 24302 3448 24308 3460
rect 22971 3420 24308 3448
rect 22971 3417 22983 3420
rect 22925 3411 22983 3417
rect 24302 3408 24308 3420
rect 24360 3408 24366 3460
rect 24578 3448 24584 3460
rect 24539 3420 24584 3448
rect 24578 3408 24584 3420
rect 24636 3408 24642 3460
rect 24673 3451 24731 3457
rect 24673 3417 24685 3451
rect 24719 3417 24731 3451
rect 24673 3411 24731 3417
rect 23106 3380 23112 3392
rect 22848 3352 23112 3380
rect 23106 3340 23112 3352
rect 23164 3380 23170 3392
rect 24688 3380 24716 3411
rect 24854 3408 24860 3460
rect 24912 3448 24918 3460
rect 25961 3451 26019 3457
rect 25961 3448 25973 3451
rect 24912 3420 25973 3448
rect 24912 3408 24918 3420
rect 25961 3417 25973 3420
rect 26007 3417 26019 3451
rect 25961 3411 26019 3417
rect 26050 3408 26056 3460
rect 26108 3448 26114 3460
rect 31202 3448 31208 3460
rect 26108 3420 31208 3448
rect 26108 3408 26114 3420
rect 31202 3408 31208 3420
rect 31260 3408 31266 3460
rect 23164 3352 24716 3380
rect 23164 3340 23170 3352
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28169 3383 28227 3389
rect 28169 3380 28181 3383
rect 27948 3352 28181 3380
rect 27948 3340 27954 3352
rect 28169 3349 28181 3352
rect 28215 3349 28227 3383
rect 28169 3343 28227 3349
rect 28534 3340 28540 3392
rect 28592 3380 28598 3392
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 28592 3352 28733 3380
rect 28592 3340 28598 3352
rect 28721 3349 28733 3352
rect 28767 3349 28779 3383
rect 29546 3380 29552 3392
rect 29507 3352 29552 3380
rect 28721 3343 28779 3349
rect 29546 3340 29552 3352
rect 29604 3340 29610 3392
rect 30469 3383 30527 3389
rect 30469 3349 30481 3383
rect 30515 3380 30527 3383
rect 30742 3380 30748 3392
rect 30515 3352 30748 3380
rect 30515 3349 30527 3352
rect 30469 3343 30527 3349
rect 30742 3340 30748 3352
rect 30800 3340 30806 3392
rect 31113 3383 31171 3389
rect 31113 3349 31125 3383
rect 31159 3380 31171 3383
rect 31386 3380 31392 3392
rect 31159 3352 31392 3380
rect 31159 3349 31171 3352
rect 31113 3343 31171 3349
rect 31386 3340 31392 3352
rect 31444 3340 31450 3392
rect 33226 3380 33232 3392
rect 33187 3352 33232 3380
rect 33226 3340 33232 3352
rect 33284 3340 33290 3392
rect 33686 3380 33692 3392
rect 33647 3352 33692 3380
rect 33686 3340 33692 3352
rect 33744 3340 33750 3392
rect 34698 3380 34704 3392
rect 34659 3352 34704 3380
rect 34698 3340 34704 3352
rect 34756 3340 34762 3392
rect 35437 3383 35495 3389
rect 35437 3349 35449 3383
rect 35483 3380 35495 3383
rect 35802 3380 35808 3392
rect 35483 3352 35808 3380
rect 35483 3349 35495 3352
rect 35437 3343 35495 3349
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 35986 3380 35992 3392
rect 35947 3352 35992 3380
rect 35986 3340 35992 3352
rect 36044 3340 36050 3392
rect 38010 3380 38016 3392
rect 37971 3352 38016 3380
rect 38010 3340 38016 3352
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 3145 3179 3203 3185
rect 3145 3176 3157 3179
rect 2924 3148 3157 3176
rect 2924 3136 2930 3148
rect 3145 3145 3157 3148
rect 3191 3145 3203 3179
rect 3145 3139 3203 3145
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3145 4767 3179
rect 4709 3139 4767 3145
rect 7009 3179 7067 3185
rect 7009 3145 7021 3179
rect 7055 3176 7067 3179
rect 7282 3176 7288 3188
rect 7055 3148 7288 3176
rect 7055 3145 7067 3148
rect 7009 3139 7067 3145
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3040 2559 3043
rect 2866 3040 2872 3052
rect 2547 3012 2872 3040
rect 2547 3009 2559 3012
rect 2501 3003 2559 3009
rect 2866 3000 2872 3012
rect 2924 3040 2930 3052
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2924 3012 3065 3040
rect 2924 3000 2930 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 3970 3040 3976 3052
rect 3927 3012 3976 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4614 3040 4620 3052
rect 4571 3012 4620 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4724 2972 4752 3139
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 10502 3136 10508 3188
rect 10560 3176 10566 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 10560 3148 10609 3176
rect 10560 3136 10566 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 13630 3176 13636 3188
rect 13591 3148 13636 3176
rect 10597 3139 10655 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 14369 3179 14427 3185
rect 14369 3145 14381 3179
rect 14415 3145 14427 3179
rect 15194 3176 15200 3188
rect 15155 3148 15200 3176
rect 14369 3139 14427 3145
rect 11606 3108 11612 3120
rect 8312 3080 11612 3108
rect 5074 3000 5080 3052
rect 5132 3040 5138 3052
rect 5169 3043 5227 3049
rect 5169 3040 5181 3043
rect 5132 3012 5181 3040
rect 5132 3000 5138 3012
rect 5169 3009 5181 3012
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 8312 2972 8340 3080
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 12989 3111 13047 3117
rect 12989 3077 13001 3111
rect 13035 3108 13047 3111
rect 14384 3108 14412 3139
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16117 3179 16175 3185
rect 16117 3145 16129 3179
rect 16163 3176 16175 3179
rect 16390 3176 16396 3188
rect 16163 3148 16396 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 16390 3136 16396 3148
rect 16448 3136 16454 3188
rect 16853 3179 16911 3185
rect 16853 3145 16865 3179
rect 16899 3176 16911 3179
rect 16942 3176 16948 3188
rect 16899 3148 16948 3176
rect 16899 3145 16911 3148
rect 16853 3139 16911 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17678 3176 17684 3188
rect 17368 3148 17684 3176
rect 17368 3136 17374 3148
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 17773 3179 17831 3185
rect 17773 3145 17785 3179
rect 17819 3176 17831 3179
rect 17862 3176 17868 3188
rect 17819 3148 17868 3176
rect 17819 3145 17831 3148
rect 17773 3139 17831 3145
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18506 3176 18512 3188
rect 18279 3148 18512 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 19518 3176 19524 3188
rect 18616 3148 19524 3176
rect 15838 3108 15844 3120
rect 13035 3080 14228 3108
rect 14384 3080 15844 3108
rect 13035 3077 13047 3080
rect 12989 3071 13047 3077
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 8444 3012 8493 3040
rect 8444 3000 8450 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 9490 3000 9496 3052
rect 9548 3040 9554 3052
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 9548 3012 9597 3040
rect 9548 3000 9554 3012
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 10594 3040 10600 3052
rect 10555 3012 10600 3040
rect 9585 3003 9643 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 11238 3040 11244 3052
rect 10827 3012 11244 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 11238 3000 11244 3012
rect 11296 3000 11302 3052
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 11756 3012 11805 3040
rect 11756 3000 11762 3012
rect 11793 3009 11805 3012
rect 11839 3009 11851 3043
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 11793 3003 11851 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 14200 3049 14228 3080
rect 15838 3068 15844 3080
rect 15896 3068 15902 3120
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 17405 3111 17463 3117
rect 17405 3108 17417 3111
rect 16356 3080 17417 3108
rect 16356 3068 16362 3080
rect 17405 3077 17417 3080
rect 17451 3077 17463 3111
rect 17405 3071 17463 3077
rect 18046 3068 18052 3120
rect 18104 3108 18110 3120
rect 18616 3108 18644 3148
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 19797 3179 19855 3185
rect 19797 3145 19809 3179
rect 19843 3176 19855 3179
rect 20070 3176 20076 3188
rect 19843 3148 20076 3176
rect 19843 3145 19855 3148
rect 19797 3139 19855 3145
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 21634 3136 21640 3188
rect 21692 3176 21698 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 21692 3148 21833 3176
rect 21692 3136 21698 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 22833 3179 22891 3185
rect 22833 3176 22845 3179
rect 22244 3148 22845 3176
rect 22244 3136 22250 3148
rect 22833 3145 22845 3148
rect 22879 3145 22891 3179
rect 24394 3176 24400 3188
rect 24355 3148 24400 3176
rect 22833 3139 22891 3145
rect 24394 3136 24400 3148
rect 24452 3136 24458 3188
rect 28353 3179 28411 3185
rect 28353 3176 28365 3179
rect 25056 3148 28365 3176
rect 18966 3108 18972 3120
rect 18104 3080 18644 3108
rect 18708 3080 18972 3108
rect 18104 3068 18110 3080
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3040 14243 3043
rect 14458 3040 14464 3052
rect 14231 3012 14464 3040
rect 14231 3009 14243 3012
rect 14185 3003 14243 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 11330 2972 11336 2984
rect 4724 2944 8340 2972
rect 8588 2944 11336 2972
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 5353 2907 5411 2913
rect 4111 2876 5304 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 5276 2836 5304 2876
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 8588 2904 8616 2944
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 14844 2972 14872 3003
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 15930 3040 15936 3052
rect 15068 3012 15113 3040
rect 15891 3012 15936 3040
rect 15068 3000 15074 3012
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 17218 3000 17224 3052
rect 17276 3040 17282 3052
rect 17313 3043 17371 3049
rect 17313 3040 17325 3043
rect 17276 3012 17325 3040
rect 17276 3000 17282 3012
rect 17313 3009 17325 3012
rect 17359 3009 17371 3043
rect 17586 3040 17592 3052
rect 17547 3012 17592 3040
rect 17313 3003 17371 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 18524 3049 18552 3080
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 18380 3012 18429 3040
rect 18380 3000 18386 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 18601 3043 18659 3049
rect 18601 3009 18613 3043
rect 18647 3040 18659 3043
rect 18708 3040 18736 3080
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 19429 3111 19487 3117
rect 19429 3077 19441 3111
rect 19475 3108 19487 3111
rect 22554 3108 22560 3120
rect 19475 3080 22560 3108
rect 19475 3077 19487 3080
rect 19429 3071 19487 3077
rect 22554 3068 22560 3080
rect 22612 3068 22618 3120
rect 23106 3108 23112 3120
rect 23067 3080 23112 3108
rect 23106 3068 23112 3080
rect 23164 3108 23170 3120
rect 24029 3111 24087 3117
rect 23164 3080 23980 3108
rect 23164 3068 23170 3080
rect 18647 3012 18736 3040
rect 18785 3043 18843 3049
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 18785 3009 18797 3043
rect 18831 3040 18843 3043
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18831 3012 19257 3040
rect 18831 3009 18843 3012
rect 18785 3003 18843 3009
rect 19245 3009 19257 3012
rect 19291 3040 19303 3043
rect 19334 3040 19340 3052
rect 19291 3012 19340 3040
rect 19291 3009 19303 3012
rect 19245 3003 19303 3009
rect 16758 2972 16764 2984
rect 12584 2944 16764 2972
rect 12584 2932 12590 2944
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 17770 2932 17776 2984
rect 17828 2972 17834 2984
rect 18800 2972 18828 3003
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19518 3040 19524 3052
rect 19479 3012 19524 3040
rect 19518 3000 19524 3012
rect 19576 3000 19582 3052
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3040 19671 3043
rect 19978 3040 19984 3052
rect 19659 3012 19984 3040
rect 19659 3009 19671 3012
rect 19613 3003 19671 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 20533 3043 20591 3049
rect 20533 3040 20545 3043
rect 20496 3012 20545 3040
rect 20496 3000 20502 3012
rect 20533 3009 20545 3012
rect 20579 3040 20591 3043
rect 20993 3043 21051 3049
rect 20993 3040 21005 3043
rect 20579 3012 21005 3040
rect 20579 3009 20591 3012
rect 20533 3003 20591 3009
rect 20993 3009 21005 3012
rect 21039 3009 21051 3043
rect 22002 3040 22008 3052
rect 21963 3012 22008 3040
rect 20993 3003 21051 3009
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3009 22155 3043
rect 22097 3003 22155 3009
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22370 3040 22376 3052
rect 22331 3012 22376 3040
rect 22189 3003 22247 3009
rect 17828 2944 18828 2972
rect 19536 2972 19564 3000
rect 20254 2972 20260 2984
rect 19536 2944 20260 2972
rect 17828 2932 17834 2944
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 21818 2972 21824 2984
rect 20772 2944 21824 2972
rect 20772 2932 20778 2944
rect 21818 2932 21824 2944
rect 21876 2972 21882 2984
rect 22112 2972 22140 3003
rect 21876 2944 22140 2972
rect 22204 2972 22232 3003
rect 22370 3000 22376 3012
rect 22428 3000 22434 3052
rect 23014 3049 23020 3052
rect 22993 3043 23020 3049
rect 22993 3009 23005 3043
rect 22993 3003 23020 3009
rect 23014 3000 23020 3003
rect 23072 3000 23078 3052
rect 23201 3043 23259 3049
rect 23201 3040 23213 3043
rect 23124 3012 23213 3040
rect 23124 2984 23152 3012
rect 23201 3009 23213 3012
rect 23247 3009 23259 3043
rect 23201 3003 23259 3009
rect 23290 3000 23296 3052
rect 23348 3040 23354 3052
rect 23385 3043 23443 3049
rect 23385 3040 23397 3043
rect 23348 3012 23397 3040
rect 23348 3000 23354 3012
rect 23385 3009 23397 3012
rect 23431 3040 23443 3043
rect 23845 3043 23903 3049
rect 23845 3040 23857 3043
rect 23431 3012 23857 3040
rect 23431 3009 23443 3012
rect 23385 3003 23443 3009
rect 23845 3009 23857 3012
rect 23891 3009 23903 3043
rect 23952 3040 23980 3080
rect 24029 3077 24041 3111
rect 24075 3108 24087 3111
rect 25056 3108 25084 3148
rect 28353 3145 28365 3148
rect 28399 3145 28411 3179
rect 28994 3176 29000 3188
rect 28955 3148 29000 3176
rect 28353 3139 28411 3145
rect 28994 3136 29000 3148
rect 29052 3136 29058 3188
rect 31202 3176 31208 3188
rect 31163 3148 31208 3176
rect 31202 3136 31208 3148
rect 31260 3136 31266 3188
rect 33318 3176 33324 3188
rect 33279 3148 33324 3176
rect 33318 3136 33324 3148
rect 33376 3136 33382 3188
rect 34425 3179 34483 3185
rect 34425 3145 34437 3179
rect 34471 3145 34483 3179
rect 34425 3139 34483 3145
rect 26329 3111 26387 3117
rect 26329 3108 26341 3111
rect 24075 3080 25084 3108
rect 25148 3080 26341 3108
rect 24075 3077 24087 3080
rect 24029 3071 24087 3077
rect 25148 3052 25176 3080
rect 26329 3077 26341 3080
rect 26375 3077 26387 3111
rect 26329 3071 26387 3077
rect 27522 3068 27528 3120
rect 27580 3108 27586 3120
rect 34440 3108 34468 3139
rect 34514 3136 34520 3188
rect 34572 3176 34578 3188
rect 36081 3179 36139 3185
rect 36081 3176 36093 3179
rect 34572 3148 36093 3176
rect 34572 3136 34578 3148
rect 36081 3145 36093 3148
rect 36127 3145 36139 3179
rect 36081 3139 36139 3145
rect 27580 3080 34468 3108
rect 27580 3068 27586 3080
rect 24121 3043 24179 3049
rect 24121 3040 24133 3043
rect 23952 3012 24133 3040
rect 23845 3003 23903 3009
rect 24121 3009 24133 3012
rect 24167 3009 24179 3043
rect 24121 3003 24179 3009
rect 24210 3000 24216 3052
rect 24268 3040 24274 3052
rect 25130 3040 25136 3052
rect 24268 3012 24313 3040
rect 25091 3012 25136 3040
rect 24268 3000 24274 3012
rect 25130 3000 25136 3012
rect 25188 3000 25194 3052
rect 25590 3040 25596 3052
rect 25551 3012 25596 3040
rect 25590 3000 25596 3012
rect 25648 3000 25654 3052
rect 26973 3043 27031 3049
rect 26973 3009 26985 3043
rect 27019 3040 27031 3043
rect 27062 3040 27068 3052
rect 27019 3012 27068 3040
rect 27019 3009 27031 3012
rect 26973 3003 27031 3009
rect 27062 3000 27068 3012
rect 27120 3000 27126 3052
rect 27154 3000 27160 3052
rect 27212 3040 27218 3052
rect 27890 3040 27896 3052
rect 27212 3012 27896 3040
rect 27212 3000 27218 3012
rect 27890 3000 27896 3012
rect 27948 3000 27954 3052
rect 28258 3000 28264 3052
rect 28316 3040 28322 3052
rect 28534 3040 28540 3052
rect 28316 3012 28540 3040
rect 28316 3000 28322 3012
rect 28534 3000 28540 3012
rect 28592 3000 28598 3052
rect 30466 3000 30472 3052
rect 30524 3040 30530 3052
rect 30742 3040 30748 3052
rect 30524 3012 30748 3040
rect 30524 3000 30530 3012
rect 30742 3000 30748 3012
rect 30800 3000 30806 3052
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 31386 3040 31392 3052
rect 31076 3012 31392 3040
rect 31076 3000 31082 3012
rect 31386 3000 31392 3012
rect 31444 3000 31450 3052
rect 33226 3000 33232 3052
rect 33284 3040 33290 3052
rect 33505 3043 33563 3049
rect 33505 3040 33517 3043
rect 33284 3012 33517 3040
rect 33284 3000 33290 3012
rect 33505 3009 33517 3012
rect 33551 3009 33563 3043
rect 33505 3003 33563 3009
rect 34330 3000 34336 3052
rect 34388 3040 34394 3052
rect 34609 3043 34667 3049
rect 34609 3040 34621 3043
rect 34388 3012 34621 3040
rect 34388 3000 34394 3012
rect 34609 3009 34621 3012
rect 34655 3040 34667 3043
rect 35069 3043 35127 3049
rect 35069 3040 35081 3043
rect 34655 3012 35081 3040
rect 34655 3009 34667 3012
rect 34609 3003 34667 3009
rect 35069 3009 35081 3012
rect 35115 3009 35127 3043
rect 35069 3003 35127 3009
rect 35986 3000 35992 3052
rect 36044 3040 36050 3052
rect 36265 3043 36323 3049
rect 36265 3040 36277 3043
rect 36044 3012 36277 3040
rect 36044 3000 36050 3012
rect 36265 3009 36277 3012
rect 36311 3009 36323 3043
rect 36265 3003 36323 3009
rect 37090 3000 37096 3052
rect 37148 3040 37154 3052
rect 37553 3043 37611 3049
rect 37553 3040 37565 3043
rect 37148 3012 37565 3040
rect 37148 3000 37154 3012
rect 37553 3009 37565 3012
rect 37599 3040 37611 3043
rect 38013 3043 38071 3049
rect 38013 3040 38025 3043
rect 37599 3012 38025 3040
rect 37599 3009 37611 3012
rect 37553 3003 37611 3009
rect 38013 3009 38025 3012
rect 38059 3009 38071 3043
rect 38013 3003 38071 3009
rect 22204 2944 22876 2972
rect 21876 2932 21882 2944
rect 5399 2876 8616 2904
rect 8665 2907 8723 2913
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 8665 2873 8677 2907
rect 8711 2904 8723 2907
rect 11882 2904 11888 2916
rect 8711 2876 11888 2904
rect 8711 2873 8723 2876
rect 8665 2867 8723 2873
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 11977 2907 12035 2913
rect 11977 2873 11989 2907
rect 12023 2904 12035 2907
rect 16022 2904 16028 2916
rect 12023 2876 16028 2904
rect 12023 2873 12035 2876
rect 11977 2867 12035 2873
rect 7374 2836 7380 2848
rect 5276 2808 7380 2836
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2836 8079 2839
rect 9674 2836 9680 2848
rect 8067 2808 9680 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9769 2839 9827 2845
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 13538 2836 13544 2848
rect 9815 2808 13544 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 14826 2836 14832 2848
rect 13780 2808 14832 2836
rect 13780 2796 13786 2808
rect 14826 2796 14832 2808
rect 14884 2796 14890 2848
rect 14936 2845 14964 2876
rect 16022 2864 16028 2876
rect 16080 2864 16086 2916
rect 16114 2864 16120 2916
rect 16172 2904 16178 2916
rect 16172 2876 19012 2904
rect 16172 2864 16178 2876
rect 14921 2839 14979 2845
rect 14921 2805 14933 2839
rect 14967 2805 14979 2839
rect 14921 2799 14979 2805
rect 15010 2796 15016 2848
rect 15068 2836 15074 2848
rect 18874 2836 18880 2848
rect 15068 2808 18880 2836
rect 15068 2796 15074 2808
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 18984 2836 19012 2876
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 20349 2907 20407 2913
rect 20349 2904 20361 2907
rect 19484 2876 20361 2904
rect 19484 2864 19490 2876
rect 20349 2873 20361 2876
rect 20395 2873 20407 2907
rect 20349 2867 20407 2873
rect 22278 2864 22284 2916
rect 22336 2904 22342 2916
rect 22848 2904 22876 2944
rect 23106 2932 23112 2984
rect 23164 2932 23170 2984
rect 23216 2944 30604 2972
rect 23216 2904 23244 2944
rect 22336 2876 22692 2904
rect 22848 2876 23244 2904
rect 22336 2864 22342 2876
rect 21450 2836 21456 2848
rect 18984 2808 21456 2836
rect 21450 2796 21456 2808
rect 21508 2796 21514 2848
rect 22186 2796 22192 2848
rect 22244 2836 22250 2848
rect 22554 2836 22560 2848
rect 22244 2808 22560 2836
rect 22244 2796 22250 2808
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 22664 2836 22692 2876
rect 23290 2864 23296 2916
rect 23348 2904 23354 2916
rect 25222 2904 25228 2916
rect 23348 2876 25228 2904
rect 23348 2864 23354 2876
rect 25222 2864 25228 2876
rect 25280 2864 25286 2916
rect 26050 2864 26056 2916
rect 26108 2904 26114 2916
rect 27157 2907 27215 2913
rect 27157 2904 27169 2907
rect 26108 2876 27169 2904
rect 26108 2864 26114 2876
rect 27157 2873 27169 2876
rect 27203 2873 27215 2907
rect 27157 2867 27215 2873
rect 28626 2864 28632 2916
rect 28684 2904 28690 2916
rect 30576 2913 30604 2944
rect 29549 2907 29607 2913
rect 29549 2904 29561 2907
rect 28684 2876 29561 2904
rect 28684 2864 28690 2876
rect 29549 2873 29561 2876
rect 29595 2873 29607 2907
rect 29549 2867 29607 2873
rect 30561 2907 30619 2913
rect 30561 2873 30573 2907
rect 30607 2873 30619 2907
rect 30561 2867 30619 2873
rect 33134 2864 33140 2916
rect 33192 2904 33198 2916
rect 37369 2907 37427 2913
rect 37369 2904 37381 2907
rect 33192 2876 37381 2904
rect 33192 2864 33198 2876
rect 37369 2873 37381 2876
rect 37415 2873 37427 2907
rect 37369 2867 37427 2873
rect 22830 2836 22836 2848
rect 22664 2808 22836 2836
rect 22830 2796 22836 2808
rect 22888 2796 22894 2848
rect 23842 2796 23848 2848
rect 23900 2836 23906 2848
rect 24949 2839 25007 2845
rect 24949 2836 24961 2839
rect 23900 2808 24961 2836
rect 23900 2796 23906 2808
rect 24949 2805 24961 2808
rect 24995 2805 25007 2839
rect 24949 2799 25007 2805
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 25777 2839 25835 2845
rect 25777 2836 25789 2839
rect 25096 2808 25789 2836
rect 25096 2796 25102 2808
rect 25777 2805 25789 2808
rect 25823 2805 25835 2839
rect 25777 2799 25835 2805
rect 26326 2796 26332 2848
rect 26384 2836 26390 2848
rect 27709 2839 27767 2845
rect 27709 2836 27721 2839
rect 26384 2808 27721 2836
rect 26384 2796 26390 2808
rect 27709 2805 27721 2808
rect 27755 2805 27767 2839
rect 27709 2799 27767 2805
rect 31478 2796 31484 2848
rect 31536 2836 31542 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31536 2808 32137 2836
rect 31536 2796 31542 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32674 2836 32680 2848
rect 32635 2808 32680 2836
rect 32125 2799 32183 2805
rect 32674 2796 32680 2808
rect 32732 2796 32738 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 9677 2635 9735 2641
rect 9677 2601 9689 2635
rect 9723 2632 9735 2635
rect 19429 2635 19487 2641
rect 9723 2604 16574 2632
rect 9723 2601 9735 2604
rect 9677 2595 9735 2601
rect 4706 2564 4712 2576
rect 3988 2536 4712 2564
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2496 2743 2499
rect 3988 2496 4016 2536
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 5810 2564 5816 2576
rect 5771 2536 5816 2564
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2533 10379 2567
rect 10321 2527 10379 2533
rect 12253 2567 12311 2573
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 13722 2564 13728 2576
rect 12299 2536 13728 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 7006 2496 7012 2508
rect 2731 2468 4016 2496
rect 4080 2468 7012 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2314 2428 2320 2440
rect 1995 2400 2320 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2314 2388 2320 2400
rect 2372 2428 2378 2440
rect 4080 2437 4108 2468
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 10042 2496 10048 2508
rect 8036 2468 10048 2496
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2372 2400 2421 2428
rect 2372 2388 2378 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5442 2428 5448 2440
rect 5031 2400 5448 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 5626 2428 5632 2440
rect 5539 2400 5632 2428
rect 5626 2388 5632 2400
rect 5684 2428 5690 2440
rect 6178 2428 6184 2440
rect 5684 2400 6184 2428
rect 5684 2388 5690 2400
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7282 2428 7288 2440
rect 6972 2400 7288 2428
rect 6972 2388 6978 2400
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 7834 2428 7840 2440
rect 7607 2400 7840 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 6457 2363 6515 2369
rect 6457 2329 6469 2363
rect 6503 2360 6515 2363
rect 8036 2360 8064 2468
rect 8202 2428 8208 2440
rect 8115 2400 8208 2428
rect 8202 2388 8208 2400
rect 8260 2428 8266 2440
rect 8938 2428 8944 2440
rect 8260 2400 8944 2428
rect 8260 2388 8266 2400
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9508 2437 9536 2468
rect 10042 2456 10048 2468
rect 10100 2456 10106 2508
rect 10336 2496 10364 2527
rect 13722 2524 13728 2536
rect 13780 2524 13786 2576
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 15194 2564 15200 2576
rect 14783 2536 15200 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 15381 2567 15439 2573
rect 15381 2533 15393 2567
rect 15427 2564 15439 2567
rect 16298 2564 16304 2576
rect 15427 2536 16304 2564
rect 15427 2533 15439 2536
rect 15381 2527 15439 2533
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 10336 2468 15332 2496
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9732 2400 10149 2428
rect 9732 2388 9738 2400
rect 10137 2397 10149 2400
rect 10183 2428 10195 2431
rect 10594 2428 10600 2440
rect 10183 2400 10600 2428
rect 10183 2397 10195 2400
rect 10137 2391 10195 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10781 2431 10839 2437
rect 10781 2397 10793 2431
rect 10827 2428 10839 2431
rect 10962 2428 10968 2440
rect 10827 2400 10968 2428
rect 10827 2397 10839 2400
rect 10781 2391 10839 2397
rect 6503 2332 8064 2360
rect 9033 2363 9091 2369
rect 6503 2329 6515 2332
rect 6457 2323 6515 2329
rect 9033 2329 9045 2363
rect 9079 2360 9091 2363
rect 10796 2360 10824 2391
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12250 2428 12256 2440
rect 12115 2400 12256 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 12802 2428 12808 2440
rect 12759 2400 12808 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 9079 2332 10824 2360
rect 11609 2363 11667 2369
rect 9079 2329 9091 2332
rect 9033 2323 9091 2329
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 12728 2360 12756 2391
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 12952 2400 13369 2428
rect 12952 2388 12958 2400
rect 13357 2397 13369 2400
rect 13403 2428 13415 2431
rect 13722 2428 13728 2440
rect 13403 2400 13728 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 14148 2400 14565 2428
rect 14148 2388 14154 2400
rect 14553 2397 14565 2400
rect 14599 2428 14611 2431
rect 15010 2428 15016 2440
rect 14599 2400 15016 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 15304 2428 15332 2468
rect 15746 2456 15752 2508
rect 15804 2496 15810 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15804 2468 15853 2496
rect 15804 2456 15810 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 16546 2496 16574 2604
rect 19429 2601 19441 2635
rect 19475 2632 19487 2635
rect 20254 2632 20260 2644
rect 19475 2604 20260 2632
rect 19475 2601 19487 2604
rect 19429 2595 19487 2601
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 25222 2632 25228 2644
rect 25183 2604 25228 2632
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 28445 2635 28503 2641
rect 28445 2632 28457 2635
rect 25332 2604 28457 2632
rect 20622 2524 20628 2576
rect 20680 2524 20686 2576
rect 21634 2524 21640 2576
rect 21692 2564 21698 2576
rect 22649 2567 22707 2573
rect 22649 2564 22661 2567
rect 21692 2536 22661 2564
rect 21692 2524 21698 2536
rect 22649 2533 22661 2536
rect 22695 2533 22707 2567
rect 22649 2527 22707 2533
rect 18322 2496 18328 2508
rect 16546 2468 18328 2496
rect 15841 2459 15899 2465
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 20640 2496 20668 2524
rect 20180 2468 20668 2496
rect 16850 2428 16856 2440
rect 15304 2400 16856 2428
rect 15197 2391 15255 2397
rect 14918 2360 14924 2372
rect 11655 2332 12756 2360
rect 12912 2332 14924 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 3881 2295 3939 2301
rect 3881 2292 3893 2295
rect 3476 2264 3893 2292
rect 3476 2252 3482 2264
rect 3881 2261 3893 2264
rect 3927 2261 3939 2295
rect 5166 2292 5172 2304
rect 5127 2264 5172 2292
rect 3881 2255 3939 2261
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7742 2292 7748 2304
rect 7703 2264 7748 2292
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 8389 2295 8447 2301
rect 8389 2261 8401 2295
rect 8435 2292 8447 2295
rect 9582 2292 9588 2304
rect 8435 2264 9588 2292
rect 8435 2261 8447 2264
rect 8389 2255 8447 2261
rect 9582 2252 9588 2264
rect 9640 2252 9646 2304
rect 10965 2295 11023 2301
rect 10965 2261 10977 2295
rect 11011 2292 11023 2295
rect 12342 2292 12348 2304
rect 11011 2264 12348 2292
rect 11011 2261 11023 2264
rect 10965 2255 11023 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 12912 2301 12940 2332
rect 14918 2320 14924 2332
rect 14976 2320 14982 2372
rect 15212 2360 15240 2391
rect 16850 2388 16856 2400
rect 16908 2388 16914 2440
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17678 2428 17684 2440
rect 17000 2400 17045 2428
rect 17639 2400 17684 2428
rect 17000 2388 17006 2400
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 18230 2388 18236 2440
rect 18288 2428 18294 2440
rect 20180 2437 20208 2468
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22152 2468 23704 2496
rect 22152 2456 22158 2468
rect 18417 2431 18475 2437
rect 18417 2428 18429 2431
rect 18288 2400 18429 2428
rect 18288 2388 18294 2400
rect 18417 2397 18429 2400
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 20165 2431 20223 2437
rect 20165 2397 20177 2431
rect 20211 2397 20223 2431
rect 20165 2391 20223 2397
rect 20254 2388 20260 2440
rect 20312 2428 20318 2440
rect 20625 2431 20683 2437
rect 20625 2428 20637 2431
rect 20312 2400 20637 2428
rect 20312 2388 20318 2400
rect 20625 2397 20637 2400
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 20898 2388 20904 2440
rect 20956 2428 20962 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 20956 2400 21833 2428
rect 20956 2388 20962 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 22278 2388 22284 2440
rect 22336 2428 22342 2440
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22336 2400 22845 2428
rect 22336 2388 22342 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22833 2391 22891 2397
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23532 2400 23581 2428
rect 23532 2388 23538 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23676 2428 23704 2468
rect 24578 2456 24584 2508
rect 24636 2496 24642 2508
rect 25332 2496 25360 2604
rect 28445 2601 28457 2604
rect 28491 2601 28503 2635
rect 35345 2635 35403 2641
rect 35345 2632 35357 2635
rect 28445 2595 28503 2601
rect 28552 2604 35357 2632
rect 25958 2564 25964 2576
rect 25919 2536 25964 2564
rect 25958 2524 25964 2536
rect 26016 2524 26022 2576
rect 26602 2524 26608 2576
rect 26660 2564 26666 2576
rect 27801 2567 27859 2573
rect 27801 2564 27813 2567
rect 26660 2536 27813 2564
rect 26660 2524 26666 2536
rect 27801 2533 27813 2536
rect 27847 2533 27859 2567
rect 28552 2564 28580 2604
rect 35345 2601 35357 2604
rect 35391 2601 35403 2635
rect 35345 2595 35403 2601
rect 27801 2527 27859 2533
rect 27908 2536 28580 2564
rect 26510 2496 26516 2508
rect 24636 2468 25360 2496
rect 25424 2468 26516 2496
rect 24636 2456 24642 2468
rect 24673 2431 24731 2437
rect 23676 2400 24624 2428
rect 23569 2391 23627 2397
rect 15286 2360 15292 2372
rect 15199 2332 15292 2360
rect 15286 2320 15292 2332
rect 15344 2360 15350 2372
rect 15562 2360 15568 2372
rect 15344 2332 15568 2360
rect 15344 2320 15350 2332
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 16025 2363 16083 2369
rect 16025 2329 16037 2363
rect 16071 2360 16083 2363
rect 16574 2360 16580 2372
rect 16071 2332 16580 2360
rect 16071 2329 16083 2332
rect 16025 2323 16083 2329
rect 16574 2320 16580 2332
rect 16632 2360 16638 2372
rect 17218 2360 17224 2372
rect 16632 2332 17224 2360
rect 16632 2320 16638 2332
rect 17218 2320 17224 2332
rect 17276 2320 17282 2372
rect 22738 2320 22744 2372
rect 22796 2360 22802 2372
rect 22796 2332 24532 2360
rect 22796 2320 22802 2332
rect 12897 2295 12955 2301
rect 12897 2261 12909 2295
rect 12943 2261 12955 2295
rect 12897 2255 12955 2261
rect 13541 2295 13599 2301
rect 13541 2261 13553 2295
rect 13587 2292 13599 2295
rect 15102 2292 15108 2304
rect 13587 2264 15108 2292
rect 13587 2261 13599 2264
rect 13541 2255 13599 2261
rect 15102 2252 15108 2264
rect 15160 2252 15166 2304
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 16206 2292 16212 2304
rect 15252 2264 16212 2292
rect 15252 2252 15258 2264
rect 16206 2252 16212 2264
rect 16264 2252 16270 2304
rect 17129 2295 17187 2301
rect 17129 2261 17141 2295
rect 17175 2292 17187 2295
rect 17770 2292 17776 2304
rect 17175 2264 17776 2292
rect 17175 2261 17187 2264
rect 17129 2255 17187 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 17865 2295 17923 2301
rect 17865 2261 17877 2295
rect 17911 2292 17923 2295
rect 18322 2292 18328 2304
rect 17911 2264 18328 2292
rect 17911 2261 17923 2264
rect 17865 2255 17923 2261
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 18874 2292 18880 2304
rect 18647 2264 18880 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 18874 2252 18880 2264
rect 18932 2252 18938 2304
rect 19978 2292 19984 2304
rect 19939 2264 19984 2292
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 20530 2252 20536 2304
rect 20588 2292 20594 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20588 2264 20821 2292
rect 20588 2252 20594 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 20809 2255 20867 2261
rect 21082 2252 21088 2304
rect 21140 2292 21146 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21140 2264 22017 2292
rect 21140 2252 21146 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 24504 2301 24532 2332
rect 23385 2295 23443 2301
rect 23385 2292 23397 2295
rect 22244 2264 23397 2292
rect 22244 2252 22250 2264
rect 23385 2261 23397 2264
rect 23431 2261 23443 2295
rect 23385 2255 23443 2261
rect 24489 2295 24547 2301
rect 24489 2261 24501 2295
rect 24535 2261 24547 2295
rect 24596 2292 24624 2400
rect 24673 2397 24685 2431
rect 24719 2428 24731 2431
rect 24854 2428 24860 2440
rect 24719 2400 24860 2428
rect 24719 2397 24731 2400
rect 24673 2391 24731 2397
rect 24854 2388 24860 2400
rect 24912 2388 24918 2440
rect 25424 2437 25452 2468
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 27908 2496 27936 2536
rect 28810 2524 28816 2576
rect 28868 2564 28874 2576
rect 30837 2567 30895 2573
rect 30837 2564 30849 2567
rect 28868 2536 30849 2564
rect 28868 2524 28874 2536
rect 30837 2533 30849 2536
rect 30883 2533 30895 2567
rect 30837 2527 30895 2533
rect 26988 2468 27936 2496
rect 28000 2468 28764 2496
rect 25409 2431 25467 2437
rect 25409 2397 25421 2431
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2428 26203 2431
rect 26234 2428 26240 2440
rect 26191 2400 26240 2428
rect 26191 2397 26203 2400
rect 26145 2391 26203 2397
rect 26234 2388 26240 2400
rect 26292 2388 26298 2440
rect 25498 2320 25504 2372
rect 25556 2360 25562 2372
rect 26878 2360 26884 2372
rect 25556 2332 26884 2360
rect 25556 2320 25562 2332
rect 26878 2320 26884 2332
rect 26936 2320 26942 2372
rect 26988 2292 27016 2468
rect 27249 2431 27307 2437
rect 27249 2397 27261 2431
rect 27295 2428 27307 2431
rect 27614 2428 27620 2440
rect 27295 2400 27620 2428
rect 27295 2397 27307 2400
rect 27249 2391 27307 2397
rect 27614 2388 27620 2400
rect 27672 2388 27678 2440
rect 28000 2437 28028 2468
rect 27985 2431 28043 2437
rect 27985 2397 27997 2431
rect 28031 2397 28043 2431
rect 28626 2428 28632 2440
rect 28539 2400 28632 2428
rect 27985 2391 28043 2397
rect 28626 2388 28632 2400
rect 28684 2388 28690 2440
rect 27706 2320 27712 2372
rect 27764 2360 27770 2372
rect 28644 2360 28672 2388
rect 27764 2332 28672 2360
rect 28736 2360 28764 2468
rect 29914 2456 29920 2508
rect 29972 2496 29978 2508
rect 31478 2496 31484 2508
rect 29972 2468 31484 2496
rect 29972 2456 29978 2468
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29546 2428 29552 2440
rect 29052 2400 29552 2428
rect 29052 2388 29058 2400
rect 29546 2388 29552 2400
rect 29604 2428 29610 2440
rect 31036 2437 31064 2468
rect 31478 2456 31484 2468
rect 31536 2456 31542 2508
rect 37642 2456 37648 2508
rect 37700 2496 37706 2508
rect 38010 2496 38016 2508
rect 37700 2468 38016 2496
rect 37700 2456 37706 2468
rect 38010 2456 38016 2468
rect 38068 2496 38074 2508
rect 38105 2499 38163 2505
rect 38105 2496 38117 2499
rect 38068 2468 38117 2496
rect 38068 2456 38074 2468
rect 38105 2465 38117 2468
rect 38151 2465 38163 2499
rect 38105 2459 38163 2465
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29604 2400 29745 2428
rect 29604 2388 29610 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30377 2431 30435 2437
rect 30377 2397 30389 2431
rect 30423 2397 30435 2431
rect 30377 2391 30435 2397
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 29086 2360 29092 2372
rect 28736 2332 29092 2360
rect 27764 2320 27770 2332
rect 29086 2320 29092 2332
rect 29144 2320 29150 2372
rect 29362 2320 29368 2372
rect 29420 2360 29426 2372
rect 30392 2360 30420 2391
rect 31754 2388 31760 2440
rect 31812 2428 31818 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 31812 2400 32321 2428
rect 31812 2388 31818 2400
rect 32309 2397 32321 2400
rect 32355 2428 32367 2431
rect 32674 2428 32680 2440
rect 32355 2400 32680 2428
rect 32355 2397 32367 2400
rect 32309 2391 32367 2397
rect 32674 2388 32680 2400
rect 32732 2388 32738 2440
rect 32953 2431 33011 2437
rect 32953 2397 32965 2431
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 31481 2363 31539 2369
rect 31481 2360 31493 2363
rect 29420 2332 31493 2360
rect 29420 2320 29426 2332
rect 31481 2329 31493 2332
rect 31527 2329 31539 2363
rect 31481 2323 31539 2329
rect 32214 2320 32220 2372
rect 32272 2360 32278 2372
rect 32968 2360 32996 2391
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33192 2400 33609 2428
rect 33192 2388 33198 2400
rect 33597 2397 33609 2400
rect 33643 2428 33655 2431
rect 33686 2428 33692 2440
rect 33643 2400 33692 2428
rect 33643 2397 33655 2400
rect 33597 2391 33655 2397
rect 33686 2388 33692 2400
rect 33744 2388 33750 2440
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34698 2428 34704 2440
rect 33836 2400 34704 2428
rect 33836 2388 33842 2400
rect 34698 2388 34704 2400
rect 34756 2428 34762 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34756 2400 34897 2428
rect 34756 2388 34762 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 34974 2388 34980 2440
rect 35032 2428 35038 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 35032 2400 35541 2428
rect 35032 2388 35038 2400
rect 35529 2397 35541 2400
rect 35575 2397 35587 2431
rect 35529 2391 35587 2397
rect 34057 2363 34115 2369
rect 34057 2360 34069 2363
rect 32272 2332 34069 2360
rect 32272 2320 32278 2332
rect 34057 2329 34069 2332
rect 34103 2329 34115 2363
rect 35544 2360 35572 2391
rect 35894 2388 35900 2440
rect 35952 2428 35958 2440
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 35952 2400 36185 2428
rect 35952 2388 35958 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 37826 2428 37832 2440
rect 37787 2400 37832 2428
rect 36173 2391 36231 2397
rect 37826 2388 37832 2400
rect 37884 2388 37890 2440
rect 36633 2363 36691 2369
rect 36633 2360 36645 2363
rect 35544 2332 36645 2360
rect 34057 2323 34115 2329
rect 36633 2329 36645 2332
rect 36679 2329 36691 2363
rect 36633 2323 36691 2329
rect 24596 2264 27016 2292
rect 24489 2255 24547 2261
rect 27062 2252 27068 2304
rect 27120 2292 27126 2304
rect 29546 2292 29552 2304
rect 27120 2264 27165 2292
rect 29507 2264 29552 2292
rect 27120 2252 27126 2264
rect 29546 2252 29552 2264
rect 29604 2252 29610 2304
rect 30190 2292 30196 2304
rect 30151 2264 30196 2292
rect 30190 2252 30196 2264
rect 30248 2252 30254 2304
rect 32122 2292 32128 2304
rect 32083 2264 32128 2292
rect 32122 2252 32128 2264
rect 32180 2252 32186 2304
rect 32766 2292 32772 2304
rect 32727 2264 32772 2292
rect 32766 2252 32772 2264
rect 32824 2252 32830 2304
rect 33410 2292 33416 2304
rect 33371 2264 33416 2292
rect 33410 2252 33416 2264
rect 33468 2252 33474 2304
rect 34514 2252 34520 2304
rect 34572 2292 34578 2304
rect 34701 2295 34759 2301
rect 34701 2292 34713 2295
rect 34572 2264 34713 2292
rect 34572 2252 34578 2264
rect 34701 2261 34713 2264
rect 34747 2261 34759 2295
rect 34701 2255 34759 2261
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35989 2295 36047 2301
rect 35989 2292 36001 2295
rect 34848 2264 36001 2292
rect 34848 2252 34854 2264
rect 35989 2261 36001 2264
rect 36035 2261 36047 2295
rect 35989 2255 36047 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 5166 2048 5172 2100
rect 5224 2088 5230 2100
rect 21910 2088 21916 2100
rect 5224 2060 21916 2088
rect 5224 2048 5230 2060
rect 21910 2048 21916 2060
rect 21968 2048 21974 2100
rect 23566 2048 23572 2100
rect 23624 2088 23630 2100
rect 29546 2088 29552 2100
rect 23624 2060 29552 2088
rect 23624 2048 23630 2060
rect 29546 2048 29552 2060
rect 29604 2048 29610 2100
rect 7098 1980 7104 2032
rect 7156 2020 7162 2032
rect 22002 2020 22008 2032
rect 7156 1992 22008 2020
rect 7156 1980 7162 1992
rect 22002 1980 22008 1992
rect 22060 1980 22066 2032
rect 23106 1980 23112 2032
rect 23164 2020 23170 2032
rect 32122 2020 32128 2032
rect 23164 1992 32128 2020
rect 23164 1980 23170 1992
rect 32122 1980 32128 1992
rect 32180 1980 32186 2032
rect 10410 1912 10416 1964
rect 10468 1952 10474 1964
rect 10468 1924 20208 1952
rect 10468 1912 10474 1924
rect 20180 1748 20208 1924
rect 20346 1912 20352 1964
rect 20404 1952 20410 1964
rect 33410 1952 33416 1964
rect 20404 1924 33416 1952
rect 20404 1912 20410 1924
rect 33410 1912 33416 1924
rect 33468 1912 33474 1964
rect 24486 1844 24492 1896
rect 24544 1884 24550 1896
rect 30190 1884 30196 1896
rect 24544 1856 30196 1884
rect 24544 1844 24550 1856
rect 30190 1844 30196 1856
rect 30248 1844 30254 1896
rect 22462 1776 22468 1828
rect 22520 1816 22526 1828
rect 32766 1816 32772 1828
rect 22520 1788 32772 1816
rect 22520 1776 22526 1788
rect 32766 1776 32772 1788
rect 32824 1776 32830 1828
rect 24854 1748 24860 1760
rect 20180 1720 24860 1748
rect 24854 1708 24860 1720
rect 24912 1708 24918 1760
rect 22646 1640 22652 1692
rect 22704 1680 22710 1692
rect 34790 1680 34796 1692
rect 22704 1652 34796 1680
rect 22704 1640 22710 1652
rect 34790 1640 34796 1652
rect 34848 1640 34854 1692
rect 24394 1368 24400 1420
rect 24452 1408 24458 1420
rect 25958 1408 25964 1420
rect 24452 1380 25964 1408
rect 24452 1368 24458 1380
rect 25958 1368 25964 1380
rect 26016 1368 26022 1420
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 8392 37451 8444 37460
rect 8392 37417 8401 37451
rect 8401 37417 8435 37451
rect 8435 37417 8444 37451
rect 8392 37408 8444 37417
rect 16120 37451 16172 37460
rect 16120 37417 16129 37451
rect 16129 37417 16163 37451
rect 16163 37417 16172 37451
rect 16120 37408 16172 37417
rect 664 37204 716 37256
rect 1308 37204 1360 37256
rect 2872 37204 2924 37256
rect 3976 37204 4028 37256
rect 5080 37204 5132 37256
rect 6184 37204 6236 37256
rect 7288 37204 7340 37256
rect 8392 37204 8444 37256
rect 9496 37204 9548 37256
rect 10600 37204 10652 37256
rect 11704 37204 11756 37256
rect 12808 37204 12860 37256
rect 13912 37204 13964 37256
rect 15016 37204 15068 37256
rect 31484 37315 31536 37324
rect 31484 37281 31493 37315
rect 31493 37281 31527 37315
rect 31527 37281 31536 37315
rect 31484 37272 31536 37281
rect 17224 37204 17276 37256
rect 18328 37204 18380 37256
rect 19432 37204 19484 37256
rect 20536 37204 20588 37256
rect 21824 37247 21876 37256
rect 21824 37213 21833 37247
rect 21833 37213 21867 37247
rect 21867 37213 21876 37247
rect 21824 37204 21876 37213
rect 23020 37204 23072 37256
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 25136 37247 25188 37256
rect 25136 37213 25145 37247
rect 25145 37213 25179 37247
rect 25179 37213 25188 37247
rect 25136 37204 25188 37213
rect 27252 37247 27304 37256
rect 4620 37136 4672 37188
rect 1952 37111 2004 37120
rect 1952 37077 1961 37111
rect 1961 37077 1995 37111
rect 1995 37077 2004 37111
rect 1952 37068 2004 37077
rect 3148 37111 3200 37120
rect 3148 37077 3157 37111
rect 3157 37077 3191 37111
rect 3191 37077 3200 37111
rect 3148 37068 3200 37077
rect 4712 37068 4764 37120
rect 10324 37136 10376 37188
rect 6368 37111 6420 37120
rect 6368 37077 6377 37111
rect 6377 37077 6411 37111
rect 6411 37077 6420 37111
rect 6368 37068 6420 37077
rect 7380 37111 7432 37120
rect 7380 37077 7389 37111
rect 7389 37077 7423 37111
rect 7423 37077 7432 37111
rect 7380 37068 7432 37077
rect 8944 37111 8996 37120
rect 8944 37077 8953 37111
rect 8953 37077 8987 37111
rect 8987 37077 8996 37111
rect 8944 37068 8996 37077
rect 9588 37111 9640 37120
rect 9588 37077 9597 37111
rect 9597 37077 9631 37111
rect 9631 37077 9640 37111
rect 9588 37068 9640 37077
rect 10692 37111 10744 37120
rect 10692 37077 10701 37111
rect 10701 37077 10735 37111
rect 10735 37077 10744 37111
rect 10692 37068 10744 37077
rect 11520 37068 11572 37120
rect 15844 37136 15896 37188
rect 14096 37111 14148 37120
rect 14096 37077 14105 37111
rect 14105 37077 14139 37111
rect 14139 37077 14148 37111
rect 14096 37068 14148 37077
rect 15108 37111 15160 37120
rect 15108 37077 15117 37111
rect 15117 37077 15151 37111
rect 15151 37077 15160 37111
rect 15108 37068 15160 37077
rect 16764 37068 16816 37120
rect 27252 37213 27261 37247
rect 27261 37213 27295 37247
rect 27295 37213 27304 37247
rect 27252 37204 27304 37213
rect 28172 37204 28224 37256
rect 29368 37204 29420 37256
rect 30380 37204 30432 37256
rect 32864 37247 32916 37256
rect 32864 37213 32873 37247
rect 32873 37213 32907 37247
rect 32907 37213 32916 37247
rect 32864 37204 32916 37213
rect 33876 37247 33928 37256
rect 33876 37213 33885 37247
rect 33885 37213 33919 37247
rect 33919 37213 33928 37247
rect 33876 37204 33928 37213
rect 34796 37204 34848 37256
rect 35900 37204 35952 37256
rect 37372 37204 37424 37256
rect 18420 37111 18472 37120
rect 18420 37077 18429 37111
rect 18429 37077 18463 37111
rect 18463 37077 18472 37111
rect 18420 37068 18472 37077
rect 19432 37068 19484 37120
rect 20628 37111 20680 37120
rect 20628 37077 20637 37111
rect 20637 37077 20671 37111
rect 20671 37077 20680 37111
rect 20628 37068 20680 37077
rect 21640 37068 21692 37120
rect 22744 37068 22796 37120
rect 23848 37068 23900 37120
rect 24952 37068 25004 37120
rect 26148 37068 26200 37120
rect 26240 37068 26292 37120
rect 27160 37068 27212 37120
rect 28264 37068 28316 37120
rect 29460 37068 29512 37120
rect 30472 37068 30524 37120
rect 31760 37068 31812 37120
rect 32680 37068 32732 37120
rect 33784 37068 33836 37120
rect 34888 37068 34940 37120
rect 35992 37068 36044 37120
rect 37096 37068 37148 37120
rect 38016 37111 38068 37120
rect 38016 37077 38025 37111
rect 38025 37077 38059 37111
rect 38059 37077 38068 37111
rect 38016 37068 38068 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 1768 36864 1820 36916
rect 2872 36907 2924 36916
rect 2872 36873 2881 36907
rect 2881 36873 2915 36907
rect 2915 36873 2924 36907
rect 2872 36864 2924 36873
rect 3976 36907 4028 36916
rect 3976 36873 3985 36907
rect 3985 36873 4019 36907
rect 4019 36873 4028 36907
rect 3976 36864 4028 36873
rect 5080 36907 5132 36916
rect 5080 36873 5089 36907
rect 5089 36873 5123 36907
rect 5123 36873 5132 36907
rect 5080 36864 5132 36873
rect 6184 36864 6236 36916
rect 7288 36907 7340 36916
rect 7288 36873 7297 36907
rect 7297 36873 7331 36907
rect 7331 36873 7340 36907
rect 7288 36864 7340 36873
rect 9496 36907 9548 36916
rect 9496 36873 9505 36907
rect 9505 36873 9539 36907
rect 9539 36873 9548 36907
rect 9496 36864 9548 36873
rect 10600 36907 10652 36916
rect 10600 36873 10609 36907
rect 10609 36873 10643 36907
rect 10643 36873 10652 36907
rect 10600 36864 10652 36873
rect 11704 36907 11756 36916
rect 11704 36873 11713 36907
rect 11713 36873 11747 36907
rect 11747 36873 11756 36907
rect 11704 36864 11756 36873
rect 12808 36907 12860 36916
rect 12808 36873 12817 36907
rect 12817 36873 12851 36907
rect 12851 36873 12860 36907
rect 12808 36864 12860 36873
rect 13912 36907 13964 36916
rect 13912 36873 13921 36907
rect 13921 36873 13955 36907
rect 13955 36873 13964 36907
rect 13912 36864 13964 36873
rect 15016 36907 15068 36916
rect 15016 36873 15025 36907
rect 15025 36873 15059 36907
rect 15059 36873 15068 36907
rect 15016 36864 15068 36873
rect 17224 36907 17276 36916
rect 17224 36873 17233 36907
rect 17233 36873 17267 36907
rect 17267 36873 17276 36907
rect 17224 36864 17276 36873
rect 18328 36907 18380 36916
rect 18328 36873 18337 36907
rect 18337 36873 18371 36907
rect 18371 36873 18380 36907
rect 18328 36864 18380 36873
rect 19340 36907 19392 36916
rect 19340 36873 19349 36907
rect 19349 36873 19383 36907
rect 19383 36873 19392 36907
rect 19340 36864 19392 36873
rect 20536 36907 20588 36916
rect 20536 36873 20545 36907
rect 20545 36873 20579 36907
rect 20579 36873 20588 36907
rect 20536 36864 20588 36873
rect 38200 36864 38252 36916
rect 2412 36728 2464 36780
rect 37832 36771 37884 36780
rect 37832 36737 37841 36771
rect 37841 36737 37875 36771
rect 37875 36737 37884 36771
rect 37832 36728 37884 36737
rect 38016 36728 38068 36780
rect 19984 36524 20036 36576
rect 21824 36567 21876 36576
rect 21824 36533 21833 36567
rect 21833 36533 21867 36567
rect 21867 36533 21876 36567
rect 21824 36524 21876 36533
rect 23020 36524 23072 36576
rect 25136 36524 25188 36576
rect 26148 36524 26200 36576
rect 27252 36524 27304 36576
rect 28172 36567 28224 36576
rect 28172 36533 28181 36567
rect 28181 36533 28215 36567
rect 28215 36533 28224 36567
rect 28172 36524 28224 36533
rect 29368 36567 29420 36576
rect 29368 36533 29377 36567
rect 29377 36533 29411 36567
rect 29411 36533 29420 36567
rect 29368 36524 29420 36533
rect 30380 36567 30432 36576
rect 30380 36533 30389 36567
rect 30389 36533 30423 36567
rect 30423 36533 30432 36567
rect 30380 36524 30432 36533
rect 32864 36524 32916 36576
rect 33876 36524 33928 36576
rect 34796 36567 34848 36576
rect 34796 36533 34805 36567
rect 34805 36533 34839 36567
rect 34839 36533 34848 36567
rect 34796 36524 34848 36533
rect 35900 36567 35952 36576
rect 35900 36533 35909 36567
rect 35909 36533 35943 36567
rect 35943 36533 35952 36567
rect 37372 36567 37424 36576
rect 35900 36524 35952 36533
rect 37372 36533 37381 36567
rect 37381 36533 37415 36567
rect 37415 36533 37424 36567
rect 37372 36524 37424 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1308 36320 1360 36372
rect 39304 36320 39356 36372
rect 2412 35980 2464 36032
rect 37280 36023 37332 36032
rect 37280 35989 37289 36023
rect 37289 35989 37323 36023
rect 37323 35989 37332 36023
rect 37280 35980 37332 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 1584 30200 1636 30252
rect 2044 30107 2096 30116
rect 2044 30073 2053 30107
rect 2053 30073 2087 30107
rect 2087 30073 2096 30107
rect 2044 30064 2096 30073
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3148 22040 3200 22092
rect 7564 22040 7616 22092
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 11428 20816 11480 20868
rect 12256 20748 12308 20800
rect 13360 20791 13412 20800
rect 13360 20757 13369 20791
rect 13369 20757 13403 20791
rect 13403 20757 13412 20791
rect 13360 20748 13412 20757
rect 16580 20791 16632 20800
rect 16580 20757 16589 20791
rect 16589 20757 16623 20791
rect 16623 20757 16632 20791
rect 16580 20748 16632 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 10324 20544 10376 20596
rect 16764 20544 16816 20596
rect 18420 20544 18472 20596
rect 10232 20408 10284 20460
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12256 20408 12308 20417
rect 13360 20383 13412 20392
rect 13360 20349 13369 20383
rect 13369 20349 13403 20383
rect 13403 20349 13412 20383
rect 13360 20340 13412 20349
rect 16304 20340 16356 20392
rect 17408 20272 17460 20324
rect 9404 20204 9456 20256
rect 10600 20204 10652 20256
rect 12900 20247 12952 20256
rect 12900 20213 12909 20247
rect 12909 20213 12943 20247
rect 12943 20213 12952 20247
rect 12900 20204 12952 20213
rect 16672 20247 16724 20256
rect 16672 20213 16681 20247
rect 16681 20213 16715 20247
rect 16715 20213 16724 20247
rect 16672 20204 16724 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4712 20000 4764 20052
rect 8300 20000 8352 20052
rect 9588 20000 9640 20052
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 15844 20000 15896 20052
rect 11704 19907 11756 19916
rect 11704 19873 11713 19907
rect 11713 19873 11747 19907
rect 11747 19873 11756 19907
rect 11704 19864 11756 19873
rect 12256 19864 12308 19916
rect 16672 19796 16724 19848
rect 19432 20000 19484 20052
rect 17408 19907 17460 19916
rect 17408 19873 17417 19907
rect 17417 19873 17451 19907
rect 17451 19873 17460 19907
rect 17408 19864 17460 19873
rect 11428 19728 11480 19780
rect 13820 19728 13872 19780
rect 16580 19728 16632 19780
rect 7656 19660 7708 19712
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10416 19660 10468 19669
rect 11152 19703 11204 19712
rect 11152 19669 11161 19703
rect 11161 19669 11195 19703
rect 11195 19669 11204 19703
rect 11152 19660 11204 19669
rect 11796 19660 11848 19712
rect 13728 19660 13780 19712
rect 15200 19703 15252 19712
rect 15200 19669 15209 19703
rect 15209 19669 15243 19703
rect 15243 19669 15252 19703
rect 15200 19660 15252 19669
rect 15660 19660 15712 19712
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 16856 19703 16908 19712
rect 16856 19669 16865 19703
rect 16865 19669 16899 19703
rect 16899 19669 16908 19703
rect 16856 19660 16908 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 2964 19456 3016 19508
rect 4712 19456 4764 19508
rect 8300 19456 8352 19508
rect 10232 19499 10284 19508
rect 10232 19465 10241 19499
rect 10241 19465 10275 19499
rect 10275 19465 10284 19499
rect 10232 19456 10284 19465
rect 11520 19456 11572 19508
rect 12808 19456 12860 19508
rect 10692 19388 10744 19440
rect 13820 19388 13872 19440
rect 15108 19388 15160 19440
rect 7656 19320 7708 19372
rect 9680 19320 9732 19372
rect 12716 19320 12768 19372
rect 13912 19320 13964 19372
rect 20628 19456 20680 19508
rect 4068 19295 4120 19304
rect 3332 19116 3384 19168
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 5540 19252 5592 19304
rect 6368 19252 6420 19304
rect 8944 19295 8996 19304
rect 8944 19261 8953 19295
rect 8953 19261 8987 19295
rect 8987 19261 8996 19295
rect 8944 19252 8996 19261
rect 10692 19295 10744 19304
rect 7932 19184 7984 19236
rect 10692 19261 10701 19295
rect 10701 19261 10735 19295
rect 10735 19261 10744 19295
rect 10692 19252 10744 19261
rect 10600 19184 10652 19236
rect 11980 19252 12032 19304
rect 11704 19184 11756 19236
rect 17316 19252 17368 19304
rect 17500 19295 17552 19304
rect 17500 19261 17509 19295
rect 17509 19261 17543 19295
rect 17543 19261 17552 19295
rect 17500 19252 17552 19261
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7288 19116 7340 19125
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 11060 19116 11112 19168
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4068 18844 4120 18896
rect 5908 18819 5960 18828
rect 5908 18785 5917 18819
rect 5917 18785 5951 18819
rect 5951 18785 5960 18819
rect 5908 18776 5960 18785
rect 5540 18708 5592 18760
rect 7380 18912 7432 18964
rect 9496 18912 9548 18964
rect 12716 18955 12768 18964
rect 12716 18921 12725 18955
rect 12725 18921 12759 18955
rect 12759 18921 12768 18955
rect 12716 18912 12768 18921
rect 17408 18912 17460 18964
rect 9312 18844 9364 18896
rect 11152 18844 11204 18896
rect 7932 18819 7984 18828
rect 3700 18640 3752 18692
rect 5172 18640 5224 18692
rect 5908 18640 5960 18692
rect 7932 18785 7941 18819
rect 7941 18785 7975 18819
rect 7975 18785 7984 18819
rect 7932 18776 7984 18785
rect 9680 18776 9732 18828
rect 8300 18708 8352 18760
rect 8852 18708 8904 18760
rect 11060 18708 11112 18760
rect 12900 18776 12952 18828
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 16856 18708 16908 18760
rect 9588 18640 9640 18692
rect 3424 18572 3476 18624
rect 5356 18615 5408 18624
rect 5356 18581 5365 18615
rect 5365 18581 5399 18615
rect 5399 18581 5408 18615
rect 5356 18572 5408 18581
rect 7104 18572 7156 18624
rect 7748 18615 7800 18624
rect 7748 18581 7757 18615
rect 7757 18581 7791 18615
rect 7791 18581 7800 18615
rect 7748 18572 7800 18581
rect 9220 18572 9272 18624
rect 14372 18572 14424 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4620 18368 4672 18420
rect 8392 18411 8444 18420
rect 8392 18377 8401 18411
rect 8401 18377 8435 18411
rect 8435 18377 8444 18411
rect 8392 18368 8444 18377
rect 8944 18368 8996 18420
rect 7748 18300 7800 18352
rect 8208 18300 8260 18352
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 7288 18232 7340 18284
rect 8484 18232 8536 18284
rect 9956 18275 10008 18284
rect 9956 18241 9965 18275
rect 9965 18241 9999 18275
rect 9999 18241 10008 18275
rect 9956 18232 10008 18241
rect 3792 18164 3844 18216
rect 5908 18164 5960 18216
rect 2596 18071 2648 18080
rect 2596 18037 2605 18071
rect 2605 18037 2639 18071
rect 2639 18037 2648 18071
rect 2596 18028 2648 18037
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 6644 18071 6696 18080
rect 6644 18037 6653 18071
rect 6653 18037 6687 18071
rect 6687 18037 6696 18071
rect 6644 18028 6696 18037
rect 6736 18028 6788 18080
rect 10140 18071 10192 18080
rect 10140 18037 10149 18071
rect 10149 18037 10183 18071
rect 10183 18037 10192 18071
rect 10140 18028 10192 18037
rect 10324 18028 10376 18080
rect 10692 18028 10744 18080
rect 11520 18028 11572 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 11980 18028 12032 18080
rect 17316 18028 17368 18080
rect 17868 18028 17920 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4620 17824 4672 17876
rect 8300 17824 8352 17876
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 5356 17620 5408 17672
rect 7104 17620 7156 17672
rect 2872 17484 2924 17536
rect 4620 17484 4672 17536
rect 6552 17527 6604 17536
rect 6552 17493 6561 17527
rect 6561 17493 6595 17527
rect 6595 17493 6604 17527
rect 6552 17484 6604 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 18052 17144 18104 17196
rect 13728 17076 13780 17128
rect 22284 16940 22336 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 5540 16575 5592 16584
rect 5540 16541 5549 16575
rect 5549 16541 5583 16575
rect 5583 16541 5592 16575
rect 5540 16532 5592 16541
rect 5908 16600 5960 16652
rect 8944 16575 8996 16584
rect 8944 16541 8953 16575
rect 8953 16541 8987 16575
rect 8987 16541 8996 16575
rect 8944 16532 8996 16541
rect 13728 16532 13780 16584
rect 9404 16464 9456 16516
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 12532 16464 12584 16516
rect 15200 16532 15252 16584
rect 19248 16464 19300 16516
rect 13544 16439 13596 16448
rect 13544 16405 13553 16439
rect 13553 16405 13587 16439
rect 13587 16405 13596 16439
rect 13544 16396 13596 16405
rect 15660 16396 15712 16448
rect 19340 16396 19392 16448
rect 19432 16396 19484 16448
rect 27252 16600 27304 16652
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2596 16192 2648 16244
rect 17868 16192 17920 16244
rect 6644 16167 6696 16176
rect 6644 16133 6678 16167
rect 6678 16133 6696 16167
rect 6644 16124 6696 16133
rect 9312 16124 9364 16176
rect 12808 16167 12860 16176
rect 12808 16133 12842 16167
rect 12842 16133 12860 16167
rect 12808 16124 12860 16133
rect 8944 16056 8996 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 6184 15988 6236 16040
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 13728 15988 13780 16040
rect 19432 15920 19484 15972
rect 21088 15988 21140 16040
rect 2780 15852 2832 15904
rect 3976 15852 4028 15904
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 11980 15852 12032 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13360 15648 13412 15700
rect 19340 15580 19392 15632
rect 8944 15512 8996 15564
rect 9312 15555 9364 15564
rect 9312 15521 9321 15555
rect 9321 15521 9355 15555
rect 9355 15521 9364 15555
rect 9312 15512 9364 15521
rect 29368 15580 29420 15632
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 4620 15444 4672 15496
rect 6184 15487 6236 15496
rect 6184 15453 6193 15487
rect 6193 15453 6227 15487
rect 6227 15453 6236 15487
rect 6184 15444 6236 15453
rect 6736 15444 6788 15496
rect 13728 15444 13780 15496
rect 2780 15376 2832 15428
rect 9588 15419 9640 15428
rect 9588 15385 9622 15419
rect 9622 15385 9640 15419
rect 9588 15376 9640 15385
rect 2872 15308 2924 15360
rect 3332 15308 3384 15360
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 8116 15308 8168 15360
rect 8392 15308 8444 15360
rect 12532 15376 12584 15428
rect 14096 15376 14148 15428
rect 16212 15376 16264 15428
rect 15016 15308 15068 15360
rect 19984 15444 20036 15496
rect 21088 15555 21140 15564
rect 21088 15521 21097 15555
rect 21097 15521 21131 15555
rect 21131 15521 21140 15555
rect 21088 15512 21140 15521
rect 20720 15444 20772 15496
rect 17684 15376 17736 15428
rect 20260 15376 20312 15428
rect 21548 15376 21600 15428
rect 17500 15351 17552 15360
rect 17500 15317 17509 15351
rect 17509 15317 17543 15351
rect 17543 15317 17552 15351
rect 17500 15308 17552 15317
rect 18696 15308 18748 15360
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 22284 15308 22336 15360
rect 31484 15308 31536 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 2780 15104 2832 15156
rect 6552 15104 6604 15156
rect 3792 15036 3844 15088
rect 9496 15104 9548 15156
rect 18052 15147 18104 15156
rect 18052 15113 18061 15147
rect 18061 15113 18095 15147
rect 18095 15113 18104 15147
rect 18052 15104 18104 15113
rect 3240 14968 3292 15020
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 15108 14968 15160 15020
rect 22284 15147 22336 15156
rect 22284 15113 22293 15147
rect 22293 15113 22327 15147
rect 22327 15113 22336 15147
rect 22284 15104 22336 15113
rect 19156 14968 19208 15020
rect 6184 14900 6236 14952
rect 12532 14943 12584 14952
rect 3884 14807 3936 14816
rect 3884 14773 3893 14807
rect 3893 14773 3927 14807
rect 3927 14773 3936 14807
rect 3884 14764 3936 14773
rect 12532 14909 12541 14943
rect 12541 14909 12575 14943
rect 12575 14909 12584 14943
rect 12532 14900 12584 14909
rect 13728 14900 13780 14952
rect 17500 14900 17552 14952
rect 30380 15036 30432 15088
rect 19984 14968 20036 15020
rect 20720 14900 20772 14952
rect 20812 14900 20864 14952
rect 21088 14943 21140 14952
rect 21088 14909 21097 14943
rect 21097 14909 21131 14943
rect 21131 14909 21140 14943
rect 21916 14968 21968 15020
rect 21088 14900 21140 14909
rect 6736 14764 6788 14816
rect 8300 14764 8352 14816
rect 13636 14764 13688 14816
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 15016 14764 15068 14816
rect 22008 14832 22060 14884
rect 22376 14943 22428 14952
rect 22376 14909 22385 14943
rect 22385 14909 22419 14943
rect 22419 14909 22428 14943
rect 22376 14900 22428 14909
rect 24400 14832 24452 14884
rect 15752 14807 15804 14816
rect 15752 14773 15761 14807
rect 15761 14773 15795 14807
rect 15795 14773 15804 14807
rect 15752 14764 15804 14773
rect 19248 14764 19300 14816
rect 20076 14764 20128 14816
rect 20812 14764 20864 14816
rect 23020 14807 23072 14816
rect 23020 14773 23029 14807
rect 23029 14773 23063 14807
rect 23063 14773 23072 14807
rect 23020 14764 23072 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3884 14560 3936 14612
rect 14004 14560 14056 14612
rect 14096 14560 14148 14612
rect 16212 14560 16264 14612
rect 19156 14560 19208 14612
rect 3792 14424 3844 14476
rect 12532 14424 12584 14476
rect 13728 14424 13780 14476
rect 6184 14356 6236 14408
rect 9312 14356 9364 14408
rect 14372 14399 14424 14408
rect 14372 14365 14406 14399
rect 14406 14365 14424 14399
rect 14372 14356 14424 14365
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 20996 14467 21048 14476
rect 20996 14433 21005 14467
rect 21005 14433 21039 14467
rect 21039 14433 21048 14467
rect 20996 14424 21048 14433
rect 21088 14467 21140 14476
rect 21088 14433 21097 14467
rect 21097 14433 21131 14467
rect 21131 14433 21140 14467
rect 21088 14424 21140 14433
rect 22376 14424 22428 14476
rect 20076 14399 20128 14408
rect 20076 14365 20085 14399
rect 20085 14365 20119 14399
rect 20119 14365 20128 14399
rect 20076 14356 20128 14365
rect 28172 14356 28224 14408
rect 5540 14288 5592 14340
rect 5724 14331 5776 14340
rect 5724 14297 5758 14331
rect 5758 14297 5776 14331
rect 10140 14331 10192 14340
rect 5724 14288 5776 14297
rect 10140 14297 10158 14331
rect 10158 14297 10192 14331
rect 10140 14288 10192 14297
rect 13912 14288 13964 14340
rect 20720 14288 20772 14340
rect 21640 14288 21692 14340
rect 24124 14288 24176 14340
rect 4436 14263 4488 14272
rect 4436 14229 4445 14263
rect 4445 14229 4479 14263
rect 4479 14229 4488 14263
rect 4436 14220 4488 14229
rect 6828 14263 6880 14272
rect 6828 14229 6837 14263
rect 6837 14229 6871 14263
rect 6871 14229 6880 14263
rect 6828 14220 6880 14229
rect 10416 14220 10468 14272
rect 10600 14220 10652 14272
rect 16488 14220 16540 14272
rect 19340 14220 19392 14272
rect 22008 14220 22060 14272
rect 22192 14263 22244 14272
rect 22192 14229 22201 14263
rect 22201 14229 22235 14263
rect 22235 14229 22244 14263
rect 22192 14220 22244 14229
rect 24308 14220 24360 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 6828 14016 6880 14068
rect 10508 14016 10560 14068
rect 17684 14016 17736 14068
rect 19432 14016 19484 14068
rect 20720 14016 20772 14068
rect 21180 14016 21232 14068
rect 22192 14016 22244 14068
rect 4436 13948 4488 14000
rect 19340 13948 19392 14000
rect 25136 13948 25188 14000
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 8208 13812 8260 13864
rect 13728 13880 13780 13932
rect 19248 13923 19300 13932
rect 19248 13889 19257 13923
rect 19257 13889 19291 13923
rect 19291 13889 19300 13923
rect 19248 13880 19300 13889
rect 20536 13880 20588 13932
rect 22376 13880 22428 13932
rect 20812 13812 20864 13864
rect 21088 13855 21140 13864
rect 21088 13821 21097 13855
rect 21097 13821 21131 13855
rect 21131 13821 21140 13855
rect 21088 13812 21140 13821
rect 20904 13744 20956 13796
rect 10416 13719 10468 13728
rect 10416 13685 10425 13719
rect 10425 13685 10459 13719
rect 10459 13685 10468 13719
rect 10416 13676 10468 13685
rect 13636 13676 13688 13728
rect 19524 13676 19576 13728
rect 20168 13676 20220 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 15108 13472 15160 13524
rect 20996 13472 21048 13524
rect 21180 13515 21232 13524
rect 21180 13481 21189 13515
rect 21189 13481 21223 13515
rect 21223 13481 21232 13515
rect 21180 13472 21232 13481
rect 10324 13404 10376 13456
rect 12532 13336 12584 13388
rect 14004 13404 14056 13456
rect 19432 13404 19484 13456
rect 19524 13404 19576 13456
rect 25136 13404 25188 13456
rect 23480 13336 23532 13388
rect 11060 13268 11112 13320
rect 11428 13268 11480 13320
rect 17224 13268 17276 13320
rect 20168 13311 20220 13320
rect 20168 13277 20177 13311
rect 20177 13277 20211 13311
rect 20211 13277 20220 13311
rect 20168 13268 20220 13277
rect 5264 13243 5316 13252
rect 5264 13209 5273 13243
rect 5273 13209 5307 13243
rect 5307 13209 5316 13243
rect 10416 13243 10468 13252
rect 5264 13200 5316 13209
rect 10416 13209 10425 13243
rect 10425 13209 10459 13243
rect 10459 13209 10468 13243
rect 10416 13200 10468 13209
rect 13544 13200 13596 13252
rect 27620 13200 27672 13252
rect 6736 13175 6788 13184
rect 6736 13141 6745 13175
rect 6745 13141 6779 13175
rect 6779 13141 6788 13175
rect 6736 13132 6788 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 11060 12928 11112 12980
rect 17224 12928 17276 12980
rect 25596 12928 25648 12980
rect 2872 12860 2924 12912
rect 6736 12860 6788 12912
rect 9220 12903 9272 12912
rect 2964 12792 3016 12844
rect 8852 12792 8904 12844
rect 9220 12869 9254 12903
rect 9254 12869 9272 12903
rect 9220 12860 9272 12869
rect 15568 12792 15620 12844
rect 7104 12767 7156 12776
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 14280 12724 14332 12776
rect 3148 12588 3200 12640
rect 9956 12588 10008 12640
rect 19340 12588 19392 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 8116 12384 8168 12436
rect 15568 12384 15620 12436
rect 20904 12384 20956 12436
rect 16304 12316 16356 12368
rect 20076 12248 20128 12300
rect 2872 12180 2924 12232
rect 7104 12180 7156 12232
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 20352 12180 20404 12232
rect 2412 12112 2464 12164
rect 7288 12112 7340 12164
rect 11336 12112 11388 12164
rect 18788 12112 18840 12164
rect 19984 12112 20036 12164
rect 20628 12112 20680 12164
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 10232 12044 10284 12096
rect 12072 12044 12124 12096
rect 20168 12044 20220 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 5172 11840 5224 11892
rect 16212 11840 16264 11892
rect 17868 11840 17920 11892
rect 18788 11883 18840 11892
rect 18788 11849 18797 11883
rect 18797 11849 18831 11883
rect 18831 11849 18840 11883
rect 18788 11840 18840 11849
rect 19340 11840 19392 11892
rect 19800 11883 19852 11892
rect 19800 11849 19809 11883
rect 19809 11849 19843 11883
rect 19843 11849 19852 11883
rect 19800 11840 19852 11849
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 2872 11747 2924 11756
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 2872 11704 2924 11713
rect 4712 11704 4764 11756
rect 7104 11772 7156 11824
rect 14004 11772 14056 11824
rect 29000 11840 29052 11892
rect 7840 11704 7892 11756
rect 10048 11704 10100 11756
rect 17868 11704 17920 11756
rect 19984 11704 20036 11756
rect 20996 11704 21048 11756
rect 14280 11679 14332 11688
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 19800 11636 19852 11688
rect 20720 11568 20772 11620
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 26148 11568 26200 11620
rect 4804 11500 4856 11552
rect 7748 11543 7800 11552
rect 7748 11509 7757 11543
rect 7757 11509 7791 11543
rect 7791 11509 7800 11543
rect 7748 11500 7800 11509
rect 11704 11500 11756 11552
rect 18236 11543 18288 11552
rect 18236 11509 18245 11543
rect 18245 11509 18279 11543
rect 18279 11509 18288 11543
rect 18236 11500 18288 11509
rect 18328 11500 18380 11552
rect 19156 11500 19208 11552
rect 37372 11772 37424 11824
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 7380 11296 7432 11348
rect 10324 11296 10376 11348
rect 19248 11296 19300 11348
rect 20168 11296 20220 11348
rect 3608 11228 3660 11280
rect 13728 11228 13780 11280
rect 18328 11228 18380 11280
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 2872 11092 2924 11144
rect 7104 11092 7156 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 20076 11160 20128 11212
rect 18696 11135 18748 11144
rect 2688 11024 2740 11076
rect 6276 11067 6328 11076
rect 6276 11033 6294 11067
rect 6294 11033 6328 11067
rect 6276 11024 6328 11033
rect 8760 11024 8812 11076
rect 10784 11024 10836 11076
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 18788 11092 18840 11144
rect 18144 11024 18196 11076
rect 18236 11024 18288 11076
rect 34796 11092 34848 11144
rect 20168 11024 20220 11076
rect 37832 11024 37884 11076
rect 17960 10956 18012 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 2872 10795 2924 10804
rect 2872 10761 2881 10795
rect 2881 10761 2915 10795
rect 2915 10761 2924 10795
rect 2872 10752 2924 10761
rect 3424 10752 3476 10804
rect 8208 10752 8260 10804
rect 8300 10752 8352 10804
rect 5264 10684 5316 10736
rect 10048 10684 10100 10736
rect 3976 10616 4028 10668
rect 10140 10616 10192 10668
rect 10968 10616 11020 10668
rect 18696 10752 18748 10804
rect 19248 10795 19300 10804
rect 19248 10761 19257 10795
rect 19257 10761 19291 10795
rect 19291 10761 19300 10795
rect 19248 10752 19300 10761
rect 19984 10795 20036 10804
rect 19984 10761 19993 10795
rect 19993 10761 20027 10795
rect 20027 10761 20036 10795
rect 19984 10752 20036 10761
rect 20168 10752 20220 10804
rect 18052 10684 18104 10736
rect 10876 10548 10928 10600
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 17960 10616 18012 10668
rect 18880 10616 18932 10668
rect 20352 10659 20404 10668
rect 20352 10625 20361 10659
rect 20361 10625 20395 10659
rect 20395 10625 20404 10659
rect 20352 10616 20404 10625
rect 18236 10480 18288 10532
rect 19984 10548 20036 10600
rect 35900 10548 35952 10600
rect 20076 10480 20128 10532
rect 11060 10412 11112 10464
rect 15752 10412 15804 10464
rect 19432 10412 19484 10464
rect 20536 10412 20588 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10968 10208 11020 10260
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 18144 10140 18196 10192
rect 18880 10208 18932 10260
rect 19984 10208 20036 10260
rect 18604 10140 18656 10192
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 19984 10072 20036 10124
rect 2872 10004 2924 10056
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 15752 10004 15804 10056
rect 3792 9936 3844 9988
rect 17960 10004 18012 10056
rect 18420 10004 18472 10056
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 18880 10004 18932 10056
rect 4620 9868 4672 9920
rect 10140 9868 10192 9920
rect 20168 9936 20220 9988
rect 32864 10004 32916 10056
rect 18420 9868 18472 9920
rect 18512 9868 18564 9920
rect 19432 9868 19484 9920
rect 20720 9868 20772 9920
rect 33876 9868 33928 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 17960 9664 18012 9716
rect 18236 9664 18288 9716
rect 18696 9664 18748 9716
rect 20720 9596 20772 9648
rect 3056 9528 3108 9580
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 10968 9571 11020 9580
rect 10968 9537 10977 9571
rect 10977 9537 11011 9571
rect 11011 9537 11020 9571
rect 10968 9528 11020 9537
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 15568 9528 15620 9580
rect 19248 9528 19300 9580
rect 19340 9528 19392 9580
rect 19156 9460 19208 9512
rect 19984 9460 20036 9512
rect 2964 9392 3016 9444
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 8760 9392 8812 9401
rect 10784 9435 10836 9444
rect 10784 9401 10793 9435
rect 10793 9401 10827 9435
rect 10827 9401 10836 9435
rect 10784 9392 10836 9401
rect 17316 9392 17368 9444
rect 37280 9392 37332 9444
rect 11980 9324 12032 9376
rect 15476 9324 15528 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 3792 9163 3844 9172
rect 3792 9129 3801 9163
rect 3801 9129 3835 9163
rect 3835 9129 3844 9163
rect 3792 9120 3844 9129
rect 5540 9120 5592 9172
rect 8852 9120 8904 9172
rect 11336 9120 11388 9172
rect 15476 9120 15528 9172
rect 26516 9120 26568 9172
rect 2504 9052 2556 9104
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 2780 8916 2832 8968
rect 3148 8984 3200 9036
rect 4620 8984 4672 9036
rect 14096 9052 14148 9104
rect 19432 9095 19484 9104
rect 19432 9061 19441 9095
rect 19441 9061 19475 9095
rect 19475 9061 19484 9095
rect 19432 9052 19484 9061
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4160 8959 4212 8968
rect 2872 8848 2924 8900
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 9956 8984 10008 9036
rect 6644 8916 6696 8968
rect 13360 8984 13412 9036
rect 26240 8984 26292 9036
rect 10324 8959 10376 8968
rect 5172 8848 5224 8900
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 10508 8916 10560 8968
rect 12348 8916 12400 8968
rect 16488 8916 16540 8968
rect 27068 8916 27120 8968
rect 11796 8848 11848 8900
rect 3240 8823 3292 8832
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 6000 8823 6052 8832
rect 6000 8789 6009 8823
rect 6009 8789 6043 8823
rect 6043 8789 6052 8823
rect 6000 8780 6052 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2872 8576 2924 8628
rect 3056 8619 3108 8628
rect 3056 8585 3065 8619
rect 3065 8585 3099 8619
rect 3099 8585 3108 8619
rect 3056 8576 3108 8585
rect 4712 8619 4764 8628
rect 2780 8508 2832 8560
rect 3240 8508 3292 8560
rect 4712 8585 4721 8619
rect 4721 8585 4755 8619
rect 4755 8585 4764 8619
rect 4712 8576 4764 8585
rect 5632 8576 5684 8628
rect 6000 8576 6052 8628
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 8944 8619 8996 8628
rect 8944 8585 8953 8619
rect 8953 8585 8987 8619
rect 8987 8585 8996 8619
rect 8944 8576 8996 8585
rect 10968 8619 11020 8628
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 11704 8619 11756 8628
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 3608 8483 3660 8492
rect 3608 8449 3618 8483
rect 3618 8449 3652 8483
rect 3652 8449 3660 8483
rect 3792 8483 3844 8492
rect 3608 8440 3660 8449
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4988 8508 5040 8560
rect 3240 8372 3292 8424
rect 4160 8440 4212 8492
rect 5080 8440 5132 8492
rect 7472 8440 7524 8492
rect 9128 8508 9180 8560
rect 11428 8508 11480 8560
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 15568 8619 15620 8628
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 12072 8483 12124 8492
rect 6092 8372 6144 8424
rect 6736 8415 6788 8424
rect 6736 8381 6745 8415
rect 6745 8381 6779 8415
rect 6779 8381 6788 8415
rect 6736 8372 6788 8381
rect 5908 8304 5960 8356
rect 7840 8372 7892 8424
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 18052 8483 18104 8492
rect 14924 8372 14976 8424
rect 18052 8449 18061 8483
rect 18061 8449 18095 8483
rect 18095 8449 18104 8483
rect 18052 8440 18104 8449
rect 19984 8372 20036 8424
rect 8944 8304 8996 8356
rect 9128 8304 9180 8356
rect 10324 8304 10376 8356
rect 6920 8236 6972 8288
rect 9956 8236 10008 8288
rect 11980 8236 12032 8288
rect 18144 8236 18196 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3516 8032 3568 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 5908 8075 5960 8084
rect 5908 8041 5917 8075
rect 5917 8041 5951 8075
rect 5951 8041 5960 8075
rect 5908 8032 5960 8041
rect 6920 8032 6972 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 3240 8007 3292 8016
rect 3240 7973 3249 8007
rect 3249 7973 3283 8007
rect 3283 7973 3292 8007
rect 3240 7964 3292 7973
rect 2044 7896 2096 7948
rect 8208 7964 8260 8016
rect 2780 7828 2832 7880
rect 3148 7828 3200 7880
rect 3608 7828 3660 7880
rect 4620 7896 4672 7948
rect 10508 8032 10560 8084
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 14096 8075 14148 8084
rect 14096 8041 14105 8075
rect 14105 8041 14139 8075
rect 14139 8041 14148 8075
rect 14096 8032 14148 8041
rect 14924 7964 14976 8016
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 4804 7828 4856 7880
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6184 7871 6236 7880
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 6644 7828 6696 7880
rect 6828 7828 6880 7880
rect 11060 7896 11112 7948
rect 10508 7828 10560 7880
rect 10140 7760 10192 7812
rect 10416 7760 10468 7812
rect 10692 7760 10744 7812
rect 5724 7692 5776 7744
rect 9680 7692 9732 7744
rect 11428 7828 11480 7880
rect 13176 7828 13228 7880
rect 13820 7896 13872 7948
rect 13912 7828 13964 7880
rect 16120 8032 16172 8084
rect 18052 7964 18104 8016
rect 17224 7871 17276 7880
rect 14924 7760 14976 7812
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17316 7871 17368 7880
rect 17316 7837 17325 7871
rect 17325 7837 17359 7871
rect 17359 7837 17368 7871
rect 18052 7871 18104 7880
rect 17316 7828 17368 7837
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 16856 7735 16908 7744
rect 11244 7692 11296 7701
rect 16856 7701 16865 7735
rect 16865 7701 16899 7735
rect 16899 7701 16908 7735
rect 16856 7692 16908 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2596 7488 2648 7540
rect 3792 7531 3844 7540
rect 3792 7497 3801 7531
rect 3801 7497 3835 7531
rect 3835 7497 3844 7531
rect 3792 7488 3844 7497
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 9404 7488 9456 7540
rect 11520 7488 11572 7540
rect 14924 7531 14976 7540
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 15752 7488 15804 7540
rect 17224 7488 17276 7540
rect 20260 7531 20312 7540
rect 20260 7497 20269 7531
rect 20269 7497 20303 7531
rect 20303 7497 20312 7531
rect 20260 7488 20312 7497
rect 2872 7420 2924 7472
rect 3148 7352 3200 7404
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 4620 7352 4672 7404
rect 6184 7352 6236 7404
rect 3056 7327 3108 7336
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 5724 7284 5776 7336
rect 7748 7352 7800 7404
rect 8024 7395 8076 7404
rect 8024 7361 8033 7395
rect 8033 7361 8067 7395
rect 8067 7361 8076 7395
rect 8024 7352 8076 7361
rect 8208 7420 8260 7472
rect 9680 7463 9732 7472
rect 9680 7429 9689 7463
rect 9689 7429 9723 7463
rect 9723 7429 9732 7463
rect 9680 7420 9732 7429
rect 9956 7420 10008 7472
rect 15844 7463 15896 7472
rect 15844 7429 15853 7463
rect 15853 7429 15887 7463
rect 15887 7429 15896 7463
rect 15844 7420 15896 7429
rect 19524 7420 19576 7472
rect 10508 7395 10560 7404
rect 10508 7361 10517 7395
rect 10517 7361 10551 7395
rect 10551 7361 10560 7395
rect 10508 7352 10560 7361
rect 13728 7395 13780 7404
rect 13728 7361 13737 7395
rect 13737 7361 13771 7395
rect 13771 7361 13780 7395
rect 13728 7352 13780 7361
rect 6828 7284 6880 7336
rect 9496 7284 9548 7336
rect 11888 7284 11940 7336
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15200 7352 15252 7404
rect 19984 7352 20036 7404
rect 14096 7284 14148 7336
rect 19800 7284 19852 7336
rect 15016 7216 15068 7268
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 13820 7148 13872 7200
rect 14188 7148 14240 7200
rect 14648 7148 14700 7200
rect 16856 7148 16908 7200
rect 21456 7148 21508 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3608 6944 3660 6996
rect 5540 6944 5592 6996
rect 4344 6876 4396 6928
rect 11796 6944 11848 6996
rect 12164 6944 12216 6996
rect 6184 6876 6236 6928
rect 12808 6876 12860 6928
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 3056 6740 3108 6792
rect 5632 6740 5684 6792
rect 6828 6808 6880 6860
rect 8944 6851 8996 6860
rect 2872 6672 2924 6724
rect 3148 6604 3200 6656
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 7840 6740 7892 6792
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 11060 6808 11112 6860
rect 11796 6808 11848 6860
rect 11980 6808 12032 6860
rect 13728 6944 13780 6996
rect 14280 6944 14332 6996
rect 14556 6944 14608 6996
rect 15016 6987 15068 6996
rect 15016 6953 15025 6987
rect 15025 6953 15059 6987
rect 15059 6953 15068 6987
rect 15016 6944 15068 6953
rect 15844 6944 15896 6996
rect 19800 6987 19852 6996
rect 19800 6953 19809 6987
rect 19809 6953 19843 6987
rect 19843 6953 19852 6987
rect 19800 6944 19852 6953
rect 6920 6715 6972 6724
rect 6920 6681 6929 6715
rect 6929 6681 6963 6715
rect 6963 6681 6972 6715
rect 6920 6672 6972 6681
rect 8024 6672 8076 6724
rect 10140 6740 10192 6792
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 14372 6808 14424 6860
rect 14556 6740 14608 6792
rect 15292 6740 15344 6792
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 9588 6672 9640 6724
rect 11704 6672 11756 6724
rect 12072 6672 12124 6724
rect 6736 6604 6788 6656
rect 11980 6604 12032 6656
rect 12348 6647 12400 6656
rect 12348 6613 12357 6647
rect 12357 6613 12391 6647
rect 12391 6613 12400 6647
rect 12348 6604 12400 6613
rect 12716 6647 12768 6656
rect 12716 6613 12725 6647
rect 12725 6613 12759 6647
rect 12759 6613 12768 6647
rect 12716 6604 12768 6613
rect 13268 6604 13320 6656
rect 14188 6604 14240 6656
rect 14280 6604 14332 6656
rect 17684 6783 17736 6792
rect 16488 6647 16540 6656
rect 16488 6613 16497 6647
rect 16497 6613 16531 6647
rect 16531 6613 16540 6647
rect 16488 6604 16540 6613
rect 17684 6749 17693 6783
rect 17693 6749 17727 6783
rect 17727 6749 17736 6783
rect 17684 6740 17736 6749
rect 18052 6876 18104 6928
rect 20996 6851 21048 6860
rect 17224 6672 17276 6724
rect 17592 6604 17644 6656
rect 20996 6817 21005 6851
rect 21005 6817 21039 6851
rect 21039 6817 21048 6851
rect 20996 6808 21048 6817
rect 19524 6672 19576 6724
rect 21088 6672 21140 6724
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 22008 6740 22060 6792
rect 21732 6672 21784 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2688 6443 2740 6452
rect 2688 6409 2697 6443
rect 2697 6409 2731 6443
rect 2731 6409 2740 6443
rect 2688 6400 2740 6409
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 10508 6400 10560 6452
rect 10784 6400 10836 6452
rect 11796 6400 11848 6452
rect 11980 6400 12032 6452
rect 2872 6307 2924 6316
rect 2872 6273 2881 6307
rect 2881 6273 2915 6307
rect 2915 6273 2924 6307
rect 2872 6264 2924 6273
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 2780 6128 2832 6180
rect 7840 6196 7892 6248
rect 9036 6264 9088 6316
rect 9956 6332 10008 6384
rect 11888 6375 11940 6384
rect 11888 6341 11897 6375
rect 11897 6341 11931 6375
rect 11931 6341 11940 6375
rect 11888 6332 11940 6341
rect 12256 6332 12308 6384
rect 14372 6332 14424 6384
rect 11244 6264 11296 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11796 6307 11848 6316
rect 11796 6273 11805 6307
rect 11805 6273 11839 6307
rect 11839 6273 11848 6307
rect 11796 6264 11848 6273
rect 11980 6307 12032 6316
rect 11980 6273 12015 6307
rect 12015 6273 12032 6307
rect 11980 6264 12032 6273
rect 12624 6264 12676 6316
rect 13912 6264 13964 6316
rect 14004 6264 14056 6316
rect 11060 6196 11112 6248
rect 12164 6239 12216 6248
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 14648 6239 14700 6248
rect 14648 6205 14657 6239
rect 14657 6205 14691 6239
rect 14691 6205 14700 6239
rect 14648 6196 14700 6205
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 4344 6128 4396 6180
rect 4712 6128 4764 6180
rect 12808 6128 12860 6180
rect 9496 6060 9548 6112
rect 10600 6060 10652 6112
rect 11428 6060 11480 6112
rect 11796 6060 11848 6112
rect 13636 6060 13688 6112
rect 13820 6060 13872 6112
rect 16396 6400 16448 6452
rect 17592 6400 17644 6452
rect 17960 6400 18012 6452
rect 19340 6443 19392 6452
rect 19340 6409 19349 6443
rect 19349 6409 19383 6443
rect 19383 6409 19392 6443
rect 19340 6400 19392 6409
rect 20444 6443 20496 6452
rect 20444 6409 20453 6443
rect 20453 6409 20487 6443
rect 20487 6409 20496 6443
rect 20444 6400 20496 6409
rect 22376 6443 22428 6452
rect 22376 6409 22385 6443
rect 22385 6409 22419 6443
rect 22419 6409 22428 6443
rect 22376 6400 22428 6409
rect 15016 6375 15068 6384
rect 15016 6341 15025 6375
rect 15025 6341 15059 6375
rect 15059 6341 15068 6375
rect 15016 6332 15068 6341
rect 16488 6332 16540 6384
rect 17684 6332 17736 6384
rect 20720 6375 20772 6384
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 19156 6307 19208 6316
rect 19156 6273 19165 6307
rect 19165 6273 19199 6307
rect 19199 6273 19208 6307
rect 19156 6264 19208 6273
rect 19340 6264 19392 6316
rect 20720 6341 20729 6375
rect 20729 6341 20763 6375
rect 20763 6341 20772 6375
rect 20720 6332 20772 6341
rect 28816 6400 28868 6452
rect 22744 6375 22796 6384
rect 22744 6341 22753 6375
rect 22753 6341 22787 6375
rect 22787 6341 22796 6375
rect 22744 6332 22796 6341
rect 15108 6128 15160 6180
rect 20904 6307 20956 6316
rect 20904 6273 20949 6307
rect 20949 6273 20956 6307
rect 20904 6264 20956 6273
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 22560 6307 22612 6316
rect 21088 6264 21140 6273
rect 22560 6273 22569 6307
rect 22569 6273 22603 6307
rect 22603 6273 22612 6307
rect 22560 6264 22612 6273
rect 22008 6196 22060 6248
rect 17224 6060 17276 6112
rect 17776 6060 17828 6112
rect 18420 6060 18472 6112
rect 37832 6060 37884 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 5724 5856 5776 5908
rect 9036 5899 9088 5908
rect 9036 5865 9045 5899
rect 9045 5865 9079 5899
rect 9079 5865 9088 5899
rect 9036 5856 9088 5865
rect 7932 5720 7984 5772
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8208 5652 8260 5704
rect 12440 5856 12492 5908
rect 12624 5899 12676 5908
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 13636 5856 13688 5908
rect 15016 5856 15068 5908
rect 20352 5856 20404 5908
rect 20720 5856 20772 5908
rect 9404 5720 9456 5772
rect 9312 5652 9364 5704
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 10600 5720 10652 5772
rect 11980 5720 12032 5772
rect 12164 5720 12216 5772
rect 12440 5720 12492 5772
rect 15200 5720 15252 5772
rect 11428 5695 11480 5704
rect 9588 5584 9640 5636
rect 10876 5584 10928 5636
rect 8300 5516 8352 5568
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 12256 5652 12308 5704
rect 11244 5584 11296 5636
rect 14096 5652 14148 5704
rect 19340 5652 19392 5704
rect 20260 5695 20312 5704
rect 19064 5584 19116 5636
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 13912 5516 13964 5568
rect 19432 5516 19484 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 7288 5355 7340 5364
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 7656 5312 7708 5364
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 20628 5312 20680 5364
rect 22008 5312 22060 5364
rect 3332 5244 3384 5296
rect 17316 5244 17368 5296
rect 21364 5244 21416 5296
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 6736 5108 6788 5160
rect 8300 5176 8352 5228
rect 19340 5176 19392 5228
rect 22100 5176 22152 5228
rect 7656 5151 7708 5160
rect 7104 5040 7156 5092
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 15384 5108 15436 5160
rect 24768 5176 24820 5228
rect 7840 5040 7892 5092
rect 20536 5040 20588 5092
rect 20904 5040 20956 5092
rect 10232 4972 10284 5024
rect 17040 4972 17092 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1952 4768 2004 4820
rect 7656 4768 7708 4820
rect 9680 4768 9732 4820
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 18788 4768 18840 4820
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 21916 4768 21968 4820
rect 23480 4811 23532 4820
rect 23480 4777 23489 4811
rect 23489 4777 23523 4811
rect 23523 4777 23532 4811
rect 23480 4768 23532 4777
rect 24400 4811 24452 4820
rect 24400 4777 24409 4811
rect 24409 4777 24443 4811
rect 24443 4777 24452 4811
rect 24400 4768 24452 4777
rect 6920 4700 6972 4752
rect 7288 4700 7340 4752
rect 15108 4700 15160 4752
rect 6736 4632 6788 4684
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 9496 4564 9548 4616
rect 10692 4632 10744 4684
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 7380 4496 7432 4548
rect 15108 4564 15160 4616
rect 15844 4632 15896 4684
rect 18880 4700 18932 4752
rect 16580 4564 16632 4616
rect 17224 4564 17276 4616
rect 17408 4564 17460 4616
rect 18512 4607 18564 4616
rect 11060 4496 11112 4548
rect 11888 4496 11940 4548
rect 16488 4496 16540 4548
rect 7012 4428 7064 4480
rect 7196 4471 7248 4480
rect 7196 4437 7205 4471
rect 7205 4437 7239 4471
rect 7239 4437 7248 4471
rect 7196 4428 7248 4437
rect 11704 4471 11756 4480
rect 11704 4437 11713 4471
rect 11713 4437 11747 4471
rect 11747 4437 11756 4471
rect 11704 4428 11756 4437
rect 15660 4428 15712 4480
rect 16672 4428 16724 4480
rect 17500 4496 17552 4548
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 20168 4632 20220 4684
rect 20352 4632 20404 4684
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 22100 4564 22152 4616
rect 24768 4564 24820 4616
rect 24952 4496 25004 4548
rect 21456 4471 21508 4480
rect 21456 4437 21465 4471
rect 21465 4437 21499 4471
rect 21499 4437 21508 4471
rect 21456 4428 21508 4437
rect 21916 4428 21968 4480
rect 23204 4428 23256 4480
rect 34428 4428 34480 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 6552 4224 6604 4276
rect 6920 4224 6972 4276
rect 7196 4088 7248 4140
rect 12256 4224 12308 4276
rect 17224 4224 17276 4276
rect 17500 4224 17552 4276
rect 17684 4224 17736 4276
rect 22100 4267 22152 4276
rect 22100 4233 22109 4267
rect 22109 4233 22143 4267
rect 22143 4233 22152 4267
rect 22100 4224 22152 4233
rect 23572 4224 23624 4276
rect 9680 4156 9732 4208
rect 18052 4156 18104 4208
rect 18972 4156 19024 4208
rect 22008 4156 22060 4208
rect 23112 4156 23164 4208
rect 7104 4063 7156 4072
rect 7104 4029 7113 4063
rect 7113 4029 7147 4063
rect 7147 4029 7156 4063
rect 7104 4020 7156 4029
rect 9588 4020 9640 4072
rect 9496 3952 9548 4004
rect 5448 3884 5500 3936
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 10692 4088 10744 4140
rect 13268 4088 13320 4140
rect 15200 4088 15252 4140
rect 10600 3952 10652 4004
rect 10784 3884 10836 3936
rect 11060 4020 11112 4072
rect 11796 4063 11848 4072
rect 11796 4029 11805 4063
rect 11805 4029 11839 4063
rect 11839 4029 11848 4063
rect 11796 4020 11848 4029
rect 11888 4063 11940 4072
rect 11888 4029 11897 4063
rect 11897 4029 11931 4063
rect 11931 4029 11940 4063
rect 11888 4020 11940 4029
rect 15660 4088 15712 4140
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 16764 4088 16816 4140
rect 17132 4020 17184 4072
rect 17776 4088 17828 4140
rect 12256 3952 12308 4004
rect 15292 3952 15344 4004
rect 11244 3884 11296 3936
rect 11888 3884 11940 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 15568 3952 15620 4004
rect 16948 3952 17000 4004
rect 17592 3952 17644 4004
rect 18880 4131 18932 4140
rect 18880 4097 18889 4131
rect 18889 4097 18923 4131
rect 18923 4097 18932 4131
rect 18880 4088 18932 4097
rect 22100 4088 22152 4140
rect 22284 4131 22336 4140
rect 22284 4097 22293 4131
rect 22293 4097 22327 4131
rect 22327 4097 22336 4131
rect 22284 4088 22336 4097
rect 21824 4020 21876 4072
rect 22468 4131 22520 4140
rect 22468 4097 22477 4131
rect 22477 4097 22511 4131
rect 22511 4097 22520 4131
rect 22468 4088 22520 4097
rect 22928 4088 22980 4140
rect 23204 4088 23256 4140
rect 23756 4156 23808 4208
rect 33324 4156 33376 4208
rect 24124 4131 24176 4140
rect 19064 3995 19116 4004
rect 19064 3961 19073 3995
rect 19073 3961 19107 3995
rect 19107 3961 19116 3995
rect 19064 3952 19116 3961
rect 22744 4020 22796 4072
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 24400 4088 24452 4140
rect 24768 4088 24820 4140
rect 25596 4131 25648 4140
rect 25596 4097 25605 4131
rect 25605 4097 25639 4131
rect 25639 4097 25648 4131
rect 25596 4088 25648 4097
rect 26240 4131 26292 4140
rect 26240 4097 26249 4131
rect 26249 4097 26283 4131
rect 26283 4097 26292 4131
rect 26240 4088 26292 4097
rect 36636 4088 36688 4140
rect 16120 3884 16172 3936
rect 16304 3884 16356 3936
rect 22560 3952 22612 4004
rect 19800 3884 19852 3936
rect 20628 3884 20680 3936
rect 22100 3884 22152 3936
rect 22652 3884 22704 3936
rect 24768 3884 24820 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 9680 3680 9732 3732
rect 11888 3680 11940 3732
rect 15384 3723 15436 3732
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 15568 3723 15620 3732
rect 15568 3689 15577 3723
rect 15577 3689 15611 3723
rect 15611 3689 15620 3723
rect 15568 3680 15620 3689
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 16212 3680 16264 3732
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 17408 3680 17460 3732
rect 19156 3680 19208 3732
rect 8392 3544 8444 3596
rect 10600 3544 10652 3596
rect 6736 3476 6788 3528
rect 9680 3476 9732 3528
rect 7840 3408 7892 3460
rect 10784 3476 10836 3528
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 11796 3544 11848 3596
rect 15752 3612 15804 3664
rect 15844 3544 15896 3596
rect 16948 3612 17000 3664
rect 19432 3680 19484 3732
rect 19984 3723 20036 3732
rect 19984 3689 19993 3723
rect 19993 3689 20027 3723
rect 20027 3689 20036 3723
rect 19984 3680 20036 3689
rect 20812 3680 20864 3732
rect 21548 3723 21600 3732
rect 21548 3689 21557 3723
rect 21557 3689 21591 3723
rect 21591 3689 21600 3723
rect 21548 3680 21600 3689
rect 22100 3680 22152 3732
rect 22744 3680 22796 3732
rect 24952 3723 25004 3732
rect 24952 3689 24961 3723
rect 24961 3689 24995 3723
rect 24995 3689 25004 3723
rect 24952 3680 25004 3689
rect 26516 3723 26568 3732
rect 26516 3689 26525 3723
rect 26525 3689 26559 3723
rect 26559 3689 26568 3723
rect 26516 3680 26568 3689
rect 27068 3723 27120 3732
rect 27068 3689 27077 3723
rect 27077 3689 27111 3723
rect 27111 3689 27120 3723
rect 27068 3680 27120 3689
rect 27620 3723 27672 3732
rect 27620 3689 27629 3723
rect 27629 3689 27663 3723
rect 27663 3689 27672 3723
rect 27620 3680 27672 3689
rect 36636 3723 36688 3732
rect 36636 3689 36645 3723
rect 36645 3689 36679 3723
rect 36679 3689 36688 3723
rect 36636 3680 36688 3689
rect 11980 3476 12032 3528
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 13636 3408 13688 3460
rect 16120 3476 16172 3528
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 16396 3476 16448 3528
rect 17960 3544 18012 3596
rect 21732 3612 21784 3664
rect 16856 3476 16908 3528
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 17776 3476 17828 3528
rect 21548 3544 21600 3596
rect 18052 3408 18104 3460
rect 3976 3383 4028 3392
rect 3976 3349 3985 3383
rect 3985 3349 4019 3383
rect 4019 3349 4028 3383
rect 3976 3340 4028 3349
rect 4620 3340 4672 3392
rect 5080 3383 5132 3392
rect 5080 3349 5089 3383
rect 5089 3349 5123 3383
rect 5123 3349 5132 3383
rect 5080 3340 5132 3349
rect 5632 3383 5684 3392
rect 5632 3349 5641 3383
rect 5641 3349 5675 3383
rect 5675 3349 5684 3383
rect 5632 3340 5684 3349
rect 6920 3340 6972 3392
rect 12900 3340 12952 3392
rect 13452 3340 13504 3392
rect 15936 3340 15988 3392
rect 16028 3340 16080 3392
rect 19432 3476 19484 3528
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 21732 3519 21784 3528
rect 21732 3485 21741 3519
rect 21741 3485 21775 3519
rect 21775 3485 21784 3519
rect 21732 3476 21784 3485
rect 20260 3451 20312 3460
rect 20260 3417 20269 3451
rect 20269 3417 20303 3451
rect 20303 3417 20312 3451
rect 20260 3408 20312 3417
rect 20352 3451 20404 3460
rect 20352 3417 20361 3451
rect 20361 3417 20395 3451
rect 20395 3417 20404 3451
rect 20352 3408 20404 3417
rect 21824 3451 21876 3460
rect 21824 3417 21833 3451
rect 21833 3417 21867 3451
rect 21867 3417 21876 3451
rect 21824 3408 21876 3417
rect 22376 3544 22428 3596
rect 22928 3544 22980 3596
rect 22744 3519 22796 3528
rect 22744 3485 22753 3519
rect 22753 3485 22787 3519
rect 22787 3485 22796 3519
rect 22744 3476 22796 3485
rect 24216 3544 24268 3596
rect 22560 3408 22612 3460
rect 23296 3476 23348 3528
rect 24768 3519 24820 3528
rect 24768 3485 24777 3519
rect 24777 3485 24811 3519
rect 24811 3485 24820 3519
rect 24768 3476 24820 3485
rect 36544 3476 36596 3528
rect 22376 3340 22428 3392
rect 24308 3408 24360 3460
rect 24584 3451 24636 3460
rect 24584 3417 24593 3451
rect 24593 3417 24627 3451
rect 24627 3417 24636 3451
rect 24584 3408 24636 3417
rect 23112 3340 23164 3392
rect 24860 3408 24912 3460
rect 26056 3408 26108 3460
rect 31208 3408 31260 3460
rect 27896 3340 27948 3392
rect 28540 3340 28592 3392
rect 29552 3383 29604 3392
rect 29552 3349 29561 3383
rect 29561 3349 29595 3383
rect 29595 3349 29604 3383
rect 29552 3340 29604 3349
rect 30748 3340 30800 3392
rect 31392 3340 31444 3392
rect 33232 3383 33284 3392
rect 33232 3349 33241 3383
rect 33241 3349 33275 3383
rect 33275 3349 33284 3383
rect 33232 3340 33284 3349
rect 33692 3383 33744 3392
rect 33692 3349 33701 3383
rect 33701 3349 33735 3383
rect 33735 3349 33744 3383
rect 33692 3340 33744 3349
rect 34704 3383 34756 3392
rect 34704 3349 34713 3383
rect 34713 3349 34747 3383
rect 34747 3349 34756 3383
rect 34704 3340 34756 3349
rect 35808 3340 35860 3392
rect 35992 3383 36044 3392
rect 35992 3349 36001 3383
rect 36001 3349 36035 3383
rect 36035 3349 36044 3383
rect 35992 3340 36044 3349
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2872 3136 2924 3188
rect 2872 3000 2924 3052
rect 3976 3000 4028 3052
rect 4620 3000 4672 3052
rect 7288 3136 7340 3188
rect 10508 3136 10560 3188
rect 13636 3179 13688 3188
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 15200 3179 15252 3188
rect 5080 3000 5132 3052
rect 6736 3000 6788 3052
rect 11612 3068 11664 3120
rect 15200 3145 15209 3179
rect 15209 3145 15243 3179
rect 15243 3145 15252 3179
rect 15200 3136 15252 3145
rect 16396 3136 16448 3188
rect 16948 3136 17000 3188
rect 17316 3136 17368 3188
rect 17684 3136 17736 3188
rect 17868 3136 17920 3188
rect 18512 3136 18564 3188
rect 8392 3000 8444 3052
rect 9496 3000 9548 3052
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11244 3000 11296 3052
rect 11704 3000 11756 3052
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 15844 3068 15896 3120
rect 16304 3068 16356 3120
rect 18052 3068 18104 3120
rect 19524 3136 19576 3188
rect 20076 3136 20128 3188
rect 21640 3136 21692 3188
rect 22192 3136 22244 3188
rect 24400 3179 24452 3188
rect 24400 3145 24409 3179
rect 24409 3145 24443 3179
rect 24443 3145 24452 3179
rect 24400 3136 24452 3145
rect 14464 3000 14516 3052
rect 11336 2932 11388 2984
rect 12532 2932 12584 2984
rect 15016 3043 15068 3052
rect 15016 3009 15025 3043
rect 15025 3009 15059 3043
rect 15059 3009 15068 3043
rect 15936 3043 15988 3052
rect 15016 3000 15068 3009
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 17224 3000 17276 3052
rect 17592 3043 17644 3052
rect 17592 3009 17601 3043
rect 17601 3009 17635 3043
rect 17635 3009 17644 3043
rect 17592 3000 17644 3009
rect 18328 3000 18380 3052
rect 18972 3068 19024 3120
rect 22560 3068 22612 3120
rect 23112 3111 23164 3120
rect 23112 3077 23121 3111
rect 23121 3077 23155 3111
rect 23155 3077 23164 3111
rect 23112 3068 23164 3077
rect 16764 2932 16816 2984
rect 17776 2932 17828 2984
rect 19340 3000 19392 3052
rect 19524 3043 19576 3052
rect 19524 3009 19533 3043
rect 19533 3009 19567 3043
rect 19567 3009 19576 3043
rect 19524 3000 19576 3009
rect 19984 3000 20036 3052
rect 20444 3000 20496 3052
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 22376 3043 22428 3052
rect 20260 2932 20312 2984
rect 20720 2932 20772 2984
rect 21824 2932 21876 2984
rect 22376 3009 22385 3043
rect 22385 3009 22419 3043
rect 22419 3009 22428 3043
rect 22376 3000 22428 3009
rect 23020 3043 23072 3052
rect 23020 3009 23039 3043
rect 23039 3009 23072 3043
rect 23020 3000 23072 3009
rect 23296 3000 23348 3052
rect 29000 3179 29052 3188
rect 29000 3145 29009 3179
rect 29009 3145 29043 3179
rect 29043 3145 29052 3179
rect 29000 3136 29052 3145
rect 31208 3179 31260 3188
rect 31208 3145 31217 3179
rect 31217 3145 31251 3179
rect 31251 3145 31260 3179
rect 31208 3136 31260 3145
rect 33324 3179 33376 3188
rect 33324 3145 33333 3179
rect 33333 3145 33367 3179
rect 33367 3145 33376 3179
rect 33324 3136 33376 3145
rect 27528 3068 27580 3120
rect 34520 3136 34572 3188
rect 24216 3043 24268 3052
rect 24216 3009 24225 3043
rect 24225 3009 24259 3043
rect 24259 3009 24268 3043
rect 25136 3043 25188 3052
rect 24216 3000 24268 3009
rect 25136 3009 25145 3043
rect 25145 3009 25179 3043
rect 25179 3009 25188 3043
rect 25136 3000 25188 3009
rect 25596 3043 25648 3052
rect 25596 3009 25605 3043
rect 25605 3009 25639 3043
rect 25639 3009 25648 3043
rect 25596 3000 25648 3009
rect 27068 3000 27120 3052
rect 27160 3000 27212 3052
rect 27896 3043 27948 3052
rect 27896 3009 27905 3043
rect 27905 3009 27939 3043
rect 27939 3009 27948 3043
rect 27896 3000 27948 3009
rect 28264 3000 28316 3052
rect 28540 3043 28592 3052
rect 28540 3009 28549 3043
rect 28549 3009 28583 3043
rect 28583 3009 28592 3043
rect 28540 3000 28592 3009
rect 30472 3000 30524 3052
rect 30748 3043 30800 3052
rect 30748 3009 30757 3043
rect 30757 3009 30791 3043
rect 30791 3009 30800 3043
rect 30748 3000 30800 3009
rect 31024 3000 31076 3052
rect 31392 3043 31444 3052
rect 31392 3009 31401 3043
rect 31401 3009 31435 3043
rect 31435 3009 31444 3043
rect 31392 3000 31444 3009
rect 33232 3000 33284 3052
rect 34336 3000 34388 3052
rect 35992 3000 36044 3052
rect 37096 3000 37148 3052
rect 11888 2864 11940 2916
rect 7380 2796 7432 2848
rect 9680 2796 9732 2848
rect 13544 2796 13596 2848
rect 13728 2796 13780 2848
rect 14832 2796 14884 2848
rect 16028 2864 16080 2916
rect 16120 2864 16172 2916
rect 15016 2796 15068 2848
rect 18880 2796 18932 2848
rect 19432 2864 19484 2916
rect 22284 2864 22336 2916
rect 23112 2932 23164 2984
rect 21456 2796 21508 2848
rect 22192 2796 22244 2848
rect 22560 2796 22612 2848
rect 23296 2864 23348 2916
rect 25228 2864 25280 2916
rect 26056 2864 26108 2916
rect 28632 2864 28684 2916
rect 33140 2864 33192 2916
rect 22836 2796 22888 2848
rect 23848 2796 23900 2848
rect 25044 2796 25096 2848
rect 26332 2796 26384 2848
rect 31484 2796 31536 2848
rect 32680 2839 32732 2848
rect 32680 2805 32689 2839
rect 32689 2805 32723 2839
rect 32723 2805 32732 2839
rect 32680 2796 32732 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4712 2524 4764 2576
rect 5816 2567 5868 2576
rect 5816 2533 5825 2567
rect 5825 2533 5859 2567
rect 5859 2533 5868 2567
rect 5816 2524 5868 2533
rect 2320 2388 2372 2440
rect 7012 2456 7064 2508
rect 5448 2388 5500 2440
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 6184 2388 6236 2440
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7288 2388 7340 2440
rect 7840 2388 7892 2440
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 8944 2388 8996 2440
rect 10048 2456 10100 2508
rect 13728 2524 13780 2576
rect 15200 2524 15252 2576
rect 16304 2524 16356 2576
rect 9680 2388 9732 2440
rect 10600 2388 10652 2440
rect 10968 2388 11020 2440
rect 12256 2388 12308 2440
rect 12808 2388 12860 2440
rect 12900 2388 12952 2440
rect 13728 2388 13780 2440
rect 14096 2388 14148 2440
rect 15016 2388 15068 2440
rect 15752 2456 15804 2508
rect 20260 2592 20312 2644
rect 25228 2635 25280 2644
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 20628 2524 20680 2576
rect 21640 2524 21692 2576
rect 18328 2456 18380 2508
rect 3424 2252 3476 2304
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 9588 2252 9640 2304
rect 12348 2252 12400 2304
rect 14924 2320 14976 2372
rect 16856 2388 16908 2440
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 17684 2431 17736 2440
rect 16948 2388 17000 2397
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 18236 2388 18288 2440
rect 22100 2456 22152 2508
rect 20260 2388 20312 2440
rect 20904 2388 20956 2440
rect 22284 2388 22336 2440
rect 23480 2388 23532 2440
rect 24584 2456 24636 2508
rect 25964 2567 26016 2576
rect 25964 2533 25973 2567
rect 25973 2533 26007 2567
rect 26007 2533 26016 2567
rect 25964 2524 26016 2533
rect 26608 2524 26660 2576
rect 15292 2320 15344 2372
rect 15568 2320 15620 2372
rect 16580 2320 16632 2372
rect 17224 2320 17276 2372
rect 22744 2320 22796 2372
rect 15108 2252 15160 2304
rect 15200 2252 15252 2304
rect 16212 2252 16264 2304
rect 17776 2252 17828 2304
rect 18328 2252 18380 2304
rect 18880 2252 18932 2304
rect 19984 2295 20036 2304
rect 19984 2261 19993 2295
rect 19993 2261 20027 2295
rect 20027 2261 20036 2295
rect 19984 2252 20036 2261
rect 20536 2252 20588 2304
rect 21088 2252 21140 2304
rect 22192 2252 22244 2304
rect 24860 2388 24912 2440
rect 26516 2456 26568 2508
rect 28816 2524 28868 2576
rect 26240 2388 26292 2440
rect 25504 2320 25556 2372
rect 26884 2320 26936 2372
rect 27620 2388 27672 2440
rect 28632 2431 28684 2440
rect 28632 2397 28641 2431
rect 28641 2397 28675 2431
rect 28675 2397 28684 2431
rect 28632 2388 28684 2397
rect 27712 2320 27764 2372
rect 29920 2456 29972 2508
rect 29000 2388 29052 2440
rect 29552 2388 29604 2440
rect 31484 2456 31536 2508
rect 37648 2456 37700 2508
rect 38016 2456 38068 2508
rect 29092 2320 29144 2372
rect 29368 2320 29420 2372
rect 31760 2388 31812 2440
rect 32680 2388 32732 2440
rect 32220 2320 32272 2372
rect 33140 2388 33192 2440
rect 33692 2388 33744 2440
rect 33784 2388 33836 2440
rect 34704 2388 34756 2440
rect 34980 2388 35032 2440
rect 35900 2388 35952 2440
rect 37832 2431 37884 2440
rect 37832 2397 37841 2431
rect 37841 2397 37875 2431
rect 37875 2397 37884 2431
rect 37832 2388 37884 2397
rect 27068 2295 27120 2304
rect 27068 2261 27077 2295
rect 27077 2261 27111 2295
rect 27111 2261 27120 2295
rect 29552 2295 29604 2304
rect 27068 2252 27120 2261
rect 29552 2261 29561 2295
rect 29561 2261 29595 2295
rect 29595 2261 29604 2295
rect 29552 2252 29604 2261
rect 30196 2295 30248 2304
rect 30196 2261 30205 2295
rect 30205 2261 30239 2295
rect 30239 2261 30248 2295
rect 30196 2252 30248 2261
rect 32128 2295 32180 2304
rect 32128 2261 32137 2295
rect 32137 2261 32171 2295
rect 32171 2261 32180 2295
rect 32128 2252 32180 2261
rect 32772 2295 32824 2304
rect 32772 2261 32781 2295
rect 32781 2261 32815 2295
rect 32815 2261 32824 2295
rect 32772 2252 32824 2261
rect 33416 2295 33468 2304
rect 33416 2261 33425 2295
rect 33425 2261 33459 2295
rect 33459 2261 33468 2295
rect 33416 2252 33468 2261
rect 34520 2252 34572 2304
rect 34796 2252 34848 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 5172 2048 5224 2100
rect 21916 2048 21968 2100
rect 23572 2048 23624 2100
rect 29552 2048 29604 2100
rect 7104 1980 7156 2032
rect 22008 1980 22060 2032
rect 23112 1980 23164 2032
rect 32128 1980 32180 2032
rect 10416 1912 10468 1964
rect 20352 1912 20404 1964
rect 33416 1912 33468 1964
rect 24492 1844 24544 1896
rect 30196 1844 30248 1896
rect 22468 1776 22520 1828
rect 32772 1776 32824 1828
rect 24860 1708 24912 1760
rect 22652 1640 22704 1692
rect 34796 1640 34848 1692
rect 24400 1368 24452 1420
rect 25964 1368 26016 1420
<< metal2 >>
rect 662 39200 718 40000
rect 1766 39200 1822 40000
rect 2870 39200 2926 40000
rect 3974 39200 4030 40000
rect 5078 39200 5134 40000
rect 6182 39200 6238 40000
rect 7286 39200 7342 40000
rect 8390 39200 8446 40000
rect 9494 39200 9550 40000
rect 10598 39200 10654 40000
rect 11702 39200 11758 40000
rect 12806 39200 12862 40000
rect 13910 39200 13966 40000
rect 15014 39200 15070 40000
rect 16118 39200 16174 40000
rect 17222 39200 17278 40000
rect 18326 39200 18382 40000
rect 19430 39200 19486 40000
rect 20534 39200 20590 40000
rect 21638 39200 21694 40000
rect 22742 39200 22798 40000
rect 23846 39200 23902 40000
rect 24950 39200 25006 40000
rect 26054 39200 26110 40000
rect 27158 39200 27214 40000
rect 28262 39200 28318 40000
rect 29366 39200 29422 40000
rect 30470 39200 30526 40000
rect 31574 39200 31630 40000
rect 32678 39200 32734 40000
rect 33782 39200 33838 40000
rect 34886 39200 34942 40000
rect 35990 39200 36046 40000
rect 37094 39200 37150 40000
rect 38198 39200 38254 40000
rect 39302 39200 39358 40000
rect 676 37262 704 39200
rect 664 37256 716 37262
rect 664 37198 716 37204
rect 1308 37256 1360 37262
rect 1308 37198 1360 37204
rect 1320 36378 1348 37198
rect 1780 36922 1808 39200
rect 2884 37262 2912 39200
rect 3988 37262 4016 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5092 37262 5120 39200
rect 6196 37262 6224 39200
rect 7300 37262 7328 39200
rect 8404 37466 8432 39200
rect 8392 37460 8444 37466
rect 8392 37402 8444 37408
rect 8404 37262 8432 37402
rect 9508 37262 9536 39200
rect 10612 37262 10640 39200
rect 11716 37262 11744 39200
rect 12820 37262 12848 39200
rect 13924 37262 13952 39200
rect 15028 37262 15056 39200
rect 16132 37466 16160 39200
rect 16120 37460 16172 37466
rect 16120 37402 16172 37408
rect 17236 37262 17264 39200
rect 18340 37262 18368 39200
rect 19444 37262 19472 39200
rect 20548 37262 20576 39200
rect 2872 37256 2924 37262
rect 2872 37198 2924 37204
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 6184 37256 6236 37262
rect 6184 37198 6236 37204
rect 7288 37256 7340 37262
rect 7288 37198 7340 37204
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 9496 37256 9548 37262
rect 9496 37198 9548 37204
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 12808 37256 12860 37262
rect 12808 37198 12860 37204
rect 13912 37256 13964 37262
rect 13912 37198 13964 37204
rect 15016 37256 15068 37262
rect 15016 37198 15068 37204
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 18328 37256 18380 37262
rect 19432 37256 19484 37262
rect 18328 37198 18380 37204
rect 19352 37204 19432 37210
rect 19352 37198 19484 37204
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 1952 37120 2004 37126
rect 1952 37062 2004 37068
rect 1768 36916 1820 36922
rect 1768 36858 1820 36864
rect 1308 36372 1360 36378
rect 1308 36314 1360 36320
rect 1584 30252 1636 30258
rect 1584 30194 1636 30200
rect 1596 30025 1624 30194
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1596 29850 1624 29951
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1964 4826 1992 37062
rect 2884 36922 2912 37198
rect 3148 37120 3200 37126
rect 3148 37062 3200 37068
rect 2872 36916 2924 36922
rect 2872 36858 2924 36864
rect 2412 36780 2464 36786
rect 2412 36722 2464 36728
rect 2424 36038 2452 36722
rect 2412 36032 2464 36038
rect 2412 35974 2464 35980
rect 2044 30116 2096 30122
rect 2044 30058 2096 30064
rect 2056 7954 2084 30058
rect 2424 14074 2452 35974
rect 3160 22098 3188 37062
rect 3988 36922 4016 37198
rect 4620 37188 4672 37194
rect 4620 37130 4672 37136
rect 3976 36916 4028 36922
rect 3976 36858 4028 36864
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2608 16250 2636 18022
rect 2976 17678 3004 19450
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2792 15434 2820 15846
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 2792 15162 2820 15370
rect 2884 15366 2912 17478
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 3252 15026 3280 18022
rect 3344 15366 3372 19110
rect 4080 18902 4108 19246
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 3700 18692 3752 18698
rect 3700 18634 3752 18640
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 18290 3464 18566
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3712 16574 3740 18634
rect 4632 18426 4660 37130
rect 4712 37120 4764 37126
rect 4712 37062 4764 37068
rect 4724 20058 4752 37062
rect 5092 36922 5120 37198
rect 6196 36922 6224 37198
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 5080 36916 5132 36922
rect 5080 36858 5132 36864
rect 6184 36916 6236 36922
rect 6184 36858 6236 36864
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4724 19514 4752 19994
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 6380 19310 6408 37062
rect 7300 36922 7328 37198
rect 7380 37120 7432 37126
rect 7380 37062 7432 37068
rect 8944 37120 8996 37126
rect 8944 37062 8996 37068
rect 7288 36916 7340 36922
rect 7288 36858 7340 36864
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 5552 18766 5580 19246
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5920 18698 5948 18770
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5908 18692 5960 18698
rect 5908 18634 5960 18640
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3804 17338 3832 18158
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18362
rect 5184 18086 5212 18634
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3804 17218 3832 17274
rect 3804 17190 4016 17218
rect 3712 16546 3924 16574
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2424 12322 2452 14010
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2424 12294 2544 12322
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2424 9178 2452 12106
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2516 9110 2544 12294
rect 2884 12238 2912 12854
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 11762 2912 12174
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2884 11150 2912 11698
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 2608 7546 2636 8910
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2700 6458 2728 11018
rect 2884 10810 2912 11086
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2884 10062 2912 10746
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2976 9450 3004 12786
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2792 8566 2820 8910
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2884 8634 2912 8842
rect 3068 8634 3096 9522
rect 3160 9042 3188 12582
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3252 8974 3280 12038
rect 3240 8968 3292 8974
rect 3160 8916 3240 8922
rect 3160 8910 3292 8916
rect 3160 8894 3280 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2792 7886 2820 8502
rect 3160 7886 3188 8894
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8566 3280 8774
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3252 8022 3280 8366
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2792 6186 2820 6734
rect 2884 6730 2912 7414
rect 3160 7410 3188 7822
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6798 3096 7278
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2884 6322 2912 6666
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6322 3188 6598
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2884 3194 2912 6258
rect 3344 5302 3372 15302
rect 3804 15094 3832 15438
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3804 14482 3832 15030
rect 3896 14822 3924 16546
rect 3988 15910 4016 17190
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 14618 3924 14758
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3804 13938 3832 14418
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3436 10033 3464 10746
rect 3422 10024 3478 10033
rect 3422 9959 3478 9968
rect 3620 8498 3648 11222
rect 3988 10674 4016 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15502 4660 17478
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 5184 15366 5212 18022
rect 5368 17678 5396 18566
rect 5920 18222 5948 18634
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5920 16658 5948 18158
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4448 14006 4476 14214
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 5184 11898 5212 15302
rect 5552 14498 5580 16526
rect 5644 16266 5672 16594
rect 5644 16238 5764 16266
rect 5552 14470 5672 14498
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 3804 9178 3832 9930
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 4632 9042 4660 9862
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4172 8498 4200 8910
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3528 8090 3556 8434
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3620 7886 3648 8434
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3620 7002 3648 7822
rect 3804 7546 3832 8434
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 8978
rect 4724 8634 4752 11698
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4816 8514 4844 11494
rect 5276 10742 5304 13194
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5552 9178 5580 14282
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 4988 8560 5040 8566
rect 4816 8508 4988 8514
rect 4816 8502 5040 8508
rect 4816 8486 5028 8502
rect 5080 8492 5132 8498
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 4448 7410 4476 7822
rect 4632 7410 4660 7890
rect 4816 7886 4844 8486
rect 5080 8434 5132 8440
rect 5092 8090 5120 8434
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 5184 7546 5212 8842
rect 5644 8634 5672 14470
rect 5736 14346 5764 16238
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6196 15502 6224 15982
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 6196 14958 6224 15438
rect 6564 15162 6592 17478
rect 6656 16182 6684 18022
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6748 15502 6776 18022
rect 7116 17678 7144 18566
rect 7300 18290 7328 19110
rect 7392 18970 7420 37062
rect 8956 26234 8984 37062
rect 9508 36922 9536 37198
rect 10324 37188 10376 37194
rect 10324 37130 10376 37136
rect 9588 37120 9640 37126
rect 9588 37062 9640 37068
rect 9496 36916 9548 36922
rect 9496 36858 9548 36864
rect 8864 26206 8984 26234
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7576 16574 7604 22034
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 19378 7696 19654
rect 8312 19514 8340 19994
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18170 7696 19314
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7944 18834 7972 19178
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7760 18358 7788 18566
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 7668 18142 7788 18170
rect 7576 16546 7696 16574
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6196 14414 6224 14894
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 6748 13190 6776 14758
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 14074 6868 14214
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12918 6776 13126
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7116 12238 7144 12718
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7116 11830 7144 12174
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7116 11150 7144 11766
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6012 8634 6040 8774
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 5276 7342 5304 8026
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5552 7002 5580 7142
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6225 3832 6598
rect 3790 6216 3846 6225
rect 4356 6186 4384 6870
rect 5644 6798 5672 8570
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5920 8090 5948 8298
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 6104 7886 6132 8366
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7342 5764 7686
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 3790 6151 3846 6160
rect 4344 6180 4396 6186
rect 3804 6118 3832 6151
rect 4344 6122 4396 6128
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3988 3058 4016 3334
rect 4632 3058 4660 3334
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2332 800 2360 2382
rect 2884 800 2912 2994
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 800 3464 2246
rect 3988 800 4016 2994
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2530 4660 2994
rect 4724 2582 4752 6122
rect 5736 5914 5764 7278
rect 6104 7018 6132 7822
rect 6196 7410 6224 7822
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6104 6990 6224 7018
rect 6196 6934 6224 6990
rect 6184 6928 6236 6934
rect 6288 6914 6316 11018
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6656 7886 6684 8910
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6656 7546 6684 7822
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6288 6886 6408 6914
rect 6184 6870 6236 6876
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 6380 5370 6408 6886
rect 6748 6662 6776 8366
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 8090 6960 8230
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7342 6868 7822
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 6866 6868 7278
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6840 6746 6868 6802
rect 6840 6730 6960 6746
rect 6840 6724 6972 6730
rect 6840 6718 6920 6724
rect 6920 6666 6972 6672
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6564 4282 6592 5170
rect 6748 5166 6776 6598
rect 7300 5370 7328 12106
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6748 4690 6776 5102
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6932 4282 6960 4694
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 5092 3058 5120 3334
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 4540 2502 4660 2530
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4540 800 4568 2502
rect 5092 800 5120 2994
rect 5460 2446 5488 3878
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5644 2446 5672 3334
rect 6748 3058 6776 3470
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 5816 2576 5868 2582
rect 5814 2544 5816 2553
rect 5868 2544 5870 2553
rect 5814 2479 5870 2488
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 2106 5212 2246
rect 5460 2122 5488 2382
rect 5172 2100 5224 2106
rect 5460 2094 5672 2122
rect 5172 2042 5224 2048
rect 5644 800 5672 2094
rect 6196 800 6224 2382
rect 6748 800 6776 2994
rect 6932 2446 6960 3334
rect 7024 2514 7052 4422
rect 7116 4078 7144 5034
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 4146 7236 4422
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7300 3194 7328 4694
rect 7392 4554 7420 11290
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7484 8090 7512 8434
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7668 5370 7696 16546
rect 7760 15910 7788 18142
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 11665 7788 15846
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 12442 8156 15302
rect 8220 14804 8248 18294
rect 8312 17882 8340 18702
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8404 15366 8432 18362
rect 8496 18290 8524 19110
rect 8864 18766 8892 26206
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8956 18426 8984 19246
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 16114 8984 16526
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8956 15570 8984 16050
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8300 14816 8352 14822
rect 8220 14776 8300 14804
rect 8300 14758 8352 14764
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7746 11656 7802 11665
rect 7746 11591 7802 11600
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7760 7410 7788 11494
rect 7852 8634 7880 11698
rect 8220 10810 8248 13806
rect 8312 10810 8340 14758
rect 9232 12918 9260 18566
rect 9324 16182 9352 18838
rect 9416 16522 9444 20198
rect 9600 20058 9628 37062
rect 10336 20602 10364 37130
rect 10612 36922 10640 37198
rect 10692 37120 10744 37126
rect 10692 37062 10744 37068
rect 11520 37120 11572 37126
rect 11520 37062 11572 37068
rect 10600 36916 10652 36922
rect 10600 36858 10652 36864
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9312 16176 9364 16182
rect 9312 16118 9364 16124
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9324 15026 9352 15506
rect 9508 15162 9536 18906
rect 9692 18834 9720 19314
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 15434 9628 18634
rect 9968 18290 9996 19654
rect 10244 19514 10272 20402
rect 10336 19854 10364 20538
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10612 19922 10640 20198
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9324 14414 9352 14962
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 10152 14346 10180 18022
rect 10336 16454 10364 18022
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10336 13462 10364 16390
rect 10428 14278 10456 19654
rect 10612 19242 10640 19858
rect 10704 19446 10732 37062
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11440 19786 11468 20810
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10704 18086 10732 19246
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18766 11100 19110
rect 11164 18902 11192 19654
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 10428 13258 10456 13670
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8772 9450 8800 11018
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8864 9178 8892 12786
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8956 8634 8984 9522
rect 9968 9042 9996 12582
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 11762 10088 12174
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 11218 10088 11698
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10742 10088 11154
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10152 9926 10180 10610
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7852 7546 7880 8366
rect 9140 8362 9168 8502
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8220 7478 8248 7958
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8036 6914 8064 7346
rect 8036 6886 8156 6914
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7852 6254 7880 6734
rect 8024 6724 8076 6730
rect 8024 6666 8076 6672
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7852 5710 7880 6190
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7668 5166 7696 5306
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7852 5098 7880 5646
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7944 4978 7972 5714
rect 8036 5710 8064 6666
rect 8128 5794 8156 6886
rect 8220 6458 8248 7414
rect 8956 6866 8984 8298
rect 9140 7546 9168 8298
rect 9968 8294 9996 8978
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9048 5914 9076 6258
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 8128 5766 8248 5794
rect 8220 5710 8248 5766
rect 9324 5710 9352 6802
rect 9416 5778 9444 7482
rect 9692 7478 9720 7686
rect 9968 7478 9996 8026
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 6118 9536 7278
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5234 8340 5510
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7852 4950 7972 4978
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7852 4622 7880 4950
rect 9508 4622 9536 6054
rect 9600 5642 9628 6666
rect 9968 6390 9996 7414
rect 10152 6798 10180 7754
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 7378 4176 7434 4185
rect 7378 4111 7434 4120
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7392 2854 7420 4111
rect 9600 4078 9628 5578
rect 10152 4826 10180 6734
rect 10244 5710 10272 12038
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10336 9058 10364 11290
rect 10428 10062 10456 13194
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10336 9030 10456 9058
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10336 8362 10364 8910
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10428 7818 10456 9030
rect 10520 8974 10548 14010
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10520 8090 10548 8910
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10520 7886 10548 8026
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10520 6458 10548 7346
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10612 6202 10640 14214
rect 11440 13326 11468 19722
rect 11532 19514 11560 37062
rect 11716 36922 11744 37198
rect 12820 36922 12848 37198
rect 13924 36922 13952 37198
rect 14096 37120 14148 37126
rect 14096 37062 14148 37068
rect 11704 36916 11756 36922
rect 11704 36858 11756 36864
rect 12808 36916 12860 36922
rect 12808 36858 12860 36864
rect 13912 36916 13964 36922
rect 13912 36858 13964 36864
rect 14108 26234 14136 37062
rect 15028 36922 15056 37198
rect 15844 37188 15896 37194
rect 15844 37130 15896 37136
rect 15108 37120 15160 37126
rect 15108 37062 15160 37068
rect 15016 36916 15068 36922
rect 15016 36858 15068 36864
rect 13924 26206 14136 26234
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 12268 20466 12296 20742
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 19922 12296 20402
rect 13372 20398 13400 20742
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11716 19242 11744 19858
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11716 18086 11744 19178
rect 11808 18766 11836 19654
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11992 18086 12020 19246
rect 12728 18970 12756 19314
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11072 12986 11100 13262
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10796 9450 10824 11018
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10428 6174 10640 6202
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10244 5030 10272 5646
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 9692 4214 9720 4762
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7852 2446 7880 3402
rect 8220 2446 8248 3878
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8404 3058 8432 3538
rect 9508 3058 9536 3946
rect 9692 3738 9720 4150
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9692 3534 9720 3674
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 2038 7144 2246
rect 7104 2032 7156 2038
rect 7104 1974 7156 1980
rect 7300 800 7328 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 2009 7788 2246
rect 7746 2000 7802 2009
rect 7746 1935 7802 1944
rect 7852 800 7880 2382
rect 8404 800 8432 2994
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8956 800 8984 2382
rect 9508 800 9536 2994
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9692 2446 9720 2790
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9588 2304 9640 2310
rect 9588 2246 9640 2252
rect 9600 1873 9628 2246
rect 9586 1864 9642 1873
rect 9586 1799 9642 1808
rect 10060 800 10088 2450
rect 10428 1970 10456 6174
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5778 10640 6054
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10704 4690 10732 7754
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10520 3194 10548 4558
rect 10704 4146 10732 4626
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10612 3602 10640 3946
rect 10796 3942 10824 6394
rect 10888 5642 10916 10542
rect 10980 10266 11008 10610
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 8634 11008 9522
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11072 7954 11100 10406
rect 11348 9178 11376 12106
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11072 6866 11100 7890
rect 11440 7886 11468 8502
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11072 6254 11100 6802
rect 11256 6322 11284 7686
rect 11532 7546 11560 18022
rect 11992 15910 12020 18022
rect 12532 16516 12584 16522
rect 12532 16458 12584 16464
rect 12544 16046 12572 16458
rect 12820 16182 12848 19450
rect 12912 18834 12940 20198
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 8634 11744 11494
rect 11992 9382 12020 15846
rect 12544 15434 12572 15982
rect 13372 15706 13400 20334
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 19292 13768 19654
rect 13832 19446 13860 19722
rect 13820 19440 13872 19446
rect 13820 19382 13872 19388
rect 13924 19378 13952 26206
rect 15120 19446 15148 37062
rect 15856 20058 15884 37130
rect 16764 37120 16816 37126
rect 16764 37062 16816 37068
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 16316 19718 16344 20334
rect 16592 19786 16620 20742
rect 16776 20602 16804 37062
rect 17236 36922 17264 37198
rect 18340 36922 18368 37198
rect 19352 37182 19472 37198
rect 18420 37120 18472 37126
rect 18420 37062 18472 37068
rect 17224 36916 17276 36922
rect 17224 36858 17276 36864
rect 18328 36916 18380 36922
rect 18328 36858 18380 36864
rect 18432 20602 18460 37062
rect 19352 36922 19380 37182
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19340 36916 19392 36922
rect 19340 36858 19392 36864
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 18420 20596 18472 20602
rect 18420 20538 18472 20544
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16684 19854 16712 20198
rect 17420 19922 17448 20266
rect 19444 20058 19472 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20548 36922 20576 37198
rect 21652 37126 21680 39200
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 20628 37120 20680 37126
rect 20628 37062 20680 37068
rect 21640 37120 21692 37126
rect 21640 37062 21692 37068
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 19984 36576 20036 36582
rect 19984 36518 20036 36524
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 15108 19440 15160 19446
rect 15108 19382 15160 19388
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13740 19264 13860 19292
rect 13832 19174 13860 19264
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13740 16590 13768 17070
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 14958 12572 15370
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12544 14482 12572 14894
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12544 13394 12572 14418
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11716 7698 11744 8570
rect 11808 8090 11836 8842
rect 12084 8498 12112 12038
rect 13372 9042 13400 15642
rect 13556 13258 13584 16390
rect 13740 16046 13768 16526
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13740 15502 13768 15982
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13832 15144 13860 19110
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 13648 15116 13860 15144
rect 13648 14822 13676 15116
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13648 13734 13676 14758
rect 13740 14482 13768 14894
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13740 13938 13768 14418
rect 13924 14346 13952 14758
rect 14108 14618 14136 15370
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 14016 13462 14044 14554
rect 14384 14414 14412 18566
rect 15212 16590 15240 19654
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 15672 16454 15700 19654
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 15028 14822 15056 15302
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 15120 13530 15148 14962
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14521 15792 14758
rect 16224 14618 16252 15370
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 15750 14512 15806 14521
rect 15750 14447 15806 14456
rect 16488 14272 16540 14278
rect 16592 14260 16620 19722
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16868 18766 16896 19654
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17420 19292 17448 19858
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 17500 19304 17552 19310
rect 17420 19264 17500 19292
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 17328 18086 17356 19246
rect 17420 18970 17448 19264
rect 17500 19246 17552 19252
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17880 16250 17908 18022
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17512 14958 17540 15302
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 16540 14232 16620 14260
rect 16488 14214 16540 14220
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14292 12238 14320 12718
rect 15580 12442 15608 12786
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11716 7670 11928 7698
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11900 7342 11928 7670
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11794 7032 11850 7041
rect 11794 6967 11796 6976
rect 11848 6967 11850 6976
rect 11796 6938 11848 6944
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 6322 11744 6666
rect 11808 6458 11836 6802
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11808 6322 11836 6394
rect 11900 6390 11928 7278
rect 11992 6866 12020 8230
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12084 6730 12112 8434
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11992 6458 12020 6598
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11256 5642 11284 6258
rect 11808 6118 11836 6258
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11440 5710 11468 6054
rect 11992 5778 12020 6258
rect 12176 6254 12204 6938
rect 12360 6662 12388 8910
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 12714 6760 12770 6769
rect 12714 6695 12770 6704
rect 12728 6662 12756 6695
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12176 5778 12204 6190
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11072 4078 11100 4490
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10612 3058 10640 3538
rect 10796 3534 10824 3878
rect 11256 3534 11284 3878
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11610 3496 11666 3505
rect 11256 3058 11284 3470
rect 11610 3431 11666 3440
rect 11624 3126 11652 3431
rect 11612 3120 11664 3126
rect 11334 3088 11390 3097
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 11244 3052 11296 3058
rect 11612 3062 11664 3068
rect 11716 3058 11744 4422
rect 11900 4078 11928 4490
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11808 3602 11836 4014
rect 11900 3942 11928 4014
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3738 11928 3878
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11992 3534 12020 5714
rect 12268 5710 12296 6326
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12636 5914 12664 6258
rect 12820 6186 12848 6870
rect 13188 6644 13216 7822
rect 13740 7410 13768 11222
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13280 6769 13308 7142
rect 13740 7002 13768 7346
rect 13832 7206 13860 7890
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13266 6760 13322 6769
rect 13266 6695 13322 6704
rect 13268 6656 13320 6662
rect 13188 6616 13268 6644
rect 13268 6598 13320 6604
rect 13280 6254 13308 6598
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12452 5778 12480 5850
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12268 4282 12296 5646
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 13280 4146 13308 6190
rect 13832 6118 13860 7142
rect 13924 6322 13952 7822
rect 14016 6322 14044 11766
rect 14292 11694 14320 12174
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14292 11150 14320 11630
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 10606 14320 11086
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14292 10130 14320 10542
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14292 9586 14320 10066
rect 15764 10062 15792 10406
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15488 9178 15516 9318
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14108 8090 14136 9046
rect 15580 8634 15608 9522
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14936 8022 14964 8366
rect 14924 8016 14976 8022
rect 14924 7958 14976 7964
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14936 7546 14964 7754
rect 15764 7546 15792 8434
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15844 7472 15896 7478
rect 15844 7414 15896 7420
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14108 7041 14136 7278
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14094 7032 14150 7041
rect 14094 6967 14150 6976
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13648 5914 13676 6054
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13924 5574 13952 6258
rect 14108 5710 14136 6734
rect 14200 6662 14228 7142
rect 14568 7002 14596 7346
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14292 6662 14320 6938
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14384 6390 14412 6802
rect 14568 6798 14596 6938
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14660 6254 14688 7142
rect 15028 7002 15056 7210
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 15212 6746 15240 7346
rect 15856 7002 15884 7414
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 16132 6798 16160 8026
rect 15292 6792 15344 6798
rect 15212 6740 15292 6746
rect 15212 6734 15344 6740
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 15212 6718 15332 6734
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 15028 5914 15056 6326
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 15120 4758 15148 6122
rect 15212 5778 15240 6718
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11334 3023 11390 3032
rect 11704 3052 11756 3058
rect 11244 2994 11296 3000
rect 11348 2990 11376 3023
rect 11704 2994 11756 3000
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10968 2440 11020 2446
rect 11020 2400 11192 2428
rect 10968 2382 11020 2388
rect 10416 1964 10468 1970
rect 10416 1906 10468 1912
rect 10612 800 10640 2382
rect 11164 800 11192 2400
rect 11716 800 11744 2994
rect 11886 2952 11942 2961
rect 11886 2887 11888 2896
rect 11940 2887 11942 2896
rect 11888 2858 11940 2864
rect 12268 2446 12296 3946
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13542 3360 13598 3369
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12544 2666 12572 2926
rect 12360 2638 12572 2666
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12268 800 12296 2382
rect 12360 2310 12388 2638
rect 12912 2446 12940 3334
rect 13464 3058 13492 3334
rect 13542 3295 13598 3304
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13464 2774 13492 2994
rect 13556 2854 13584 3295
rect 13648 3194 13676 3402
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13372 2746 13492 2774
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12820 800 12848 2382
rect 13372 800 13400 2746
rect 13740 2582 13768 2790
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 14108 2446 14136 3878
rect 15120 3534 15148 4558
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 13728 2440 13780 2446
rect 14096 2440 14148 2446
rect 13780 2400 13952 2428
rect 13728 2382 13780 2388
rect 13924 800 13952 2400
rect 14096 2382 14148 2388
rect 14476 800 14504 2994
rect 15028 2938 15056 2994
rect 14844 2910 15056 2938
rect 14844 2854 14872 2910
rect 15028 2854 15056 2910
rect 14832 2848 14884 2854
rect 15016 2848 15068 2854
rect 14832 2790 14884 2796
rect 14922 2816 14978 2825
rect 15016 2790 15068 2796
rect 14922 2751 14978 2760
rect 14936 2378 14964 2751
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 15028 800 15056 2382
rect 15120 2310 15148 3470
rect 15212 3194 15240 4082
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15212 2310 15240 2518
rect 15304 2378 15332 3946
rect 15396 3738 15424 5102
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15672 4146 15700 4422
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15672 4049 15700 4082
rect 15658 4040 15714 4049
rect 15568 4004 15620 4010
rect 15658 3975 15714 3984
rect 15568 3946 15620 3952
rect 15580 3738 15608 3946
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15396 2825 15424 3674
rect 15764 3670 15792 4082
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 15382 2816 15438 2825
rect 15382 2751 15438 2760
rect 15764 2514 15792 3606
rect 15856 3602 15884 4626
rect 16120 3936 16172 3942
rect 16224 3913 16252 11834
rect 16316 3942 16344 12310
rect 16500 8974 16528 14214
rect 17696 14074 17724 15370
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17236 12986 17264 13262
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17880 11898 17908 16186
rect 18064 15162 18092 17138
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 19260 15450 19288 16458
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19352 15638 19380 16390
rect 19444 15978 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19996 15502 20024 36518
rect 20640 19514 20668 37062
rect 21836 36582 21864 37198
rect 22756 37126 22784 39200
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 22744 37120 22796 37126
rect 22744 37062 22796 37068
rect 23032 36582 23060 37198
rect 23860 37126 23888 39200
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 23848 37120 23900 37126
rect 23848 37062 23900 37068
rect 21824 36576 21876 36582
rect 21824 36518 21876 36524
rect 23020 36576 23072 36582
rect 23020 36518 23072 36524
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 19984 15496 20036 15502
rect 19260 15422 19472 15450
rect 19984 15438 20036 15444
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18708 14414 18736 15302
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19168 14618 19196 14962
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 19260 13938 19288 14758
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19352 14006 19380 14214
rect 19444 14074 19472 15422
rect 20260 15428 20312 15434
rect 20260 15370 20312 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13462 19564 13670
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19524 13456 19576 13462
rect 19524 13398 19576 13404
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18800 11898 18828 12106
rect 19352 11898 19380 12582
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17880 10266 17908 11698
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18248 11082 18276 11494
rect 18340 11286 18368 11494
rect 18328 11280 18380 11286
rect 18328 11222 18380 11228
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18144 11076 18196 11082
rect 18144 11018 18196 11024
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10674 18000 10950
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9722 18000 9998
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 17328 7886 17356 9386
rect 18064 8650 18092 10678
rect 18156 10198 18184 11018
rect 18248 10538 18276 11018
rect 18708 10810 18736 11086
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18420 10056 18472 10062
rect 18616 10044 18644 10134
rect 18472 10016 18644 10044
rect 18696 10056 18748 10062
rect 18420 9998 18472 10004
rect 18696 9998 18748 10004
rect 18420 9920 18472 9926
rect 18512 9920 18564 9926
rect 18472 9880 18512 9908
rect 18420 9862 18472 9868
rect 18512 9862 18564 9868
rect 18708 9722 18736 9998
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 17880 8622 18092 8650
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16868 7206 16896 7686
rect 17236 7546 17264 7822
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16408 6225 16436 6394
rect 16500 6390 16528 6598
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16394 6216 16450 6225
rect 16394 6151 16450 6160
rect 17236 6118 17264 6666
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17604 6458 17632 6598
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17696 6390 17724 6734
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17316 5296 17368 5302
rect 17316 5238 17368 5244
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16304 3936 16356 3942
rect 16120 3878 16172 3884
rect 16210 3904 16266 3913
rect 16132 3738 16160 3878
rect 16304 3878 16356 3884
rect 16210 3839 16266 3848
rect 16500 3738 16528 4490
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15856 3126 15884 3538
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 15844 3120 15896 3126
rect 15844 3062 15896 3068
rect 15948 3058 15976 3334
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15948 2774 15976 2994
rect 16040 2922 16068 3334
rect 16132 2922 16160 3470
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 15948 2746 16160 2774
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15580 800 15608 2314
rect 16132 800 16160 2746
rect 16224 2310 16252 3674
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16316 3126 16344 3470
rect 16408 3194 16436 3470
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16316 2582 16344 3062
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16592 2378 16620 4558
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16684 3058 16712 4422
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 16684 800 16712 2994
rect 16776 2990 16804 4082
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16960 3777 16988 3946
rect 16946 3768 17002 3777
rect 16946 3703 17002 3712
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16868 2446 16896 3470
rect 16960 3194 16988 3606
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17052 2774 17080 4966
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17236 4282 17264 4558
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 16960 2746 17080 2774
rect 16960 2446 16988 2746
rect 17144 2689 17172 4014
rect 17236 3058 17264 4218
rect 17328 3194 17356 5238
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 3738 17448 4558
rect 17500 4548 17552 4554
rect 17500 4490 17552 4496
rect 17512 4282 17540 4490
rect 17696 4282 17724 6326
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17788 4146 17816 6054
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17498 3768 17554 3777
rect 17408 3732 17460 3738
rect 17498 3703 17554 3712
rect 17408 3674 17460 3680
rect 17512 3534 17540 3703
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17130 2680 17186 2689
rect 17130 2615 17186 2624
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 16948 2440 17000 2446
rect 17512 2417 17540 3470
rect 17604 3058 17632 3946
rect 17788 3534 17816 4082
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17696 2446 17724 3130
rect 17788 2990 17816 3470
rect 17880 3194 17908 8622
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18064 8022 18092 8434
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 18052 7880 18104 7886
rect 18156 7868 18184 8230
rect 18104 7840 18184 7868
rect 18052 7822 18104 7828
rect 18064 6934 18092 7822
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17972 3602 18000 6394
rect 18248 5370 18276 9658
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18432 6118 18460 6258
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 18064 3466 18092 4150
rect 18052 3460 18104 3466
rect 18052 3402 18104 3408
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 18064 3126 18092 3402
rect 18052 3120 18104 3126
rect 18052 3062 18104 3068
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 18248 2446 18276 5306
rect 18800 4826 18828 11086
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18892 10266 18920 10610
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18892 4758 18920 9998
rect 19168 9518 19196 11494
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19260 10810 19288 11290
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19260 9586 19288 10746
rect 19444 10470 19472 13398
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12170 20024 14962
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 20088 14414 20116 14758
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 13326 20208 13670
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19812 11694 19840 11834
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10810 20024 11698
rect 20088 11218 20116 12242
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11354 20208 12038
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 20088 10690 20116 11154
rect 20180 11082 20208 11290
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20180 10810 20208 11018
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 19996 10662 20116 10690
rect 19996 10606 20024 10662
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19996 10266 20024 10542
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19996 10130 20024 10202
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19432 9920 19484 9926
rect 19432 9862 19484 9868
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19352 6458 19380 9522
rect 19444 9110 19472 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9518 20024 10066
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8430 20024 9454
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19524 7472 19576 7478
rect 20088 7449 20116 10474
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19524 7414 19576 7420
rect 20074 7440 20130 7449
rect 19536 6730 19564 7414
rect 19984 7404 20036 7410
rect 20074 7375 20130 7384
rect 19984 7346 20036 7352
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19812 7002 19840 7278
rect 19800 6996 19852 7002
rect 19800 6938 19852 6944
rect 19524 6724 19576 6730
rect 19444 6684 19524 6712
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19340 6316 19392 6322
rect 19444 6304 19472 6684
rect 19524 6666 19576 6672
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19392 6276 19472 6304
rect 19340 6258 19392 6264
rect 19064 5636 19116 5642
rect 19064 5578 19116 5584
rect 18880 4752 18932 4758
rect 18880 4694 18932 4700
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 3194 18552 4558
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 18880 4140 18932 4146
rect 18880 4082 18932 4088
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18340 2514 18368 2994
rect 18892 2854 18920 4082
rect 18984 3126 19012 4150
rect 19076 4010 19104 5578
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 19168 3738 19196 6258
rect 19352 5710 19380 6258
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 19352 3058 19380 5170
rect 19444 3738 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19996 4706 20024 7346
rect 20180 4826 20208 9930
rect 20272 7546 20300 15370
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20364 11898 20392 12174
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20258 7440 20314 7449
rect 20258 7375 20314 7384
rect 20272 5794 20300 7375
rect 20364 5914 20392 10610
rect 20456 6458 20484 16050
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21100 15570 21128 15982
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 13938 20576 15302
rect 20732 14958 20760 15438
rect 21100 14958 21128 15506
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 20824 14822 20852 14894
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20720 14340 20772 14346
rect 20720 14282 20772 14288
rect 20732 14074 20760 14282
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20824 13870 20852 14758
rect 20994 14512 21050 14521
rect 21100 14482 21128 14894
rect 20994 14447 20996 14456
rect 21048 14447 21050 14456
rect 21088 14476 21140 14482
rect 20996 14418 21048 14424
rect 21088 14418 21140 14424
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20916 12442 20944 13738
rect 21008 13530 21036 14418
rect 21100 13870 21128 14418
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 21192 13530 21220 14010
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20548 6304 20576 10406
rect 20456 6276 20576 6304
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20272 5766 20392 5794
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 19996 4678 20116 4706
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19890 4176 19946 4185
rect 19890 4111 19946 4120
rect 19800 3936 19852 3942
rect 19798 3904 19800 3913
rect 19852 3904 19854 3913
rect 19798 3839 19854 3848
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19904 3618 19932 4111
rect 19996 3738 20024 4558
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19904 3590 20024 3618
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 3369 19472 3470
rect 19430 3360 19486 3369
rect 19430 3295 19486 3304
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19536 3058 19564 3130
rect 19996 3058 20024 3590
rect 20088 3194 20116 4678
rect 20168 4684 20220 4690
rect 20168 4626 20220 4632
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 17684 2440 17736 2446
rect 16948 2382 17000 2388
rect 17498 2408 17554 2417
rect 17224 2372 17276 2378
rect 17684 2382 17736 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 17498 2343 17554 2352
rect 17224 2314 17276 2320
rect 17236 800 17264 2314
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 17788 800 17816 2246
rect 18340 800 18368 2246
rect 18892 800 18920 2246
rect 19444 800 19472 2858
rect 20180 2774 20208 4626
rect 20272 3466 20300 5646
rect 20364 4690 20392 5766
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 20260 3460 20312 3466
rect 20260 3402 20312 3408
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20272 2990 20300 3402
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20180 2746 20300 2774
rect 20272 2650 20300 2746
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20272 2446 20300 2586
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2246
rect 20364 1970 20392 3402
rect 20456 3058 20484 6276
rect 20640 5370 20668 12106
rect 20916 11694 20944 12378
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20904 11688 20956 11694
rect 20810 11656 20866 11665
rect 20720 11620 20772 11626
rect 20904 11630 20956 11636
rect 20810 11591 20866 11600
rect 20720 11562 20772 11568
rect 20732 9926 20760 11562
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20732 9654 20760 9862
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20732 5914 20760 6326
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20536 5092 20588 5098
rect 20536 5034 20588 5040
rect 20548 3534 20576 5034
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20640 2582 20668 3878
rect 20732 2990 20760 5850
rect 20824 3738 20852 11591
rect 21008 6866 21036 11698
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21468 6798 21496 7142
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 21100 6322 21128 6666
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20916 5098 20944 6258
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 20904 5092 20956 5098
rect 20904 5034 20956 5040
rect 21376 4622 21404 5238
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20824 2774 20852 3674
rect 21468 2854 21496 4422
rect 21560 3738 21588 15370
rect 22296 15366 22324 16934
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22296 15162 22324 15302
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21546 3632 21602 3641
rect 21546 3567 21548 3576
rect 21600 3567 21602 3576
rect 21548 3538 21600 3544
rect 21652 3194 21680 14282
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21744 3670 21772 6666
rect 21928 4826 21956 14962
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 22020 14278 22048 14826
rect 22388 14482 22416 14894
rect 23032 14822 23060 36518
rect 24412 16574 24440 37198
rect 24964 37126 24992 39200
rect 25136 37256 25188 37262
rect 25136 37198 25188 37204
rect 26068 37210 26096 39200
rect 24952 37120 25004 37126
rect 24952 37062 25004 37068
rect 25148 36582 25176 37198
rect 26068 37182 26280 37210
rect 26252 37126 26280 37182
rect 27172 37126 27200 39200
rect 27252 37256 27304 37262
rect 27252 37198 27304 37204
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 26148 37120 26200 37126
rect 26148 37062 26200 37068
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 26160 36582 26188 37062
rect 27264 36582 27292 37198
rect 28184 36582 28212 37198
rect 28276 37126 28304 39200
rect 29380 37346 29408 39200
rect 29380 37318 29500 37346
rect 29368 37256 29420 37262
rect 29368 37198 29420 37204
rect 28264 37120 28316 37126
rect 28264 37062 28316 37068
rect 29380 36582 29408 37198
rect 29472 37126 29500 37318
rect 30380 37256 30432 37262
rect 30380 37198 30432 37204
rect 29460 37120 29512 37126
rect 29460 37062 29512 37068
rect 30392 36582 30420 37198
rect 30484 37126 30512 39200
rect 31484 37324 31536 37330
rect 31484 37266 31536 37272
rect 30472 37120 30524 37126
rect 30472 37062 30524 37068
rect 25136 36576 25188 36582
rect 25136 36518 25188 36524
rect 26148 36576 26200 36582
rect 26148 36518 26200 36524
rect 27252 36576 27304 36582
rect 27252 36518 27304 36524
rect 28172 36576 28224 36582
rect 28172 36518 28224 36524
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 30380 36576 30432 36582
rect 30380 36518 30432 36524
rect 24320 16546 24440 16574
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 24124 14340 24176 14346
rect 24124 14282 24176 14288
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22204 14074 22232 14214
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 22020 6254 22048 6734
rect 22388 6458 22416 13874
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 22742 6760 22798 6769
rect 22742 6695 22798 6704
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22756 6390 22784 6695
rect 22744 6384 22796 6390
rect 22744 6326 22796 6332
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22020 5370 22048 6190
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 22112 4706 22140 5170
rect 22112 4678 22232 4706
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21732 3664 21784 3670
rect 21732 3606 21784 3612
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 20824 2746 20944 2774
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20916 2446 20944 2746
rect 21640 2576 21692 2582
rect 21640 2518 21692 2524
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 20536 2304 20588 2310
rect 20536 2246 20588 2252
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 20352 1964 20404 1970
rect 20352 1906 20404 1912
rect 20548 800 20576 2246
rect 21100 800 21128 2246
rect 21652 800 21680 2518
rect 21744 2009 21772 3470
rect 21836 3466 21864 4014
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21836 3369 21864 3402
rect 21822 3360 21878 3369
rect 21822 3295 21878 3304
rect 21836 2990 21864 3295
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21928 2106 21956 4422
rect 22112 4282 22140 4558
rect 22100 4276 22152 4282
rect 22100 4218 22152 4224
rect 22008 4208 22060 4214
rect 22006 4176 22008 4185
rect 22060 4176 22062 4185
rect 22006 4111 22062 4120
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22112 3942 22140 4082
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 21916 2100 21968 2106
rect 21916 2042 21968 2048
rect 22020 2038 22048 2994
rect 22112 2514 22140 3674
rect 22204 3194 22232 4678
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22296 3040 22324 4082
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 22388 3398 22416 3538
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22388 3058 22416 3334
rect 22204 3012 22324 3040
rect 22376 3052 22428 3058
rect 22204 2854 22232 3012
rect 22376 2994 22428 3000
rect 22284 2916 22336 2922
rect 22284 2858 22336 2864
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22296 2446 22324 2858
rect 22284 2440 22336 2446
rect 22284 2382 22336 2388
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22008 2032 22060 2038
rect 21730 2000 21786 2009
rect 22008 1974 22060 1980
rect 21730 1935 21786 1944
rect 22204 800 22232 2246
rect 22480 1834 22508 4082
rect 22572 4010 22600 6258
rect 23492 4826 23520 13330
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23112 4208 23164 4214
rect 23112 4150 23164 4156
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 22744 4072 22796 4078
rect 22744 4014 22796 4020
rect 22560 4004 22612 4010
rect 22560 3946 22612 3952
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 22572 3369 22600 3402
rect 22558 3360 22614 3369
rect 22558 3295 22614 3304
rect 22558 3224 22614 3233
rect 22558 3159 22614 3168
rect 22572 3126 22600 3159
rect 22560 3120 22612 3126
rect 22560 3062 22612 3068
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22572 1873 22600 2790
rect 22558 1864 22614 1873
rect 22468 1828 22520 1834
rect 22558 1799 22614 1808
rect 22468 1770 22520 1776
rect 22664 1698 22692 3878
rect 22756 3738 22784 4014
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22756 3618 22784 3674
rect 22756 3590 22876 3618
rect 22940 3602 22968 4082
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22756 2553 22784 3470
rect 22848 2854 22876 3590
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 23124 3398 23152 4150
rect 23216 4146 23244 4422
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23124 3126 23152 3334
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 23308 3058 23336 3470
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23032 2961 23060 2994
rect 23112 2984 23164 2990
rect 23018 2952 23074 2961
rect 23112 2926 23164 2932
rect 23018 2887 23074 2896
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22742 2544 22798 2553
rect 22742 2479 22798 2488
rect 22744 2372 22796 2378
rect 22744 2314 22796 2320
rect 22652 1692 22704 1698
rect 22652 1634 22704 1640
rect 22756 800 22784 2314
rect 23124 2038 23152 2926
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23112 2032 23164 2038
rect 23112 1974 23164 1980
rect 23308 800 23336 2858
rect 23492 2446 23520 4762
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23584 2106 23612 4218
rect 23756 4208 23808 4214
rect 23754 4176 23756 4185
rect 23808 4176 23810 4185
rect 24136 4146 24164 14282
rect 24320 14278 24348 16546
rect 24400 14884 24452 14890
rect 24400 14826 24452 14832
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24412 4826 24440 14826
rect 25148 14006 25176 36518
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 25136 13456 25188 13462
rect 25136 13398 25188 13404
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24780 4622 24808 5170
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24780 4146 24808 4558
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 23754 4111 23810 4120
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 24228 3097 24256 3538
rect 24308 3460 24360 3466
rect 24308 3402 24360 3408
rect 24214 3088 24270 3097
rect 24214 3023 24216 3032
rect 24268 3023 24270 3032
rect 24216 2994 24268 3000
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23572 2100 23624 2106
rect 23572 2042 23624 2048
rect 23860 800 23888 2790
rect 24320 2774 24348 3402
rect 24412 3194 24440 4082
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24780 3534 24808 3878
rect 24964 3738 24992 4490
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 24768 3528 24820 3534
rect 24766 3496 24768 3505
rect 24820 3496 24822 3505
rect 24584 3460 24636 3466
rect 24766 3431 24822 3440
rect 24860 3460 24912 3466
rect 24584 3402 24636 3408
rect 24860 3402 24912 3408
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24320 2746 24532 2774
rect 24504 1902 24532 2746
rect 24596 2514 24624 3402
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24872 2446 24900 3402
rect 25148 3058 25176 13398
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25608 4146 25636 12922
rect 26160 11626 26188 36518
rect 27264 16658 27292 36518
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 28184 14414 28212 36518
rect 29380 15638 29408 36518
rect 29368 15632 29420 15638
rect 29368 15574 29420 15580
rect 30392 15094 30420 36518
rect 31496 15366 31524 37266
rect 31588 37108 31616 39200
rect 32692 37126 32720 39200
rect 32864 37256 32916 37262
rect 32864 37198 32916 37204
rect 31760 37120 31812 37126
rect 31588 37080 31760 37108
rect 31760 37062 31812 37068
rect 32680 37120 32732 37126
rect 32680 37062 32732 37068
rect 32876 36582 32904 37198
rect 33796 37126 33824 39200
rect 34900 37754 34928 39200
rect 34808 37726 34928 37754
rect 34808 37346 34836 37726
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34808 37318 34928 37346
rect 33876 37256 33928 37262
rect 33876 37198 33928 37204
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 33784 37120 33836 37126
rect 33784 37062 33836 37068
rect 33888 36582 33916 37198
rect 34808 36582 34836 37198
rect 34900 37126 34928 37318
rect 35900 37256 35952 37262
rect 35900 37198 35952 37204
rect 34888 37120 34940 37126
rect 34888 37062 34940 37068
rect 35912 36582 35940 37198
rect 36004 37126 36032 39200
rect 37108 37126 37136 39200
rect 37372 37256 37424 37262
rect 37372 37198 37424 37204
rect 35992 37120 36044 37126
rect 35992 37062 36044 37068
rect 37096 37120 37148 37126
rect 37096 37062 37148 37068
rect 37384 36582 37412 37198
rect 38016 37120 38068 37126
rect 38016 37062 38068 37068
rect 38028 36786 38056 37062
rect 38212 36922 38240 39200
rect 38200 36916 38252 36922
rect 38200 36858 38252 36864
rect 37832 36780 37884 36786
rect 37832 36722 37884 36728
rect 38016 36780 38068 36786
rect 38016 36722 38068 36728
rect 32864 36576 32916 36582
rect 32864 36518 32916 36524
rect 33876 36576 33928 36582
rect 33876 36518 33928 36524
rect 34796 36576 34848 36582
rect 34796 36518 34848 36524
rect 35900 36576 35952 36582
rect 35900 36518 35952 36524
rect 37372 36576 37424 36582
rect 37372 36518 37424 36524
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 30380 15088 30432 15094
rect 30380 15030 30432 15036
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 27620 13252 27672 13258
rect 27620 13194 27672 13200
rect 26148 11620 26200 11626
rect 26148 11562 26200 11568
rect 26516 9172 26568 9178
rect 26516 9114 26568 9120
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 26252 4146 26280 8978
rect 25596 4140 25648 4146
rect 25596 4082 25648 4088
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 25608 3058 25636 4082
rect 26054 3632 26110 3641
rect 26054 3567 26110 3576
rect 26068 3466 26096 3567
rect 26056 3460 26108 3466
rect 26056 3402 26108 3408
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 26056 2916 26108 2922
rect 26056 2858 26108 2864
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 24492 1896 24544 1902
rect 24492 1838 24544 1844
rect 24872 1766 24900 2382
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 25056 1442 25084 2790
rect 25240 2650 25268 2858
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25964 2576 26016 2582
rect 25964 2518 26016 2524
rect 25504 2372 25556 2378
rect 25504 2314 25556 2320
rect 24400 1420 24452 1426
rect 24400 1362 24452 1368
rect 24964 1414 25084 1442
rect 24412 800 24440 1362
rect 24964 800 24992 1414
rect 25516 800 25544 2314
rect 25976 1426 26004 2518
rect 25964 1420 26016 1426
rect 25964 1362 26016 1368
rect 26068 800 26096 2858
rect 26252 2446 26280 4082
rect 26528 3738 26556 9114
rect 27068 8968 27120 8974
rect 27068 8910 27120 8916
rect 27080 3738 27108 8910
rect 27632 3738 27660 13194
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 26516 3732 26568 3738
rect 26516 3674 26568 3680
rect 27068 3732 27120 3738
rect 27068 3674 27120 3680
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 26330 3224 26386 3233
rect 26330 3159 26386 3168
rect 26344 2854 26372 3159
rect 26332 2848 26384 2854
rect 26332 2790 26384 2796
rect 26528 2514 26556 3674
rect 27080 3058 27108 3674
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 26608 2576 26660 2582
rect 26608 2518 26660 2524
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 26620 800 26648 2518
rect 26896 2378 27108 2394
rect 26884 2372 27108 2378
rect 26936 2366 27108 2372
rect 26884 2314 26936 2320
rect 27080 2310 27108 2366
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27172 800 27200 2994
rect 27540 2689 27568 3062
rect 27526 2680 27582 2689
rect 27526 2615 27582 2624
rect 27632 2446 27660 3674
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 27908 3058 27936 3334
rect 28552 3058 28580 3334
rect 27896 3052 27948 3058
rect 27896 2994 27948 3000
rect 28264 3052 28316 3058
rect 28264 2994 28316 3000
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 27724 800 27752 2314
rect 28276 800 28304 2994
rect 28632 2916 28684 2922
rect 28632 2858 28684 2864
rect 28644 2446 28672 2858
rect 28828 2582 28856 6394
rect 29012 3194 29040 11834
rect 32876 10062 32904 36518
rect 32864 10056 32916 10062
rect 32864 9998 32916 10004
rect 33888 9926 33916 36518
rect 34808 11150 34836 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 35912 10606 35940 36518
rect 37280 36032 37332 36038
rect 37280 35974 37332 35980
rect 35900 10600 35952 10606
rect 35900 10542 35952 10548
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 33876 9920 33928 9926
rect 33876 9862 33928 9868
rect 37292 9450 37320 35974
rect 37384 11830 37412 36518
rect 37372 11824 37424 11830
rect 37372 11766 37424 11772
rect 37844 11082 37872 36722
rect 39316 36378 39344 39200
rect 39304 36372 39356 36378
rect 39304 36314 39356 36320
rect 37832 11076 37884 11082
rect 37832 11018 37884 11024
rect 37280 9444 37332 9450
rect 37280 9386 37332 9392
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34428 4480 34480 4486
rect 34428 4422 34480 4428
rect 33324 4208 33376 4214
rect 33324 4150 33376 4156
rect 33138 4040 33194 4049
rect 33138 3975 33194 3984
rect 31208 3460 31260 3466
rect 31208 3402 31260 3408
rect 29552 3392 29604 3398
rect 29552 3334 29604 3340
rect 30748 3392 30800 3398
rect 30748 3334 30800 3340
rect 29000 3188 29052 3194
rect 29000 3130 29052 3136
rect 28816 2576 28868 2582
rect 29012 2564 29040 3130
rect 29012 2536 29132 2564
rect 28816 2518 28868 2524
rect 28632 2440 28684 2446
rect 29000 2440 29052 2446
rect 28632 2382 28684 2388
rect 28828 2400 29000 2428
rect 28828 800 28856 2400
rect 29000 2382 29052 2388
rect 29104 2378 29132 2536
rect 29564 2446 29592 3334
rect 30760 3058 30788 3334
rect 31220 3194 31248 3402
rect 31392 3392 31444 3398
rect 31392 3334 31444 3340
rect 31208 3188 31260 3194
rect 31208 3130 31260 3136
rect 31404 3058 31432 3334
rect 30472 3052 30524 3058
rect 30472 2994 30524 3000
rect 30748 3052 30800 3058
rect 30748 2994 30800 3000
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 31392 3052 31444 3058
rect 31392 2994 31444 3000
rect 29920 2508 29972 2514
rect 29920 2450 29972 2456
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29092 2372 29144 2378
rect 29092 2314 29144 2320
rect 29368 2372 29420 2378
rect 29368 2314 29420 2320
rect 29380 800 29408 2314
rect 29552 2304 29604 2310
rect 29552 2246 29604 2252
rect 29564 2106 29592 2246
rect 29552 2100 29604 2106
rect 29552 2042 29604 2048
rect 29932 800 29960 2450
rect 30196 2304 30248 2310
rect 30196 2246 30248 2252
rect 30208 1902 30236 2246
rect 30196 1896 30248 1902
rect 30196 1838 30248 1844
rect 30484 800 30512 2994
rect 31036 800 31064 2994
rect 33152 2922 33180 3975
rect 33232 3392 33284 3398
rect 33232 3334 33284 3340
rect 33244 3058 33272 3334
rect 33336 3194 33364 4150
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33324 3188 33376 3194
rect 33324 3130 33376 3136
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 33140 2916 33192 2922
rect 33140 2858 33192 2864
rect 31484 2848 31536 2854
rect 31484 2790 31536 2796
rect 32680 2848 32732 2854
rect 32680 2790 32732 2796
rect 31496 2514 31524 2790
rect 31484 2508 31536 2514
rect 31484 2450 31536 2456
rect 32692 2446 32720 2790
rect 31760 2440 31812 2446
rect 31588 2400 31760 2428
rect 31588 800 31616 2400
rect 31760 2382 31812 2388
rect 32680 2440 32732 2446
rect 33140 2440 33192 2446
rect 32680 2382 32732 2388
rect 33060 2400 33140 2428
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 32128 2304 32180 2310
rect 32128 2246 32180 2252
rect 32140 2038 32168 2246
rect 32128 2032 32180 2038
rect 32128 1974 32180 1980
rect 32232 1850 32260 2314
rect 32772 2304 32824 2310
rect 32772 2246 32824 2252
rect 32140 1822 32260 1850
rect 32784 1834 32812 2246
rect 32772 1828 32824 1834
rect 32140 800 32168 1822
rect 32772 1770 32824 1776
rect 32692 870 32812 898
rect 32692 800 32720 870
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11702 0 11758 800
rect 12254 0 12310 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23294 0 23350 800
rect 23846 0 23902 800
rect 24398 0 24454 800
rect 24950 0 25006 800
rect 25502 0 25558 800
rect 26054 0 26110 800
rect 26606 0 26662 800
rect 27158 0 27214 800
rect 27710 0 27766 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29366 0 29422 800
rect 29918 0 29974 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 32784 762 32812 870
rect 33060 762 33088 2400
rect 33140 2382 33192 2388
rect 33244 800 33272 2994
rect 33704 2446 33732 3334
rect 34440 3210 34468 4422
rect 36636 4140 36688 4146
rect 36636 4082 36688 4088
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36648 3738 36676 4082
rect 36636 3732 36688 3738
rect 36636 3674 36688 3680
rect 36544 3528 36596 3534
rect 36544 3470 36596 3476
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35992 3392 36044 3398
rect 35992 3334 36044 3340
rect 34440 3194 34560 3210
rect 34440 3188 34572 3194
rect 34440 3182 34520 3188
rect 34520 3130 34572 3136
rect 34336 3052 34388 3058
rect 34336 2994 34388 3000
rect 33692 2440 33744 2446
rect 33692 2382 33744 2388
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33416 2304 33468 2310
rect 33416 2246 33468 2252
rect 33428 1970 33456 2246
rect 33416 1964 33468 1970
rect 33416 1906 33468 1912
rect 33796 800 33824 2382
rect 34348 800 34376 2994
rect 34716 2446 34744 3334
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34704 2440 34756 2446
rect 34518 2408 34574 2417
rect 34980 2440 35032 2446
rect 34704 2382 34756 2388
rect 34900 2400 34980 2428
rect 34518 2343 34574 2352
rect 34532 2310 34560 2343
rect 34520 2304 34572 2310
rect 34520 2246 34572 2252
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 34808 1698 34836 2246
rect 34796 1692 34848 1698
rect 34796 1634 34848 1640
rect 34900 800 34928 2400
rect 34980 2382 35032 2388
rect 35820 2394 35848 3334
rect 36004 3058 36032 3334
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 35900 2440 35952 2446
rect 35820 2388 35900 2394
rect 35820 2382 35952 2388
rect 35820 2366 35940 2382
rect 35452 870 35572 898
rect 35452 800 35480 870
rect 32784 734 33088 762
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35438 0 35494 800
rect 35544 762 35572 870
rect 35820 762 35848 2366
rect 36004 800 36032 2994
rect 36556 800 36584 3470
rect 37096 3052 37148 3058
rect 37096 2994 37148 3000
rect 37108 800 37136 2994
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 37660 800 37688 2450
rect 37844 2446 37872 6054
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 38028 2514 38056 3334
rect 38016 2508 38068 2514
rect 38016 2450 38068 2456
rect 37832 2440 37884 2446
rect 37832 2382 37884 2388
rect 35544 734 35848 762
rect 35990 0 36046 800
rect 36542 0 36598 800
rect 37094 0 37150 800
rect 37646 0 37702 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1582 29960 1638 30016
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 3422 9968 3478 10024
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3790 6160 3846 6216
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5814 2524 5816 2544
rect 5816 2524 5868 2544
rect 5868 2524 5870 2544
rect 5814 2488 5870 2524
rect 7746 11600 7802 11656
rect 7378 4120 7434 4176
rect 7746 1944 7802 2000
rect 9586 1808 9642 1864
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 15750 14456 15806 14512
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 11794 6996 11850 7032
rect 11794 6976 11796 6996
rect 11796 6976 11848 6996
rect 11848 6976 11850 6996
rect 12714 6704 12770 6760
rect 11610 3440 11666 3496
rect 11334 3032 11390 3088
rect 13266 6704 13322 6760
rect 14094 6976 14150 7032
rect 11886 2916 11942 2952
rect 11886 2896 11888 2916
rect 11888 2896 11940 2916
rect 11940 2896 11942 2916
rect 13542 3304 13598 3360
rect 14922 2760 14978 2816
rect 15658 3984 15714 4040
rect 15382 2760 15438 2816
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 16394 6160 16450 6216
rect 16210 3848 16266 3904
rect 16946 3712 17002 3768
rect 17498 3712 17554 3768
rect 17130 2624 17186 2680
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 20074 7384 20130 7440
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 20258 7384 20314 7440
rect 20994 14476 21050 14512
rect 20994 14456 20996 14476
rect 20996 14456 21048 14476
rect 21048 14456 21050 14476
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19890 4120 19946 4176
rect 19798 3884 19800 3904
rect 19800 3884 19852 3904
rect 19852 3884 19854 3904
rect 19798 3848 19854 3884
rect 19430 3304 19486 3360
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 17498 2352 17554 2408
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20810 11600 20866 11656
rect 21546 3596 21602 3632
rect 21546 3576 21548 3596
rect 21548 3576 21600 3596
rect 21600 3576 21602 3596
rect 22742 6704 22798 6760
rect 21822 3304 21878 3360
rect 22006 4156 22008 4176
rect 22008 4156 22060 4176
rect 22060 4156 22062 4176
rect 22006 4120 22062 4156
rect 21730 1944 21786 2000
rect 22558 3304 22614 3360
rect 22558 3168 22614 3224
rect 22558 1808 22614 1864
rect 23018 2896 23074 2952
rect 22742 2488 22798 2544
rect 23754 4156 23756 4176
rect 23756 4156 23808 4176
rect 23808 4156 23810 4176
rect 23754 4120 23810 4156
rect 24214 3052 24270 3088
rect 24214 3032 24216 3052
rect 24216 3032 24268 3052
rect 24268 3032 24270 3052
rect 24766 3476 24768 3496
rect 24768 3476 24820 3496
rect 24820 3476 24822 3496
rect 24766 3440 24822 3476
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 26054 3576 26110 3632
rect 26330 3168 26386 3224
rect 27526 2624 27582 2680
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 33138 3984 33194 4040
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 34518 2352 34574 2408
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 0 30018 800 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 800 29958
rect 1577 29955 1643 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 15745 14514 15811 14517
rect 20989 14514 21055 14517
rect 15745 14512 21055 14514
rect 15745 14456 15750 14512
rect 15806 14456 20994 14512
rect 21050 14456 21055 14512
rect 15745 14454 21055 14456
rect 15745 14451 15811 14454
rect 20989 14451 21055 14454
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 7741 11658 7807 11661
rect 20805 11658 20871 11661
rect 7741 11656 20871 11658
rect 7741 11600 7746 11656
rect 7802 11600 20810 11656
rect 20866 11600 20871 11656
rect 7741 11598 20871 11600
rect 7741 11595 7807 11598
rect 20805 11595 20871 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 0 10026 800 10056
rect 3417 10026 3483 10029
rect 0 10024 3483 10026
rect 0 9968 3422 10024
rect 3478 9968 3483 10024
rect 0 9966 3483 9968
rect 0 9936 800 9966
rect 3417 9963 3483 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 20069 7442 20135 7445
rect 20253 7442 20319 7445
rect 20069 7440 20319 7442
rect 20069 7384 20074 7440
rect 20130 7384 20258 7440
rect 20314 7384 20319 7440
rect 20069 7382 20319 7384
rect 20069 7379 20135 7382
rect 20253 7379 20319 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 11789 7034 11855 7037
rect 14089 7034 14155 7037
rect 11789 7032 14155 7034
rect 11789 6976 11794 7032
rect 11850 6976 14094 7032
rect 14150 6976 14155 7032
rect 11789 6974 14155 6976
rect 11789 6971 11855 6974
rect 14089 6971 14155 6974
rect 12709 6762 12775 6765
rect 13261 6762 13327 6765
rect 22737 6762 22803 6765
rect 12709 6760 22803 6762
rect 12709 6704 12714 6760
rect 12770 6704 13266 6760
rect 13322 6704 22742 6760
rect 22798 6704 22803 6760
rect 12709 6702 22803 6704
rect 12709 6699 12775 6702
rect 13261 6699 13327 6702
rect 22737 6699 22803 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 3785 6218 3851 6221
rect 16389 6218 16455 6221
rect 3785 6216 16455 6218
rect 3785 6160 3790 6216
rect 3846 6160 16394 6216
rect 16450 6160 16455 6216
rect 3785 6158 16455 6160
rect 3785 6155 3851 6158
rect 16389 6155 16455 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 7373 4178 7439 4181
rect 19885 4178 19951 4181
rect 7373 4176 19951 4178
rect 7373 4120 7378 4176
rect 7434 4120 19890 4176
rect 19946 4120 19951 4176
rect 7373 4118 19951 4120
rect 7373 4115 7439 4118
rect 19885 4115 19951 4118
rect 22001 4178 22067 4181
rect 23749 4178 23815 4181
rect 22001 4176 23815 4178
rect 22001 4120 22006 4176
rect 22062 4120 23754 4176
rect 23810 4120 23815 4176
rect 22001 4118 23815 4120
rect 22001 4115 22067 4118
rect 23749 4115 23815 4118
rect 15653 4042 15719 4045
rect 33133 4042 33199 4045
rect 15653 4040 33199 4042
rect 15653 3984 15658 4040
rect 15714 3984 33138 4040
rect 33194 3984 33199 4040
rect 15653 3982 33199 3984
rect 15653 3979 15719 3982
rect 33133 3979 33199 3982
rect 16205 3906 16271 3909
rect 19793 3906 19859 3909
rect 16205 3904 19859 3906
rect 16205 3848 16210 3904
rect 16266 3848 19798 3904
rect 19854 3848 19859 3904
rect 16205 3846 19859 3848
rect 16205 3843 16271 3846
rect 19793 3843 19859 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 16941 3770 17007 3773
rect 17493 3770 17559 3773
rect 16941 3768 17559 3770
rect 16941 3712 16946 3768
rect 17002 3712 17498 3768
rect 17554 3712 17559 3768
rect 16941 3710 17559 3712
rect 16941 3707 17007 3710
rect 17493 3707 17559 3710
rect 21541 3634 21607 3637
rect 26049 3634 26115 3637
rect 21541 3632 26115 3634
rect 21541 3576 21546 3632
rect 21602 3576 26054 3632
rect 26110 3576 26115 3632
rect 21541 3574 26115 3576
rect 21541 3571 21607 3574
rect 26049 3571 26115 3574
rect 11605 3498 11671 3501
rect 24761 3498 24827 3501
rect 11605 3496 24827 3498
rect 11605 3440 11610 3496
rect 11666 3440 24766 3496
rect 24822 3440 24827 3496
rect 11605 3438 24827 3440
rect 11605 3435 11671 3438
rect 24761 3435 24827 3438
rect 13537 3362 13603 3365
rect 19425 3362 19491 3365
rect 13537 3360 19491 3362
rect 13537 3304 13542 3360
rect 13598 3304 19430 3360
rect 19486 3304 19491 3360
rect 13537 3302 19491 3304
rect 13537 3299 13603 3302
rect 19425 3299 19491 3302
rect 21817 3362 21883 3365
rect 22553 3362 22619 3365
rect 21817 3360 22619 3362
rect 21817 3304 21822 3360
rect 21878 3304 22558 3360
rect 22614 3304 22619 3360
rect 21817 3302 22619 3304
rect 21817 3299 21883 3302
rect 22553 3299 22619 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 22553 3226 22619 3229
rect 26325 3226 26391 3229
rect 22553 3224 26391 3226
rect 22553 3168 22558 3224
rect 22614 3168 26330 3224
rect 26386 3168 26391 3224
rect 22553 3166 26391 3168
rect 22553 3163 22619 3166
rect 26325 3163 26391 3166
rect 11329 3090 11395 3093
rect 24209 3090 24275 3093
rect 11329 3088 24275 3090
rect 11329 3032 11334 3088
rect 11390 3032 24214 3088
rect 24270 3032 24275 3088
rect 11329 3030 24275 3032
rect 11329 3027 11395 3030
rect 24209 3027 24275 3030
rect 11881 2954 11947 2957
rect 23013 2954 23079 2957
rect 11881 2952 23079 2954
rect 11881 2896 11886 2952
rect 11942 2896 23018 2952
rect 23074 2896 23079 2952
rect 11881 2894 23079 2896
rect 11881 2891 11947 2894
rect 23013 2891 23079 2894
rect 14917 2818 14983 2821
rect 15377 2818 15443 2821
rect 14917 2816 15443 2818
rect 14917 2760 14922 2816
rect 14978 2760 15382 2816
rect 15438 2760 15443 2816
rect 14917 2758 15443 2760
rect 14917 2755 14983 2758
rect 15377 2755 15443 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 17125 2682 17191 2685
rect 27521 2682 27587 2685
rect 17125 2680 27587 2682
rect 17125 2624 17130 2680
rect 17186 2624 27526 2680
rect 27582 2624 27587 2680
rect 17125 2622 27587 2624
rect 17125 2619 17191 2622
rect 27521 2619 27587 2622
rect 5809 2546 5875 2549
rect 22737 2546 22803 2549
rect 5809 2544 22803 2546
rect 5809 2488 5814 2544
rect 5870 2488 22742 2544
rect 22798 2488 22803 2544
rect 5809 2486 22803 2488
rect 5809 2483 5875 2486
rect 22737 2483 22803 2486
rect 17493 2410 17559 2413
rect 34513 2410 34579 2413
rect 17493 2408 34579 2410
rect 17493 2352 17498 2408
rect 17554 2352 34518 2408
rect 34574 2352 34579 2408
rect 17493 2350 34579 2352
rect 17493 2347 17559 2350
rect 34513 2347 34579 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 7741 2002 7807 2005
rect 21725 2002 21791 2005
rect 7741 2000 21791 2002
rect 7741 1944 7746 2000
rect 7802 1944 21730 2000
rect 21786 1944 21791 2000
rect 7741 1942 21791 1944
rect 7741 1939 7807 1942
rect 21725 1939 21791 1942
rect 9581 1866 9647 1869
rect 22553 1866 22619 1869
rect 9581 1864 22619 1866
rect 9581 1808 9586 1864
rect 9642 1808 22558 1864
rect 22614 1808 22619 1864
rect 9581 1806 22619 1808
rect 9581 1803 9647 1806
rect 22553 1803 22619 1806
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A2
timestamp 1649977179
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__B1
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__C
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A1
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A2
timestamp 1649977179
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__C1
timestamp 1649977179
transform 1 0 11960 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A2
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__B
timestamp 1649977179
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A1
timestamp 1649977179
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A2
timestamp 1649977179
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__C1
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__B
timestamp 1649977179
transform -1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1649977179
transform -1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1649977179
transform -1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1649977179
transform -1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__B1
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A1
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__B2
timestamp 1649977179
transform 1 0 6072 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A0
timestamp 1649977179
transform -1 0 4416 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A1
timestamp 1649977179
transform -1 0 3036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A0
timestamp 1649977179
transform -1 0 4968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A1
timestamp 1649977179
transform -1 0 3864 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A0
timestamp 1649977179
transform 1 0 4968 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A1
timestamp 1649977179
transform -1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A0
timestamp 1649977179
transform 1 0 6532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__233__A1
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A0
timestamp 1649977179
transform -1 0 8280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__A1
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A0
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A1
timestamp 1649977179
transform -1 0 8464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A0
timestamp 1649977179
transform -1 0 9292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A1
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A0
timestamp 1649977179
transform -1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__A1
timestamp 1649977179
transform 1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A0
timestamp 1649977179
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A1
timestamp 1649977179
transform -1 0 9568 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A0
timestamp 1649977179
transform -1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A1
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__S
timestamp 1649977179
transform 1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A0
timestamp 1649977179
transform -1 0 13340 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A1
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__S
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A0
timestamp 1649977179
transform -1 0 14260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A1
timestamp 1649977179
transform -1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__S
timestamp 1649977179
transform -1 0 12880 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A0
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A1
timestamp 1649977179
transform -1 0 10580 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__S
timestamp 1649977179
transform -1 0 11132 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A0
timestamp 1649977179
transform -1 0 18032 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__S
timestamp 1649977179
transform 1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A0
timestamp 1649977179
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A1
timestamp 1649977179
transform -1 0 16652 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__S
timestamp 1649977179
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A0
timestamp 1649977179
transform -1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A1
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__S
timestamp 1649977179
transform 1 0 17204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__B
timestamp 1649977179
transform 1 0 9384 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A1
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__290__A2
timestamp 1649977179
transform -1 0 25208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A1
timestamp 1649977179
transform -1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A2
timestamp 1649977179
transform -1 0 25576 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A1
timestamp 1649977179
transform -1 0 21988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A2
timestamp 1649977179
transform -1 0 23092 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A1
timestamp 1649977179
transform 1 0 23276 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A1
timestamp 1649977179
transform -1 0 21344 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__303__A1
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__304__A1
timestamp 1649977179
transform -1 0 19964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__A_N
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__B
timestamp 1649977179
transform -1 0 19412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__308__A1
timestamp 1649977179
transform 1 0 19872 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__311__A1
timestamp 1649977179
transform -1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__314__A1
timestamp 1649977179
transform 1 0 21712 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__318__A1
timestamp 1649977179
transform -1 0 17664 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__322__A1
timestamp 1649977179
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__A1
timestamp 1649977179
transform -1 0 19504 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__A1
timestamp 1649977179
transform -1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__332__B1
timestamp 1649977179
transform -1 0 16928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__334__A1
timestamp 1649977179
transform 1 0 18216 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A1
timestamp 1649977179
transform -1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__B1
timestamp 1649977179
transform -1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1
timestamp 1649977179
transform -1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__B1
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A1
timestamp 1649977179
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A
timestamp 1649977179
transform -1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A1
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A1
timestamp 1649977179
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A2
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A0
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A0
timestamp 1649977179
transform -1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_i_clk_A
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2944 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 4048 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 15088 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 16192 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 17296 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 18400 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 19504 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 20608 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 5152 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 6532 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 7360 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 8464 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 9568 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 10672 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 11776 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 12880 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 14076 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 1748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 12880 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 13064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 4600 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 14168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 14720 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 5428 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 5704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 6256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 15456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 28336 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 33856 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 33304 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 34868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 35236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 36800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 35512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 29716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 28888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 29716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 32292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 30544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 31188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 32844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 36064 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 37444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 38180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output67_A
timestamp 1649977179
transform 1 0 2208 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1649977179
transform -1 0 21988 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output69_A
timestamp 1649977179
transform 1 0 32660 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform 1 0 33672 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1649977179
transform 1 0 34776 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform 1 0 35880 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1649977179
transform -1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output74_A
timestamp 1649977179
transform -1 0 38180 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1649977179
transform 1 0 22632 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform -1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1649977179
transform 1 0 24932 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1649977179
transform 1 0 25944 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1649977179
transform 1 0 27048 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output80_A
timestamp 1649977179
transform 1 0 28152 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1649977179
transform 1 0 29348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1649977179
transform 1 0 30360 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1649977179
transform -1 0 31648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1649977179
transform -1 0 37444 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1649977179
transform 1 0 16744 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform -1 0 26496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1649977179
transform -1 0 26312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1649977179
transform -1 0 25760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1649977179
transform -1 0 27784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1649977179
transform -1 0 27232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1649977179
transform -1 0 29164 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1649977179
transform 1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1649977179
transform -1 0 21160 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1649977179
transform -1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform 1 0 19320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1649977179
transform 1 0 20976 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output99_A
timestamp 1649977179
transform -1 0 23736 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output100_A
timestamp 1649977179
transform -1 0 23644 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1649977179
transform -1 0 26128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output102_A
timestamp 1649977179
transform -1 0 26680 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1649977179
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1649977179
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_200
timestamp 1649977179
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1649977179
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1649977179
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_229
timestamp 1649977179
transform 1 0 22172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1649977179
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1649977179
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285
timestamp 1649977179
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1649977179
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_312
timestamp 1649977179
transform 1 0 29808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_319
timestamp 1649977179
transform 1 0 30452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_326
timestamp 1649977179
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_340
timestamp 1649977179
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_354
timestamp 1649977179
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_11
timestamp 1649977179
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_16
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_24
timestamp 1649977179
transform 1 0 3312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1649977179
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_65
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_83
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_91
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_95
timestamp 1649977179
transform 1 0 9844 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1649977179
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1649977179
transform 1 0 12788 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_130
timestamp 1649977179
transform 1 0 13064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_154
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_160
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_182
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_212
timestamp 1649977179
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1649977179
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1649977179
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1649977179
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1649977179
transform 1 0 24472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_270
timestamp 1649977179
transform 1 0 25944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_292
timestamp 1649977179
transform 1 0 27968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1649977179
transform 1 0 28612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_311
timestamp 1649977179
transform 1 0 29716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_319
timestamp 1649977179
transform 1 0 30452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_323
timestamp 1649977179
transform 1 0 30820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_330
timestamp 1649977179
transform 1 0 31464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_339
timestamp 1649977179
transform 1 0 32292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_345
timestamp 1649977179
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_353
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_365
timestamp 1649977179
transform 1 0 34684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_371
timestamp 1649977179
transform 1 0 35236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_379
timestamp 1649977179
transform 1 0 35972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_383
timestamp 1649977179
transform 1 0 36340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_397
timestamp 1649977179
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1649977179
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_38
timestamp 1649977179
transform 1 0 4600 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_56
timestamp 1649977179
transform 1 0 6256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1649977179
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_92
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_96
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_114
timestamp 1649977179
transform 1 0 11592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_120
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_134
timestamp 1649977179
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1649977179
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_162
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_169
timestamp 1649977179
transform 1 0 16652 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1649977179
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_199
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_212
timestamp 1649977179
transform 1 0 20608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1649977179
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1649977179
transform 1 0 22172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1649977179
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1649977179
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_260
timestamp 1649977179
transform 1 0 25024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_266
timestamp 1649977179
transform 1 0 25576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_272
timestamp 1649977179
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_278
timestamp 1649977179
transform 1 0 26680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_284
timestamp 1649977179
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_290
timestamp 1649977179
transform 1 0 27784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_296
timestamp 1649977179
transform 1 0 28336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1649977179
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_311
timestamp 1649977179
transform 1 0 29716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_317
timestamp 1649977179
transform 1 0 30268 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_320
timestamp 1649977179
transform 1 0 30544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_324
timestamp 1649977179
transform 1 0 30912 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_327
timestamp 1649977179
transform 1 0 31188 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_339
timestamp 1649977179
transform 1 0 32292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_347
timestamp 1649977179
transform 1 0 33028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_350
timestamp 1649977179
transform 1 0 33304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1649977179
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_367
timestamp 1649977179
transform 1 0 34868 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_371
timestamp 1649977179
transform 1 0 35236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_374
timestamp 1649977179
transform 1 0 35512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_380
timestamp 1649977179
transform 1 0 36064 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_395
timestamp 1649977179
transform 1 0 37444 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1649977179
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_66
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1649977179
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1649977179
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1649977179
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_102
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_121
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_139
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_183
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_208
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_235
timestamp 1649977179
transform 1 0 22724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_246
timestamp 1649977179
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_256
timestamp 1649977179
transform 1 0 24656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_262
timestamp 1649977179
transform 1 0 25208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_268
timestamp 1649977179
transform 1 0 25760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1649977179
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp 1649977179
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1649977179
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_116
timestamp 1649977179
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_128
timestamp 1649977179
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_156
timestamp 1649977179
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_162
timestamp 1649977179
transform 1 0 16008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_201
timestamp 1649977179
transform 1 0 19596 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_208
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_226
timestamp 1649977179
transform 1 0 21896 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_234
timestamp 1649977179
transform 1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_239
timestamp 1649977179
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_259
timestamp 1649977179
transform 1 0 24932 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_271
timestamp 1649977179
transform 1 0 26036 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_283
timestamp 1649977179
transform 1 0 27140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_295
timestamp 1649977179
transform 1 0 28244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_60
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1649977179
transform 1 0 7912 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_80
timestamp 1649977179
transform 1 0 8464 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_92
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_97
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1649977179
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_172
timestamp 1649977179
transform 1 0 16928 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_180
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_188
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_200
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_208
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_231
timestamp 1649977179
transform 1 0 22356 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_243
timestamp 1649977179
transform 1 0 23460 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_255
timestamp 1649977179
transform 1 0 24564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_267
timestamp 1649977179
transform 1 0 25668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_76
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_89
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_103
timestamp 1649977179
transform 1 0 10580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_115
timestamp 1649977179
transform 1 0 11684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_126
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_146
timestamp 1649977179
transform 1 0 14536 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_158
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_170
timestamp 1649977179
transform 1 0 16744 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_182
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_203
timestamp 1649977179
transform 1 0 19780 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_207
timestamp 1649977179
transform 1 0 20148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_212
timestamp 1649977179
transform 1 0 20608 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_224
timestamp 1649977179
transform 1 0 21712 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_236
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1649977179
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1649977179
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_36
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1649977179
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_85
timestamp 1649977179
transform 1 0 8924 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_89
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_95
timestamp 1649977179
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_101
timestamp 1649977179
transform 1 0 10396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_121
timestamp 1649977179
transform 1 0 12236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_129
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_141
timestamp 1649977179
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_145
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_152
timestamp 1649977179
transform 1 0 15088 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_173
timestamp 1649977179
transform 1 0 17020 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_199
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_206
timestamp 1649977179
transform 1 0 20056 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_218
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_243
timestamp 1649977179
transform 1 0 23460 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_255
timestamp 1649977179
transform 1 0 24564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_267
timestamp 1649977179
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_43
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_51
timestamp 1649977179
transform 1 0 5796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_55
timestamp 1649977179
transform 1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_66
timestamp 1649977179
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_78
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_92
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_104
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_116
timestamp 1649977179
transform 1 0 11776 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_131
timestamp 1649977179
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_146
timestamp 1649977179
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1649977179
transform 1 0 15640 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_176
timestamp 1649977179
transform 1 0 17296 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_183
timestamp 1649977179
transform 1 0 17940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_212
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_234
timestamp 1649977179
transform 1 0 22632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1649977179
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1649977179
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_31
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_79
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1649977179
transform 1 0 9292 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_95
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_142
timestamp 1649977179
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1649977179
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_174
timestamp 1649977179
transform 1 0 17112 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_186
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_194
timestamp 1649977179
transform 1 0 18952 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_199
timestamp 1649977179
transform 1 0 19412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_203
timestamp 1649977179
transform 1 0 19780 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1649977179
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_57
timestamp 1649977179
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_71
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_92
timestamp 1649977179
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_111
timestamp 1649977179
transform 1 0 11316 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_118
timestamp 1649977179
transform 1 0 11960 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_149
timestamp 1649977179
transform 1 0 14812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_161
timestamp 1649977179
transform 1 0 15916 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1649977179
transform 1 0 16468 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1649977179
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1649977179
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_72
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_91
timestamp 1649977179
transform 1 0 9476 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1649977179
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_126
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_138
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_150
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_192
timestamp 1649977179
transform 1 0 18768 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_204
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1649977179
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_11
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_17
timestamp 1649977179
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_35
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_45
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_58
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_70
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_102
timestamp 1649977179
transform 1 0 10488 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_127
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_200
timestamp 1649977179
transform 1 0 19504 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_212
timestamp 1649977179
transform 1 0 20608 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_224
timestamp 1649977179
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_236
timestamp 1649977179
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1649977179
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_21
timestamp 1649977179
transform 1 0 3036 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_33
timestamp 1649977179
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_86
timestamp 1649977179
transform 1 0 9016 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_98
timestamp 1649977179
transform 1 0 10120 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_104
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_160
timestamp 1649977179
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_192
timestamp 1649977179
transform 1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_213
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_160
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_172
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_180
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_185
timestamp 1649977179
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_222
timestamp 1649977179
transform 1 0 21528 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_234
timestamp 1649977179
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_246
timestamp 1649977179
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_36
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_177
timestamp 1649977179
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1649977179
transform 1 0 18400 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1649977179
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1649977179
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1649977179
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1649977179
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_113
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_125
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_160
timestamp 1649977179
transform 1 0 15824 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_181
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1649977179
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_212
timestamp 1649977179
transform 1 0 20608 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_224
timestamp 1649977179
transform 1 0 21712 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_236
timestamp 1649977179
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_74
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_90
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1649977179
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1649977179
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_195
timestamp 1649977179
transform 1 0 19044 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_218
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_72
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_113
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_125
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1649977179
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_160
timestamp 1649977179
transform 1 0 15824 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_172
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_184
timestamp 1649977179
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_204
timestamp 1649977179
transform 1 0 19872 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_208
timestamp 1649977179
transform 1 0 20240 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_215
timestamp 1649977179
transform 1 0 20884 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_227
timestamp 1649977179
transform 1 0 21988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_239
timestamp 1649977179
transform 1 0 23092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_11
timestamp 1649977179
transform 1 0 2116 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_30
timestamp 1649977179
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_42
timestamp 1649977179
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_101
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_143
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1649977179
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_214
timestamp 1649977179
transform 1 0 20792 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_220
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_232
timestamp 1649977179
transform 1 0 22448 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1649977179
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_11
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_30
timestamp 1649977179
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_42
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1649977179
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_227
timestamp 1649977179
transform 1 0 21988 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_239
timestamp 1649977179
transform 1 0 23092 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_251
timestamp 1649977179
transform 1 0 24196 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_263
timestamp 1649977179
transform 1 0 25300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1649977179
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_35
timestamp 1649977179
transform 1 0 4324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_39
timestamp 1649977179
transform 1 0 4692 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_63
timestamp 1649977179
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_114
timestamp 1649977179
transform 1 0 11592 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_126
timestamp 1649977179
transform 1 0 12696 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_200
timestamp 1649977179
transform 1 0 19504 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_207
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_31
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_85
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_121
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_160
timestamp 1649977179
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1649977179
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1649977179
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1649977179
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_234
timestamp 1649977179
transform 1 0 22632 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_240
timestamp 1649977179
transform 1 0 23184 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_252
timestamp 1649977179
transform 1 0 24288 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_264
timestamp 1649977179
transform 1 0 25392 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1649977179
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_71
timestamp 1649977179
transform 1 0 7636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_105
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_117
timestamp 1649977179
transform 1 0 11868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1649977179
transform 1 0 15732 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_179
timestamp 1649977179
transform 1 0 17572 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_187
timestamp 1649977179
transform 1 0 18308 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1649977179
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_220
timestamp 1649977179
transform 1 0 21344 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1649977179
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_232
timestamp 1649977179
transform 1 0 22448 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1649977179
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_30
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1649977179
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_73
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_121
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1649977179
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1649977179
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_51
timestamp 1649977179
transform 1 0 5796 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_63
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1649977179
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_101
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_113
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_119
timestamp 1649977179
transform 1 0 12052 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_160
timestamp 1649977179
transform 1 0 15824 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_172
timestamp 1649977179
transform 1 0 16928 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_184
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_206
timestamp 1649977179
transform 1 0 20056 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_218
timestamp 1649977179
transform 1 0 21160 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_230
timestamp 1649977179
transform 1 0 22264 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_242
timestamp 1649977179
transform 1 0 23368 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1649977179
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_30
timestamp 1649977179
transform 1 0 3864 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_42
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_21
timestamp 1649977179
transform 1 0 3036 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_36
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_42
timestamp 1649977179
transform 1 0 4968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1649977179
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_58
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_62
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1649977179
transform 1 0 7912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1649977179
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_26
timestamp 1649977179
transform 1 0 3496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp 1649977179
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_63
timestamp 1649977179
transform 1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_70
timestamp 1649977179
transform 1 0 7544 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_80
timestamp 1649977179
transform 1 0 8464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_86
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_99
timestamp 1649977179
transform 1 0 10212 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_123
timestamp 1649977179
transform 1 0 12420 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_135
timestamp 1649977179
transform 1 0 13524 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_147
timestamp 1649977179
transform 1 0 14628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_171
timestamp 1649977179
transform 1 0 16836 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_183
timestamp 1649977179
transform 1 0 17940 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_195
timestamp 1649977179
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_207
timestamp 1649977179
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_21
timestamp 1649977179
transform 1 0 3036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1649977179
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_55
timestamp 1649977179
transform 1 0 6164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_61
timestamp 1649977179
transform 1 0 6716 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1649977179
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_89
timestamp 1649977179
transform 1 0 9292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_96
timestamp 1649977179
transform 1 0 9936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_103
timestamp 1649977179
transform 1 0 10580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_110
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_117
timestamp 1649977179
transform 1 0 11868 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1649977179
transform 1 0 12604 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_128
timestamp 1649977179
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_171
timestamp 1649977179
transform 1 0 16836 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1649977179
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_34
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_44
timestamp 1649977179
transform 1 0 5152 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_65
timestamp 1649977179
transform 1 0 7084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_76
timestamp 1649977179
transform 1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_89
timestamp 1649977179
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_95
timestamp 1649977179
transform 1 0 9844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_126
timestamp 1649977179
transform 1 0 12696 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_130
timestamp 1649977179
transform 1 0 13064 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_133
timestamp 1649977179
transform 1 0 13340 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_151
timestamp 1649977179
transform 1 0 14996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1649977179
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_187
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_199
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_211
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_33
timestamp 1649977179
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_36
timestamp 1649977179
transform 1 0 4416 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_48
timestamp 1649977179
transform 1 0 5520 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_60
timestamp 1649977179
transform 1 0 6624 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_74
timestamp 1649977179
transform 1 0 7912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1649977179
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp 1649977179
transform 1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_105
timestamp 1649977179
transform 1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_118
timestamp 1649977179
transform 1 0 11960 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1649977179
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_143
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1649977179
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_156
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_164
timestamp 1649977179
transform 1 0 16192 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1649977179
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_98
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1649977179
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_127
timestamp 1649977179
transform 1 0 12788 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_143
timestamp 1649977179
transform 1 0 14260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1649977179
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1649977179
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_184
timestamp 1649977179
transform 1 0 18032 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_196
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_208
timestamp 1649977179
transform 1 0 20240 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1649977179
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_117
timestamp 1649977179
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1649977179
transform 1 0 12604 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_128
timestamp 1649977179
transform 1 0 12880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1649977179
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_169
timestamp 1649977179
transform 1 0 16652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_181
timestamp 1649977179
transform 1 0 17756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1649977179
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1649977179
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1649977179
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_11
timestamp 1649977179
transform 1 0 2116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_23
timestamp 1649977179
transform 1 0 3220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_35
timestamp 1649977179
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1649977179
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_7
timestamp 1649977179
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_11
timestamp 1649977179
transform 1 0 2116 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_14
timestamp 1649977179
transform 1 0 2392 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 1649977179
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_395
timestamp 1649977179
transform 1 0 37444 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1649977179
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_7
timestamp 1649977179
transform 1 0 1748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_12
timestamp 1649977179
transform 1 0 2208 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_20
timestamp 1649977179
transform 1 0 2944 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_28
timestamp 1649977179
transform 1 0 3680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_32
timestamp 1649977179
transform 1 0 4048 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_40
timestamp 1649977179
transform 1 0 4784 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_44
timestamp 1649977179
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_59
timestamp 1649977179
transform 1 0 6532 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_65
timestamp 1649977179
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_68
timestamp 1649977179
transform 1 0 7360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_80
timestamp 1649977179
transform 1 0 8464 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_88
timestamp 1649977179
transform 1 0 9200 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_92
timestamp 1649977179
transform 1 0 9568 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_100
timestamp 1649977179
transform 1 0 10304 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_104
timestamp 1649977179
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_116
timestamp 1649977179
transform 1 0 11776 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_124
timestamp 1649977179
transform 1 0 12512 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_128
timestamp 1649977179
transform 1 0 12880 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_136
timestamp 1649977179
transform 1 0 13616 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_141
timestamp 1649977179
transform 1 0 14076 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_152
timestamp 1649977179
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1649977179
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_173
timestamp 1649977179
transform 1 0 17020 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_176
timestamp 1649977179
transform 1 0 17296 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_184
timestamp 1649977179
transform 1 0 18032 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_188
timestamp 1649977179
transform 1 0 18400 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_196
timestamp 1649977179
transform 1 0 19136 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_200
timestamp 1649977179
transform 1 0 19504 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_208
timestamp 1649977179
transform 1 0 20240 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_212
timestamp 1649977179
transform 1 0 20608 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_227
timestamp 1649977179
transform 1 0 21988 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_233
timestamp 1649977179
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_236
timestamp 1649977179
transform 1 0 22816 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_248
timestamp 1649977179
transform 1 0 23920 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_256
timestamp 1649977179
transform 1 0 24656 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_269
timestamp 1649977179
transform 1 0 25852 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1649977179
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_284
timestamp 1649977179
transform 1 0 27232 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_292
timestamp 1649977179
transform 1 0 27968 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_296
timestamp 1649977179
transform 1 0 28336 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_304
timestamp 1649977179
transform 1 0 29072 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_309
timestamp 1649977179
transform 1 0 29532 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_320
timestamp 1649977179
transform 1 0 30544 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1649977179
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_345
timestamp 1649977179
transform 1 0 32844 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_353
timestamp 1649977179
transform 1 0 33580 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_356
timestamp 1649977179
transform 1 0 33856 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_364
timestamp 1649977179
transform 1 0 34592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_368
timestamp 1649977179
transform 1 0 34960 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_376
timestamp 1649977179
transform 1 0 35696 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_380
timestamp 1649977179
transform 1 0 36064 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_395
timestamp 1649977179
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1649977179
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_13
timestamp 1649977179
transform 1 0 2300 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_19
timestamp 1649977179
transform 1 0 2852 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1649977179
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_35
timestamp 1649977179
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_43
timestamp 1649977179
transform 1 0 5060 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_47
timestamp 1649977179
transform 1 0 5428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1649977179
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_60
timestamp 1649977179
transform 1 0 6624 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_71
timestamp 1649977179
transform 1 0 7636 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1649977179
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_88
timestamp 1649977179
transform 1 0 9200 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_95
timestamp 1649977179
transform 1 0 9844 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_103
timestamp 1649977179
transform 1 0 10580 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_107
timestamp 1649977179
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1649977179
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1649977179
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_119
timestamp 1649977179
transform 1 0 12052 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_127
timestamp 1649977179
transform 1 0 12788 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_131
timestamp 1649977179
transform 1 0 13156 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_144
timestamp 1649977179
transform 1 0 14352 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_155
timestamp 1649977179
transform 1 0 15364 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_161
timestamp 1649977179
transform 1 0 15916 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_164
timestamp 1649977179
transform 1 0 16192 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_172
timestamp 1649977179
transform 1 0 16928 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_179
timestamp 1649977179
transform 1 0 17572 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_187
timestamp 1649977179
transform 1 0 18308 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_191
timestamp 1649977179
transform 1 0 18676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_203
timestamp 1649977179
transform 1 0 19780 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_211
timestamp 1649977179
transform 1 0 20516 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_215
timestamp 1649977179
transform 1 0 20884 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1649977179
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_229
timestamp 1649977179
transform 1 0 22172 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_235
timestamp 1649977179
transform 1 0 22724 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_240
timestamp 1649977179
transform 1 0 23184 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1649977179
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_257
timestamp 1649977179
transform 1 0 24748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_271
timestamp 1649977179
transform 1 0 26036 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1649977179
transform 1 0 26496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_281
timestamp 1649977179
transform 1 0 26956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_288
timestamp 1649977179
transform 1 0 27600 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_300
timestamp 1649977179
transform 1 0 28704 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_64_313
timestamp 1649977179
transform 1 0 29900 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_319
timestamp 1649977179
transform 1 0 30452 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_324
timestamp 1649977179
transform 1 0 30912 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_332
timestamp 1649977179
transform 1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_341
timestamp 1649977179
transform 1 0 32476 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_349
timestamp 1649977179
transform 1 0 33212 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_355
timestamp 1649977179
transform 1 0 33764 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1649977179
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_372
timestamp 1649977179
transform 1 0 35328 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_384
timestamp 1649977179
transform 1 0 36432 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_397
timestamp 1649977179
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1649977179
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _181_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _182_
timestamp 1649977179
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _183_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _184_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _185_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _186_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15088 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _187_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _188_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _189_
timestamp 1649977179
transform 1 0 15088 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _190_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1649977179
transform -1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _192_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9844 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _193_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_4  _194_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__a32o_1  _195_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _196_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10948 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _197_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12144 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _198_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _199_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _200_
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _201_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _202_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _203_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _204_
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _205_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _206_
timestamp 1649977179
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _207_
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _208_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _209_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _210_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _211_
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 1649977179
transform 1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _214_
timestamp 1649977179
transform 1 0 9384 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _215_
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _216_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12420 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 1649977179
transform -1 0 5796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _218_
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _219_
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _220_
timestamp 1649977179
transform -1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _221_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _222_
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _223_
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _224_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _225_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7176 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _227_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _228_
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _229_
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _230_
timestamp 1649977179
transform 1 0 2576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _231_
timestamp 1649977179
transform 1 0 4140 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp 1649977179
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _233_
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _234_
timestamp 1649977179
transform 1 0 4140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _235_
timestamp 1649977179
transform 1 0 7268 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp 1649977179
transform 1 0 6532 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _237_
timestamp 1649977179
transform 1 0 7268 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1649977179
transform 1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _239_
timestamp 1649977179
transform 1 0 8464 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1649977179
transform 1 0 7268 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _241_
timestamp 1649977179
transform 1 0 10212 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1649977179
transform 1 0 9844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _243_
timestamp 1649977179
transform 1 0 9936 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1649977179
transform -1 0 10212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _245_
timestamp 1649977179
transform 1 0 11868 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1649977179
transform 1 0 10304 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _247_
timestamp 1649977179
transform 1 0 12328 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1649977179
transform 1 0 11592 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1649977179
transform 1 0 12880 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1649977179
transform 1 0 10948 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1649977179
transform 1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _253_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1649977179
transform 1 0 15640 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1649977179
transform 1 0 16928 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _259_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7176 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _260_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _261_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14536 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _262_
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _263_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5520 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _264_
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1649977179
transform -1 0 6164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _267_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _268_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _269_
timestamp 1649977179
transform -1 0 6348 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _270_
timestamp 1649977179
transform -1 0 3128 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1649977179
transform 1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1649977179
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1649977179
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _274_
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _275_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _276_
timestamp 1649977179
transform 1 0 15456 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _278_
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _279_
timestamp 1649977179
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _280_
timestamp 1649977179
transform -1 0 18492 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _281_
timestamp 1649977179
transform 1 0 19228 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _282_
timestamp 1649977179
transform 1 0 19872 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _283_
timestamp 1649977179
transform 1 0 9936 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_4  _284_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__clkbuf_4  _285_
timestamp 1649977179
transform -1 0 20884 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _286_
timestamp 1649977179
transform 1 0 19320 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _288_
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _289_
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _290_
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _291_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _292_
timestamp 1649977179
transform 1 0 20516 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1649977179
transform 1 0 19872 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _294_
timestamp 1649977179
transform 1 0 23828 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _295_
timestamp 1649977179
transform 1 0 24104 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp 1649977179
transform 1 0 21712 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _298_
timestamp 1649977179
transform -1 0 23736 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _299_
timestamp 1649977179
transform 1 0 22356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _300_
timestamp 1649977179
transform 1 0 20516 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _302_
timestamp 1649977179
transform -1 0 23184 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _303_
timestamp 1649977179
transform 1 0 20976 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _304_
timestamp 1649977179
transform 1 0 20332 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _306_
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _307_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21160 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _309_
timestamp 1649977179
transform 1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _310_
timestamp 1649977179
transform -1 0 22448 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _311_
timestamp 1649977179
transform 1 0 20516 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _312_
timestamp 1649977179
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _313_
timestamp 1649977179
transform -1 0 22172 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _314_
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1649977179
transform 1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _316_
timestamp 1649977179
transform -1 0 23460 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _317_
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1649977179
transform 1 0 19320 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _319_
timestamp 1649977179
transform 1 0 19044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _320_
timestamp 1649977179
transform -1 0 22724 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _321_
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _322_
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _323_
timestamp 1649977179
transform 1 0 18032 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _324_
timestamp 1649977179
transform -1 0 20608 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _325_
timestamp 1649977179
transform -1 0 20240 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _327_
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _328_
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _329_
timestamp 1649977179
transform -1 0 18768 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _330_
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _331_
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _332_
timestamp 1649977179
transform -1 0 17756 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _333_
timestamp 1649977179
transform -1 0 17848 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _334_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _335_
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _336_
timestamp 1649977179
transform -1 0 17940 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _337_
timestamp 1649977179
transform -1 0 17848 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1649977179
transform 1 0 18768 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _339_
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _340_
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _341_
timestamp 1649977179
transform -1 0 19412 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1649977179
transform 1 0 19136 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _343_
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _344_
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _345_
timestamp 1649977179
transform -1 0 19780 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _346_
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _347_
timestamp 1649977179
transform 1 0 18768 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp 1649977179
transform 1 0 6716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1649977179
transform -1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _350_
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _351_
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _352_
timestamp 1649977179
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1649977179
transform 1 0 5612 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1649977179
transform 1 0 4416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_2  _355_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13156 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _356_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _357_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _358_
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _359_
timestamp 1649977179
transform 1 0 2392 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _360_
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _361_
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _362_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _363_
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _364_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9476 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _365_
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _366_
timestamp 1649977179
transform -1 0 10764 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _367_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _368_
timestamp 1649977179
transform 1 0 6992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _369_
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _370_
timestamp 1649977179
transform -1 0 6624 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _371_
timestamp 1649977179
transform 1 0 1840 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _372_
timestamp 1649977179
transform 1 0 2392 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _373_
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _374_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _377_
timestamp 1649977179
transform 1 0 6164 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp 1649977179
transform -1 0 10488 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp 1649977179
transform 1 0 9200 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp 1649977179
transform 1 0 9292 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp 1649977179
transform 1 0 8924 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _385_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _386_
timestamp 1649977179
transform 1 0 12512 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _387_
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _388_
timestamp 1649977179
transform 1 0 1840 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _389_
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _390_
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _391_
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _392_
timestamp 1649977179
transform 1 0 14352 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _393_
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _394_
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _395_
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _396_
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _397_
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _398_
timestamp 1649977179
transform 1 0 14352 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _399_
timestamp 1649977179
transform 1 0 16100 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _400_
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _401_
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _402_
timestamp 1649977179
transform 1 0 14260 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _403_
timestamp 1649977179
transform 1 0 14260 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _404_
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _405_
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _406_
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _407_
timestamp 1649977179
transform -1 0 3864 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _408_
timestamp 1649977179
transform 1 0 1840 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _409_
timestamp 1649977179
transform 1 0 1840 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _410_
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_clk opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_i_clk
timestamp 1649977179
transform -1 0 4416 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_i_clk
timestamp 1649977179
transform 1 0 5244 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_i_clk
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_i_clk
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1649977179
transform 1 0 1748 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1649977179
transform 1 0 2944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 4324 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 15088 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 16652 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 17296 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 18400 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 19504 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 20608 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 5152 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 6348 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 7360 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 9568 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 10672 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 11776 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 12880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2392 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 4140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 16192 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 5428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform 1 0 33396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform 1 0 34408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform 1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 35972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform 1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 30176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform 1 0 30544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform 1 0 31188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform 1 0 32752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform 1 0 36064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform 1 0 36616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1649977179
transform -1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 2208 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 33856 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 34960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 36064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 37260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 23184 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 25116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 26128 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 27232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 28336 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 30544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 37812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 25484 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal2 s 662 39200 718 40000 0 FreeSans 224 90 0 0 cw_ack
port 0 nsew signal input
flabel metal2 s 1766 39200 1822 40000 0 FreeSans 224 90 0 0 cw_dir
port 1 nsew signal tristate
flabel metal2 s 2870 39200 2926 40000 0 FreeSans 224 90 0 0 cw_err
port 2 nsew signal input
flabel metal2 s 3974 39200 4030 40000 0 FreeSans 224 90 0 0 cw_io_i[0]
port 3 nsew signal input
flabel metal2 s 15014 39200 15070 40000 0 FreeSans 224 90 0 0 cw_io_i[10]
port 4 nsew signal input
flabel metal2 s 16118 39200 16174 40000 0 FreeSans 224 90 0 0 cw_io_i[11]
port 5 nsew signal input
flabel metal2 s 17222 39200 17278 40000 0 FreeSans 224 90 0 0 cw_io_i[12]
port 6 nsew signal input
flabel metal2 s 18326 39200 18382 40000 0 FreeSans 224 90 0 0 cw_io_i[13]
port 7 nsew signal input
flabel metal2 s 19430 39200 19486 40000 0 FreeSans 224 90 0 0 cw_io_i[14]
port 8 nsew signal input
flabel metal2 s 20534 39200 20590 40000 0 FreeSans 224 90 0 0 cw_io_i[15]
port 9 nsew signal input
flabel metal2 s 5078 39200 5134 40000 0 FreeSans 224 90 0 0 cw_io_i[1]
port 10 nsew signal input
flabel metal2 s 6182 39200 6238 40000 0 FreeSans 224 90 0 0 cw_io_i[2]
port 11 nsew signal input
flabel metal2 s 7286 39200 7342 40000 0 FreeSans 224 90 0 0 cw_io_i[3]
port 12 nsew signal input
flabel metal2 s 8390 39200 8446 40000 0 FreeSans 224 90 0 0 cw_io_i[4]
port 13 nsew signal input
flabel metal2 s 9494 39200 9550 40000 0 FreeSans 224 90 0 0 cw_io_i[5]
port 14 nsew signal input
flabel metal2 s 10598 39200 10654 40000 0 FreeSans 224 90 0 0 cw_io_i[6]
port 15 nsew signal input
flabel metal2 s 11702 39200 11758 40000 0 FreeSans 224 90 0 0 cw_io_i[7]
port 16 nsew signal input
flabel metal2 s 12806 39200 12862 40000 0 FreeSans 224 90 0 0 cw_io_i[8]
port 17 nsew signal input
flabel metal2 s 13910 39200 13966 40000 0 FreeSans 224 90 0 0 cw_io_i[9]
port 18 nsew signal input
flabel metal2 s 21638 39200 21694 40000 0 FreeSans 224 90 0 0 cw_io_o[0]
port 19 nsew signal tristate
flabel metal2 s 32678 39200 32734 40000 0 FreeSans 224 90 0 0 cw_io_o[10]
port 20 nsew signal tristate
flabel metal2 s 33782 39200 33838 40000 0 FreeSans 224 90 0 0 cw_io_o[11]
port 21 nsew signal tristate
flabel metal2 s 34886 39200 34942 40000 0 FreeSans 224 90 0 0 cw_io_o[12]
port 22 nsew signal tristate
flabel metal2 s 35990 39200 36046 40000 0 FreeSans 224 90 0 0 cw_io_o[13]
port 23 nsew signal tristate
flabel metal2 s 37094 39200 37150 40000 0 FreeSans 224 90 0 0 cw_io_o[14]
port 24 nsew signal tristate
flabel metal2 s 38198 39200 38254 40000 0 FreeSans 224 90 0 0 cw_io_o[15]
port 25 nsew signal tristate
flabel metal2 s 22742 39200 22798 40000 0 FreeSans 224 90 0 0 cw_io_o[1]
port 26 nsew signal tristate
flabel metal2 s 23846 39200 23902 40000 0 FreeSans 224 90 0 0 cw_io_o[2]
port 27 nsew signal tristate
flabel metal2 s 24950 39200 25006 40000 0 FreeSans 224 90 0 0 cw_io_o[3]
port 28 nsew signal tristate
flabel metal2 s 26054 39200 26110 40000 0 FreeSans 224 90 0 0 cw_io_o[4]
port 29 nsew signal tristate
flabel metal2 s 27158 39200 27214 40000 0 FreeSans 224 90 0 0 cw_io_o[5]
port 30 nsew signal tristate
flabel metal2 s 28262 39200 28318 40000 0 FreeSans 224 90 0 0 cw_io_o[6]
port 31 nsew signal tristate
flabel metal2 s 29366 39200 29422 40000 0 FreeSans 224 90 0 0 cw_io_o[7]
port 32 nsew signal tristate
flabel metal2 s 30470 39200 30526 40000 0 FreeSans 224 90 0 0 cw_io_o[8]
port 33 nsew signal tristate
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 cw_io_o[9]
port 34 nsew signal tristate
flabel metal2 s 39302 39200 39358 40000 0 FreeSans 224 90 0 0 cw_req
port 35 nsew signal tristate
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 i_clk
port 36 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 i_rst
port 37 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 38 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 38 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 39 nsew ground bidirectional
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 wb_4_burst
port 40 nsew signal input
flabel metal2 s 2870 0 2926 800 0 FreeSans 224 90 0 0 wb_8_burst
port 41 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 wb_ack
port 42 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 wb_adr[0]
port 43 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wb_adr[10]
port 44 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wb_adr[11]
port 45 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wb_adr[12]
port 46 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wb_adr[13]
port 47 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wb_adr[14]
port 48 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wb_adr[15]
port 49 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wb_adr[16]
port 50 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wb_adr[17]
port 51 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wb_adr[18]
port 52 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wb_adr[19]
port 53 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wb_adr[1]
port 54 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wb_adr[20]
port 55 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wb_adr[21]
port 56 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wb_adr[22]
port 57 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wb_adr[23]
port 58 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 wb_adr[2]
port 59 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wb_adr[3]
port 60 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wb_adr[4]
port 61 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wb_adr[5]
port 62 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wb_adr[6]
port 63 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wb_adr[7]
port 64 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wb_adr[8]
port 65 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wb_adr[9]
port 66 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wb_cyc
port 67 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 wb_err
port 68 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wb_i_dat[0]
port 69 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 wb_i_dat[10]
port 70 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 wb_i_dat[11]
port 71 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 wb_i_dat[12]
port 72 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 wb_i_dat[13]
port 73 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 wb_i_dat[14]
port 74 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 wb_i_dat[15]
port 75 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 wb_i_dat[1]
port 76 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wb_i_dat[2]
port 77 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 wb_i_dat[3]
port 78 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 wb_i_dat[4]
port 79 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 wb_i_dat[5]
port 80 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 wb_i_dat[6]
port 81 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 wb_i_dat[7]
port 82 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 wb_i_dat[8]
port 83 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 wb_i_dat[9]
port 84 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 wb_o_dat[0]
port 85 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 wb_o_dat[10]
port 86 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 wb_o_dat[11]
port 87 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 wb_o_dat[12]
port 88 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 wb_o_dat[13]
port 89 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 wb_o_dat[14]
port 90 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 wb_o_dat[15]
port 91 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 wb_o_dat[1]
port 92 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 wb_o_dat[2]
port 93 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 wb_o_dat[3]
port 94 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 wb_o_dat[4]
port 95 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 wb_o_dat[5]
port 96 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 wb_o_dat[6]
port 97 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 wb_o_dat[7]
port 98 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 wb_o_dat[8]
port 99 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 wb_o_dat[9]
port 100 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 wb_sel[0]
port 101 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 wb_sel[1]
port 102 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 wb_stb
port 103 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 wb_we
port 104 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
