magic
tech sky130B
magscale 1 2
timestamp 1663051598
<< obsli1 >>
rect 1104 2159 48852 47345
<< obsm1 >>
rect 14 1776 49666 47524
<< metal2 >>
rect 662 49200 718 50000
rect 1950 49200 2006 50000
rect 3238 49200 3294 50000
rect 5170 49200 5226 50000
rect 6458 49200 6514 50000
rect 7746 49200 7802 50000
rect 9034 49200 9090 50000
rect 10322 49200 10378 50000
rect 12254 49200 12310 50000
rect 13542 49200 13598 50000
rect 14830 49200 14886 50000
rect 16118 49200 16174 50000
rect 18050 49200 18106 50000
rect 19338 49200 19394 50000
rect 20626 49200 20682 50000
rect 21914 49200 21970 50000
rect 23202 49200 23258 50000
rect 25134 49200 25190 50000
rect 26422 49200 26478 50000
rect 27710 49200 27766 50000
rect 28998 49200 29054 50000
rect 30930 49200 30986 50000
rect 32218 49200 32274 50000
rect 33506 49200 33562 50000
rect 34794 49200 34850 50000
rect 36082 49200 36138 50000
rect 38014 49200 38070 50000
rect 39302 49200 39358 50000
rect 40590 49200 40646 50000
rect 41878 49200 41934 50000
rect 43810 49200 43866 50000
rect 45098 49200 45154 50000
rect 46386 49200 46442 50000
rect 47674 49200 47730 50000
rect 48962 49200 49018 50000
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36726 0 36782 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 49606 0 49662 800
<< obsm2 >>
rect 20 49144 606 49745
rect 774 49144 1894 49745
rect 2062 49144 3182 49745
rect 3350 49144 5114 49745
rect 5282 49144 6402 49745
rect 6570 49144 7690 49745
rect 7858 49144 8978 49745
rect 9146 49144 10266 49745
rect 10434 49144 12198 49745
rect 12366 49144 13486 49745
rect 13654 49144 14774 49745
rect 14942 49144 16062 49745
rect 16230 49144 17994 49745
rect 18162 49144 19282 49745
rect 19450 49144 20570 49745
rect 20738 49144 21858 49745
rect 22026 49144 23146 49745
rect 23314 49144 25078 49745
rect 25246 49144 26366 49745
rect 26534 49144 27654 49745
rect 27822 49144 28942 49745
rect 29110 49144 30874 49745
rect 31042 49144 32162 49745
rect 32330 49144 33450 49745
rect 33618 49144 34738 49745
rect 34906 49144 36026 49745
rect 36194 49144 37958 49745
rect 38126 49144 39246 49745
rect 39414 49144 40534 49745
rect 40702 49144 41822 49745
rect 41990 49144 43754 49745
rect 43922 49144 45042 49745
rect 45210 49144 46330 49745
rect 46498 49144 47618 49745
rect 47786 49144 48906 49745
rect 49074 49144 49660 49745
rect 20 856 49660 49144
rect 130 711 1250 856
rect 1418 711 2538 856
rect 2706 711 3826 856
rect 3994 711 5114 856
rect 5282 711 7046 856
rect 7214 711 8334 856
rect 8502 711 9622 856
rect 9790 711 10910 856
rect 11078 711 12198 856
rect 12366 711 14130 856
rect 14298 711 15418 856
rect 15586 711 16706 856
rect 16874 711 17994 856
rect 18162 711 19926 856
rect 20094 711 21214 856
rect 21382 711 22502 856
rect 22670 711 23790 856
rect 23958 711 25078 856
rect 25246 711 27010 856
rect 27178 711 28298 856
rect 28466 711 29586 856
rect 29754 711 30874 856
rect 31042 711 32806 856
rect 32974 711 34094 856
rect 34262 711 35382 856
rect 35550 711 36670 856
rect 36838 711 37958 856
rect 38126 711 39890 856
rect 40058 711 41178 856
rect 41346 711 42466 856
rect 42634 711 43754 856
rect 43922 711 45686 856
rect 45854 711 46974 856
rect 47142 711 48262 856
rect 48430 711 49550 856
<< metal3 >>
rect 0 49648 800 49768
rect 49200 48968 50000 49088
rect 0 48288 800 48408
rect 49200 47608 50000 47728
rect 0 46248 800 46368
rect 49200 46248 50000 46368
rect 0 44888 800 45008
rect 49200 44888 50000 45008
rect 0 43528 800 43648
rect 49200 43528 50000 43648
rect 0 42168 800 42288
rect 49200 41488 50000 41608
rect 0 40128 800 40248
rect 49200 40128 50000 40248
rect 0 38768 800 38888
rect 49200 38768 50000 38888
rect 0 37408 800 37528
rect 49200 37408 50000 37528
rect 0 36048 800 36168
rect 49200 35368 50000 35488
rect 0 34688 800 34808
rect 49200 34008 50000 34128
rect 0 32648 800 32768
rect 49200 32648 50000 32768
rect 0 31288 800 31408
rect 49200 31288 50000 31408
rect 0 29928 800 30048
rect 49200 29928 50000 30048
rect 0 28568 800 28688
rect 49200 27888 50000 28008
rect 0 26528 800 26648
rect 49200 26528 50000 26648
rect 0 25168 800 25288
rect 49200 25168 50000 25288
rect 0 23808 800 23928
rect 49200 23808 50000 23928
rect 0 22448 800 22568
rect 49200 21768 50000 21888
rect 0 21088 800 21208
rect 49200 20408 50000 20528
rect 0 19048 800 19168
rect 49200 19048 50000 19168
rect 0 17688 800 17808
rect 49200 17688 50000 17808
rect 0 16328 800 16448
rect 49200 16328 50000 16448
rect 0 14968 800 15088
rect 49200 14288 50000 14408
rect 0 12928 800 13048
rect 49200 12928 50000 13048
rect 0 11568 800 11688
rect 49200 11568 50000 11688
rect 0 10208 800 10328
rect 49200 10208 50000 10328
rect 0 8848 800 8968
rect 49200 8168 50000 8288
rect 0 7488 800 7608
rect 49200 6808 50000 6928
rect 0 5448 800 5568
rect 49200 5448 50000 5568
rect 0 4088 800 4208
rect 49200 4088 50000 4208
rect 0 2728 800 2848
rect 49200 2728 50000 2848
rect 0 1368 800 1488
rect 49200 688 50000 808
<< obsm3 >>
rect 880 49568 49200 49741
rect 800 49168 49200 49568
rect 800 48888 49120 49168
rect 800 48488 49200 48888
rect 880 48208 49200 48488
rect 800 47808 49200 48208
rect 800 47528 49120 47808
rect 800 46448 49200 47528
rect 880 46168 49120 46448
rect 800 45088 49200 46168
rect 880 44808 49120 45088
rect 800 43728 49200 44808
rect 880 43448 49120 43728
rect 800 42368 49200 43448
rect 880 42088 49200 42368
rect 800 41688 49200 42088
rect 800 41408 49120 41688
rect 800 40328 49200 41408
rect 880 40048 49120 40328
rect 800 38968 49200 40048
rect 880 38688 49120 38968
rect 800 37608 49200 38688
rect 880 37328 49120 37608
rect 800 36248 49200 37328
rect 880 35968 49200 36248
rect 800 35568 49200 35968
rect 800 35288 49120 35568
rect 800 34888 49200 35288
rect 880 34608 49200 34888
rect 800 34208 49200 34608
rect 800 33928 49120 34208
rect 800 32848 49200 33928
rect 880 32568 49120 32848
rect 800 31488 49200 32568
rect 880 31208 49120 31488
rect 800 30128 49200 31208
rect 880 29848 49120 30128
rect 800 28768 49200 29848
rect 880 28488 49200 28768
rect 800 28088 49200 28488
rect 800 27808 49120 28088
rect 800 26728 49200 27808
rect 880 26448 49120 26728
rect 800 25368 49200 26448
rect 880 25088 49120 25368
rect 800 24008 49200 25088
rect 880 23728 49120 24008
rect 800 22648 49200 23728
rect 880 22368 49200 22648
rect 800 21968 49200 22368
rect 800 21688 49120 21968
rect 800 21288 49200 21688
rect 880 21008 49200 21288
rect 800 20608 49200 21008
rect 800 20328 49120 20608
rect 800 19248 49200 20328
rect 880 18968 49120 19248
rect 800 17888 49200 18968
rect 880 17608 49120 17888
rect 800 16528 49200 17608
rect 880 16248 49120 16528
rect 800 15168 49200 16248
rect 880 14888 49200 15168
rect 800 14488 49200 14888
rect 800 14208 49120 14488
rect 800 13128 49200 14208
rect 880 12848 49120 13128
rect 800 11768 49200 12848
rect 880 11488 49120 11768
rect 800 10408 49200 11488
rect 880 10128 49120 10408
rect 800 9048 49200 10128
rect 880 8768 49200 9048
rect 800 8368 49200 8768
rect 800 8088 49120 8368
rect 800 7688 49200 8088
rect 880 7408 49200 7688
rect 800 7008 49200 7408
rect 800 6728 49120 7008
rect 800 5648 49200 6728
rect 880 5368 49120 5648
rect 800 4288 49200 5368
rect 880 4008 49120 4288
rect 800 2928 49200 4008
rect 880 2648 49120 2928
rect 800 1568 49200 2648
rect 880 1288 49200 1568
rect 800 888 49200 1288
rect 800 715 49120 888
<< metal4 >>
rect 4208 2128 4528 47376
rect 19568 2128 19888 47376
rect 34928 2128 35248 47376
<< obsm4 >>
rect 4659 2347 19488 47021
rect 19968 2347 34848 47021
rect 35328 2347 48149 47021
<< labels >>
rlabel metal3 s 0 28568 800 28688 6 cc_data_page
port 1 nsew signal input
rlabel metal2 s 7746 49200 7802 50000 6 cc_instr_page
port 2 nsew signal input
rlabel metal3 s 49200 34008 50000 34128 6 data_cacheable
port 3 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 data_mem_addr[0]
port 4 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 data_mem_addr[10]
port 5 nsew signal input
rlabel metal2 s 34794 49200 34850 50000 6 data_mem_addr[11]
port 6 nsew signal input
rlabel metal2 s 28998 49200 29054 50000 6 data_mem_addr[12]
port 7 nsew signal input
rlabel metal2 s 26422 49200 26478 50000 6 data_mem_addr[13]
port 8 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 data_mem_addr[14]
port 9 nsew signal input
rlabel metal2 s 40590 49200 40646 50000 6 data_mem_addr[15]
port 10 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 data_mem_addr[1]
port 11 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 data_mem_addr[2]
port 12 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 data_mem_addr[3]
port 13 nsew signal input
rlabel metal2 s 47674 49200 47730 50000 6 data_mem_addr[4]
port 14 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 data_mem_addr[5]
port 15 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 data_mem_addr[6]
port 16 nsew signal input
rlabel metal2 s 5170 49200 5226 50000 6 data_mem_addr[7]
port 17 nsew signal input
rlabel metal2 s 43810 49200 43866 50000 6 data_mem_addr[8]
port 18 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 data_mem_addr[9]
port 19 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 data_mem_addr_paged[0]
port 20 nsew signal output
rlabel metal2 s 46386 49200 46442 50000 6 data_mem_addr_paged[10]
port 21 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 data_mem_addr_paged[11]
port 22 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 data_mem_addr_paged[12]
port 23 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 data_mem_addr_paged[13]
port 24 nsew signal output
rlabel metal2 s 6458 49200 6514 50000 6 data_mem_addr_paged[14]
port 25 nsew signal output
rlabel metal3 s 49200 37408 50000 37528 6 data_mem_addr_paged[15]
port 26 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 data_mem_addr_paged[16]
port 27 nsew signal output
rlabel metal2 s 18050 49200 18106 50000 6 data_mem_addr_paged[17]
port 28 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 data_mem_addr_paged[18]
port 29 nsew signal output
rlabel metal3 s 49200 688 50000 808 6 data_mem_addr_paged[19]
port 30 nsew signal output
rlabel metal3 s 49200 14288 50000 14408 6 data_mem_addr_paged[1]
port 31 nsew signal output
rlabel metal3 s 49200 19048 50000 19168 6 data_mem_addr_paged[20]
port 32 nsew signal output
rlabel metal3 s 49200 21768 50000 21888 6 data_mem_addr_paged[21]
port 33 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 data_mem_addr_paged[22]
port 34 nsew signal output
rlabel metal2 s 25134 49200 25190 50000 6 data_mem_addr_paged[23]
port 35 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 data_mem_addr_paged[2]
port 36 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 data_mem_addr_paged[3]
port 37 nsew signal output
rlabel metal3 s 49200 25168 50000 25288 6 data_mem_addr_paged[4]
port 38 nsew signal output
rlabel metal2 s 23202 49200 23258 50000 6 data_mem_addr_paged[5]
port 39 nsew signal output
rlabel metal2 s 21914 49200 21970 50000 6 data_mem_addr_paged[6]
port 40 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 data_mem_addr_paged[7]
port 41 nsew signal output
rlabel metal2 s 32218 49200 32274 50000 6 data_mem_addr_paged[8]
port 42 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 data_mem_addr_paged[9]
port 43 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 fetch_wb_adr[0]
port 44 nsew signal input
rlabel metal2 s 10322 49200 10378 50000 6 fetch_wb_adr[10]
port 45 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 fetch_wb_adr[11]
port 46 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 fetch_wb_adr[12]
port 47 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 fetch_wb_adr[13]
port 48 nsew signal input
rlabel metal2 s 41878 49200 41934 50000 6 fetch_wb_adr[14]
port 49 nsew signal input
rlabel metal3 s 49200 43528 50000 43648 6 fetch_wb_adr[15]
port 50 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 fetch_wb_adr[1]
port 51 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 fetch_wb_adr[2]
port 52 nsew signal input
rlabel metal2 s 662 49200 718 50000 6 fetch_wb_adr[3]
port 53 nsew signal input
rlabel metal3 s 49200 12928 50000 13048 6 fetch_wb_adr[4]
port 54 nsew signal input
rlabel metal2 s 16118 49200 16174 50000 6 fetch_wb_adr[5]
port 55 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 fetch_wb_adr[6]
port 56 nsew signal input
rlabel metal3 s 49200 40128 50000 40248 6 fetch_wb_adr[7]
port 57 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 fetch_wb_adr[8]
port 58 nsew signal input
rlabel metal2 s 48962 49200 49018 50000 6 fetch_wb_adr[9]
port 59 nsew signal input
rlabel metal3 s 49200 38768 50000 38888 6 fetch_wb_adr_paged[0]
port 60 nsew signal output
rlabel metal3 s 49200 8168 50000 8288 6 fetch_wb_adr_paged[10]
port 61 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 fetch_wb_adr_paged[11]
port 62 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 fetch_wb_adr_paged[12]
port 63 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 fetch_wb_adr_paged[13]
port 64 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 fetch_wb_adr_paged[14]
port 65 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 fetch_wb_adr_paged[15]
port 66 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 fetch_wb_adr_paged[16]
port 67 nsew signal output
rlabel metal2 s 12254 49200 12310 50000 6 fetch_wb_adr_paged[17]
port 68 nsew signal output
rlabel metal3 s 49200 46248 50000 46368 6 fetch_wb_adr_paged[18]
port 69 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 fetch_wb_adr_paged[19]
port 70 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 fetch_wb_adr_paged[1]
port 71 nsew signal output
rlabel metal2 s 3238 49200 3294 50000 6 fetch_wb_adr_paged[20]
port 72 nsew signal output
rlabel metal2 s 14830 49200 14886 50000 6 fetch_wb_adr_paged[21]
port 73 nsew signal output
rlabel metal2 s 19338 49200 19394 50000 6 fetch_wb_adr_paged[22]
port 74 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 fetch_wb_adr_paged[23]
port 75 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 fetch_wb_adr_paged[2]
port 76 nsew signal output
rlabel metal3 s 49200 16328 50000 16448 6 fetch_wb_adr_paged[3]
port 77 nsew signal output
rlabel metal3 s 49200 47608 50000 47728 6 fetch_wb_adr_paged[4]
port 78 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 fetch_wb_adr_paged[5]
port 79 nsew signal output
rlabel metal3 s 49200 2728 50000 2848 6 fetch_wb_adr_paged[6]
port 80 nsew signal output
rlabel metal3 s 49200 17688 50000 17808 6 fetch_wb_adr_paged[7]
port 81 nsew signal output
rlabel metal2 s 33506 49200 33562 50000 6 fetch_wb_adr_paged[8]
port 82 nsew signal output
rlabel metal3 s 49200 10208 50000 10328 6 fetch_wb_adr_paged[9]
port 83 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 fetch_wb_o_dat[0]
port 84 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 fetch_wb_o_dat[10]
port 85 nsew signal output
rlabel metal3 s 49200 26528 50000 26648 6 fetch_wb_o_dat[11]
port 86 nsew signal output
rlabel metal3 s 49200 48968 50000 49088 6 fetch_wb_o_dat[12]
port 87 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 fetch_wb_o_dat[13]
port 88 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 fetch_wb_o_dat[14]
port 89 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 fetch_wb_o_dat[15]
port 90 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 fetch_wb_o_dat[1]
port 91 nsew signal output
rlabel metal2 s 20626 49200 20682 50000 6 fetch_wb_o_dat[2]
port 92 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 fetch_wb_o_dat[3]
port 93 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 fetch_wb_o_dat[4]
port 94 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 fetch_wb_o_dat[5]
port 95 nsew signal output
rlabel metal3 s 49200 4088 50000 4208 6 fetch_wb_o_dat[6]
port 96 nsew signal output
rlabel metal3 s 49200 35368 50000 35488 6 fetch_wb_o_dat[7]
port 97 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 fetch_wb_o_dat[8]
port 98 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 fetch_wb_o_dat[9]
port 99 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 i_clk
port 100 nsew signal input
rlabel metal3 s 49200 11568 50000 11688 6 i_rst
port 101 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 sr_bus_addr[0]
port 102 nsew signal input
rlabel metal3 s 49200 27888 50000 28008 6 sr_bus_addr[10]
port 103 nsew signal input
rlabel metal3 s 49200 41488 50000 41608 6 sr_bus_addr[11]
port 104 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 sr_bus_addr[12]
port 105 nsew signal input
rlabel metal3 s 49200 44888 50000 45008 6 sr_bus_addr[13]
port 106 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 sr_bus_addr[14]
port 107 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 sr_bus_addr[15]
port 108 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 sr_bus_addr[1]
port 109 nsew signal input
rlabel metal2 s 18 0 74 800 6 sr_bus_addr[2]
port 110 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 sr_bus_addr[3]
port 111 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 sr_bus_addr[4]
port 112 nsew signal input
rlabel metal2 s 13542 49200 13598 50000 6 sr_bus_addr[5]
port 113 nsew signal input
rlabel metal2 s 30930 49200 30986 50000 6 sr_bus_addr[6]
port 114 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 sr_bus_addr[7]
port 115 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 sr_bus_addr[8]
port 116 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 sr_bus_addr[9]
port 117 nsew signal input
rlabel metal2 s 39302 49200 39358 50000 6 sr_bus_data_o[0]
port 118 nsew signal input
rlabel metal2 s 27710 49200 27766 50000 6 sr_bus_data_o[10]
port 119 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 sr_bus_data_o[11]
port 120 nsew signal input
rlabel metal2 s 45098 49200 45154 50000 6 sr_bus_data_o[12]
port 121 nsew signal input
rlabel metal3 s 49200 6808 50000 6928 6 sr_bus_data_o[13]
port 122 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 sr_bus_data_o[14]
port 123 nsew signal input
rlabel metal3 s 49200 31288 50000 31408 6 sr_bus_data_o[15]
port 124 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 sr_bus_data_o[1]
port 125 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 sr_bus_data_o[2]
port 126 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 sr_bus_data_o[3]
port 127 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 sr_bus_data_o[4]
port 128 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 sr_bus_data_o[5]
port 129 nsew signal input
rlabel metal2 s 38014 49200 38070 50000 6 sr_bus_data_o[6]
port 130 nsew signal input
rlabel metal2 s 36082 49200 36138 50000 6 sr_bus_data_o[7]
port 131 nsew signal input
rlabel metal2 s 1950 49200 2006 50000 6 sr_bus_data_o[8]
port 132 nsew signal input
rlabel metal2 s 9034 49200 9090 50000 6 sr_bus_data_o[9]
port 133 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 sr_bus_we
port 134 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 135 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 135 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 136 nsew ground bidirectional
rlabel metal3 s 0 12928 800 13048 6 wb0_8_burst
port 137 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 wb1_4_burst
port 138 nsew signal output
rlabel metal3 s 49200 23808 50000 23928 6 wb1_8_burst
port 139 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 50000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5939022
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/upper_core_logic/runs/22_09_13_08_44/results/signoff/upper_core_logic.magic.gds
string GDS_START 333974
<< end >>

