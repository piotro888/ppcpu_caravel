magic
tech sky130A
magscale 1 2
timestamp 1672257255
<< obsli1 >>
rect 1104 2159 78844 157777
<< obsm1 >>
rect 750 1912 79658 157808
<< metal2 >>
rect 754 0 810 800
rect 1858 0 1914 800
rect 2962 0 3018 800
rect 4066 0 4122 800
rect 5170 0 5226 800
rect 6274 0 6330 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10690 0 10746 800
rect 11794 0 11850 800
rect 12898 0 12954 800
rect 14002 0 14058 800
rect 15106 0 15162 800
rect 16210 0 16266 800
rect 17314 0 17370 800
rect 18418 0 18474 800
rect 19522 0 19578 800
rect 20626 0 20682 800
rect 21730 0 21786 800
rect 22834 0 22890 800
rect 23938 0 23994 800
rect 25042 0 25098 800
rect 26146 0 26202 800
rect 27250 0 27306 800
rect 28354 0 28410 800
rect 29458 0 29514 800
rect 30562 0 30618 800
rect 31666 0 31722 800
rect 32770 0 32826 800
rect 33874 0 33930 800
rect 34978 0 35034 800
rect 36082 0 36138 800
rect 37186 0 37242 800
rect 38290 0 38346 800
rect 39394 0 39450 800
rect 40498 0 40554 800
rect 41602 0 41658 800
rect 42706 0 42762 800
rect 43810 0 43866 800
rect 44914 0 44970 800
rect 46018 0 46074 800
rect 47122 0 47178 800
rect 48226 0 48282 800
rect 49330 0 49386 800
rect 50434 0 50490 800
rect 51538 0 51594 800
rect 52642 0 52698 800
rect 53746 0 53802 800
rect 54850 0 54906 800
rect 55954 0 56010 800
rect 57058 0 57114 800
rect 58162 0 58218 800
rect 59266 0 59322 800
rect 60370 0 60426 800
rect 61474 0 61530 800
rect 62578 0 62634 800
rect 63682 0 63738 800
rect 64786 0 64842 800
rect 65890 0 65946 800
rect 66994 0 67050 800
rect 68098 0 68154 800
rect 69202 0 69258 800
rect 70306 0 70362 800
rect 71410 0 71466 800
rect 72514 0 72570 800
rect 73618 0 73674 800
rect 74722 0 74778 800
rect 75826 0 75882 800
rect 76930 0 76986 800
rect 78034 0 78090 800
rect 79138 0 79194 800
<< obsm2 >>
rect 756 856 79652 157797
rect 866 800 1802 856
rect 1970 800 2906 856
rect 3074 800 4010 856
rect 4178 800 5114 856
rect 5282 800 6218 856
rect 6386 800 7322 856
rect 7490 800 8426 856
rect 8594 800 9530 856
rect 9698 800 10634 856
rect 10802 800 11738 856
rect 11906 800 12842 856
rect 13010 800 13946 856
rect 14114 800 15050 856
rect 15218 800 16154 856
rect 16322 800 17258 856
rect 17426 800 18362 856
rect 18530 800 19466 856
rect 19634 800 20570 856
rect 20738 800 21674 856
rect 21842 800 22778 856
rect 22946 800 23882 856
rect 24050 800 24986 856
rect 25154 800 26090 856
rect 26258 800 27194 856
rect 27362 800 28298 856
rect 28466 800 29402 856
rect 29570 800 30506 856
rect 30674 800 31610 856
rect 31778 800 32714 856
rect 32882 800 33818 856
rect 33986 800 34922 856
rect 35090 800 36026 856
rect 36194 800 37130 856
rect 37298 800 38234 856
rect 38402 800 39338 856
rect 39506 800 40442 856
rect 40610 800 41546 856
rect 41714 800 42650 856
rect 42818 800 43754 856
rect 43922 800 44858 856
rect 45026 800 45962 856
rect 46130 800 47066 856
rect 47234 800 48170 856
rect 48338 800 49274 856
rect 49442 800 50378 856
rect 50546 800 51482 856
rect 51650 800 52586 856
rect 52754 800 53690 856
rect 53858 800 54794 856
rect 54962 800 55898 856
rect 56066 800 57002 856
rect 57170 800 58106 856
rect 58274 800 59210 856
rect 59378 800 60314 856
rect 60482 800 61418 856
rect 61586 800 62522 856
rect 62690 800 63626 856
rect 63794 800 64730 856
rect 64898 800 65834 856
rect 66002 800 66938 856
rect 67106 800 68042 856
rect 68210 800 69146 856
rect 69314 800 70250 856
rect 70418 800 71354 856
rect 71522 800 72458 856
rect 72626 800 73562 856
rect 73730 800 74666 856
rect 74834 800 75770 856
rect 75938 800 76874 856
rect 77042 800 77978 856
rect 78146 800 79082 856
rect 79250 800 79652 856
<< metal3 >>
rect 79200 152872 80000 152992
rect 79200 152056 80000 152176
rect 79200 151240 80000 151360
rect 79200 150424 80000 150544
rect 79200 149608 80000 149728
rect 79200 148792 80000 148912
rect 79200 147976 80000 148096
rect 79200 147160 80000 147280
rect 79200 146344 80000 146464
rect 79200 145528 80000 145648
rect 79200 144712 80000 144832
rect 79200 143896 80000 144016
rect 79200 143080 80000 143200
rect 79200 142264 80000 142384
rect 79200 141448 80000 141568
rect 79200 140632 80000 140752
rect 79200 139816 80000 139936
rect 79200 139000 80000 139120
rect 79200 138184 80000 138304
rect 79200 137368 80000 137488
rect 79200 136552 80000 136672
rect 79200 135736 80000 135856
rect 79200 134920 80000 135040
rect 79200 134104 80000 134224
rect 79200 133288 80000 133408
rect 79200 132472 80000 132592
rect 79200 131656 80000 131776
rect 79200 130840 80000 130960
rect 79200 130024 80000 130144
rect 79200 129208 80000 129328
rect 79200 128392 80000 128512
rect 79200 127576 80000 127696
rect 79200 126760 80000 126880
rect 79200 125944 80000 126064
rect 79200 125128 80000 125248
rect 79200 124312 80000 124432
rect 79200 123496 80000 123616
rect 79200 122680 80000 122800
rect 79200 121864 80000 121984
rect 79200 121048 80000 121168
rect 79200 120232 80000 120352
rect 79200 119416 80000 119536
rect 79200 118600 80000 118720
rect 79200 117784 80000 117904
rect 79200 116968 80000 117088
rect 79200 116152 80000 116272
rect 79200 115336 80000 115456
rect 79200 114520 80000 114640
rect 79200 113704 80000 113824
rect 79200 112888 80000 113008
rect 79200 112072 80000 112192
rect 79200 111256 80000 111376
rect 79200 110440 80000 110560
rect 79200 109624 80000 109744
rect 79200 108808 80000 108928
rect 79200 107992 80000 108112
rect 79200 107176 80000 107296
rect 79200 106360 80000 106480
rect 79200 105544 80000 105664
rect 79200 104728 80000 104848
rect 79200 103912 80000 104032
rect 79200 103096 80000 103216
rect 79200 102280 80000 102400
rect 79200 101464 80000 101584
rect 79200 100648 80000 100768
rect 79200 99832 80000 99952
rect 79200 99016 80000 99136
rect 79200 98200 80000 98320
rect 79200 97384 80000 97504
rect 79200 96568 80000 96688
rect 79200 95752 80000 95872
rect 79200 94936 80000 95056
rect 79200 94120 80000 94240
rect 79200 93304 80000 93424
rect 79200 92488 80000 92608
rect 79200 91672 80000 91792
rect 79200 90856 80000 90976
rect 79200 90040 80000 90160
rect 79200 89224 80000 89344
rect 79200 88408 80000 88528
rect 79200 87592 80000 87712
rect 79200 86776 80000 86896
rect 79200 85960 80000 86080
rect 79200 85144 80000 85264
rect 79200 84328 80000 84448
rect 79200 83512 80000 83632
rect 79200 82696 80000 82816
rect 79200 81880 80000 82000
rect 79200 81064 80000 81184
rect 79200 80248 80000 80368
rect 79200 79432 80000 79552
rect 79200 78616 80000 78736
rect 79200 77800 80000 77920
rect 79200 76984 80000 77104
rect 79200 76168 80000 76288
rect 79200 75352 80000 75472
rect 79200 74536 80000 74656
rect 79200 73720 80000 73840
rect 79200 72904 80000 73024
rect 79200 72088 80000 72208
rect 79200 71272 80000 71392
rect 79200 70456 80000 70576
rect 79200 69640 80000 69760
rect 79200 68824 80000 68944
rect 79200 68008 80000 68128
rect 79200 67192 80000 67312
rect 79200 66376 80000 66496
rect 79200 65560 80000 65680
rect 79200 64744 80000 64864
rect 79200 63928 80000 64048
rect 79200 63112 80000 63232
rect 79200 62296 80000 62416
rect 79200 61480 80000 61600
rect 79200 60664 80000 60784
rect 79200 59848 80000 59968
rect 79200 59032 80000 59152
rect 79200 58216 80000 58336
rect 79200 57400 80000 57520
rect 79200 56584 80000 56704
rect 79200 55768 80000 55888
rect 79200 54952 80000 55072
rect 79200 54136 80000 54256
rect 79200 53320 80000 53440
rect 79200 52504 80000 52624
rect 79200 51688 80000 51808
rect 79200 50872 80000 50992
rect 79200 50056 80000 50176
rect 79200 49240 80000 49360
rect 79200 48424 80000 48544
rect 79200 47608 80000 47728
rect 79200 46792 80000 46912
rect 79200 45976 80000 46096
rect 79200 45160 80000 45280
rect 79200 44344 80000 44464
rect 79200 43528 80000 43648
rect 79200 42712 80000 42832
rect 79200 41896 80000 42016
rect 79200 41080 80000 41200
rect 79200 40264 80000 40384
rect 79200 39448 80000 39568
rect 79200 38632 80000 38752
rect 79200 37816 80000 37936
rect 79200 37000 80000 37120
rect 79200 36184 80000 36304
rect 79200 35368 80000 35488
rect 79200 34552 80000 34672
rect 79200 33736 80000 33856
rect 79200 32920 80000 33040
rect 79200 32104 80000 32224
rect 79200 31288 80000 31408
rect 79200 30472 80000 30592
rect 79200 29656 80000 29776
rect 79200 28840 80000 28960
rect 79200 28024 80000 28144
rect 79200 27208 80000 27328
rect 79200 26392 80000 26512
rect 79200 25576 80000 25696
rect 79200 24760 80000 24880
rect 79200 23944 80000 24064
rect 79200 23128 80000 23248
rect 79200 22312 80000 22432
rect 79200 21496 80000 21616
rect 79200 20680 80000 20800
rect 79200 19864 80000 19984
rect 79200 19048 80000 19168
rect 79200 18232 80000 18352
rect 79200 17416 80000 17536
rect 79200 16600 80000 16720
rect 79200 15784 80000 15904
rect 79200 14968 80000 15088
rect 79200 14152 80000 14272
rect 79200 13336 80000 13456
rect 79200 12520 80000 12640
rect 79200 11704 80000 11824
rect 79200 10888 80000 11008
rect 79200 10072 80000 10192
rect 79200 9256 80000 9376
rect 79200 8440 80000 8560
rect 79200 7624 80000 7744
rect 79200 6808 80000 6928
<< obsm3 >>
rect 3601 153072 79200 157793
rect 3601 152792 79120 153072
rect 3601 152256 79200 152792
rect 3601 151976 79120 152256
rect 3601 151440 79200 151976
rect 3601 151160 79120 151440
rect 3601 150624 79200 151160
rect 3601 150344 79120 150624
rect 3601 149808 79200 150344
rect 3601 149528 79120 149808
rect 3601 148992 79200 149528
rect 3601 148712 79120 148992
rect 3601 148176 79200 148712
rect 3601 147896 79120 148176
rect 3601 147360 79200 147896
rect 3601 147080 79120 147360
rect 3601 146544 79200 147080
rect 3601 146264 79120 146544
rect 3601 145728 79200 146264
rect 3601 145448 79120 145728
rect 3601 144912 79200 145448
rect 3601 144632 79120 144912
rect 3601 144096 79200 144632
rect 3601 143816 79120 144096
rect 3601 143280 79200 143816
rect 3601 143000 79120 143280
rect 3601 142464 79200 143000
rect 3601 142184 79120 142464
rect 3601 141648 79200 142184
rect 3601 141368 79120 141648
rect 3601 140832 79200 141368
rect 3601 140552 79120 140832
rect 3601 140016 79200 140552
rect 3601 139736 79120 140016
rect 3601 139200 79200 139736
rect 3601 138920 79120 139200
rect 3601 138384 79200 138920
rect 3601 138104 79120 138384
rect 3601 137568 79200 138104
rect 3601 137288 79120 137568
rect 3601 136752 79200 137288
rect 3601 136472 79120 136752
rect 3601 135936 79200 136472
rect 3601 135656 79120 135936
rect 3601 135120 79200 135656
rect 3601 134840 79120 135120
rect 3601 134304 79200 134840
rect 3601 134024 79120 134304
rect 3601 133488 79200 134024
rect 3601 133208 79120 133488
rect 3601 132672 79200 133208
rect 3601 132392 79120 132672
rect 3601 131856 79200 132392
rect 3601 131576 79120 131856
rect 3601 131040 79200 131576
rect 3601 130760 79120 131040
rect 3601 130224 79200 130760
rect 3601 129944 79120 130224
rect 3601 129408 79200 129944
rect 3601 129128 79120 129408
rect 3601 128592 79200 129128
rect 3601 128312 79120 128592
rect 3601 127776 79200 128312
rect 3601 127496 79120 127776
rect 3601 126960 79200 127496
rect 3601 126680 79120 126960
rect 3601 126144 79200 126680
rect 3601 125864 79120 126144
rect 3601 125328 79200 125864
rect 3601 125048 79120 125328
rect 3601 124512 79200 125048
rect 3601 124232 79120 124512
rect 3601 123696 79200 124232
rect 3601 123416 79120 123696
rect 3601 122880 79200 123416
rect 3601 122600 79120 122880
rect 3601 122064 79200 122600
rect 3601 121784 79120 122064
rect 3601 121248 79200 121784
rect 3601 120968 79120 121248
rect 3601 120432 79200 120968
rect 3601 120152 79120 120432
rect 3601 119616 79200 120152
rect 3601 119336 79120 119616
rect 3601 118800 79200 119336
rect 3601 118520 79120 118800
rect 3601 117984 79200 118520
rect 3601 117704 79120 117984
rect 3601 117168 79200 117704
rect 3601 116888 79120 117168
rect 3601 116352 79200 116888
rect 3601 116072 79120 116352
rect 3601 115536 79200 116072
rect 3601 115256 79120 115536
rect 3601 114720 79200 115256
rect 3601 114440 79120 114720
rect 3601 113904 79200 114440
rect 3601 113624 79120 113904
rect 3601 113088 79200 113624
rect 3601 112808 79120 113088
rect 3601 112272 79200 112808
rect 3601 111992 79120 112272
rect 3601 111456 79200 111992
rect 3601 111176 79120 111456
rect 3601 110640 79200 111176
rect 3601 110360 79120 110640
rect 3601 109824 79200 110360
rect 3601 109544 79120 109824
rect 3601 109008 79200 109544
rect 3601 108728 79120 109008
rect 3601 108192 79200 108728
rect 3601 107912 79120 108192
rect 3601 107376 79200 107912
rect 3601 107096 79120 107376
rect 3601 106560 79200 107096
rect 3601 106280 79120 106560
rect 3601 105744 79200 106280
rect 3601 105464 79120 105744
rect 3601 104928 79200 105464
rect 3601 104648 79120 104928
rect 3601 104112 79200 104648
rect 3601 103832 79120 104112
rect 3601 103296 79200 103832
rect 3601 103016 79120 103296
rect 3601 102480 79200 103016
rect 3601 102200 79120 102480
rect 3601 101664 79200 102200
rect 3601 101384 79120 101664
rect 3601 100848 79200 101384
rect 3601 100568 79120 100848
rect 3601 100032 79200 100568
rect 3601 99752 79120 100032
rect 3601 99216 79200 99752
rect 3601 98936 79120 99216
rect 3601 98400 79200 98936
rect 3601 98120 79120 98400
rect 3601 97584 79200 98120
rect 3601 97304 79120 97584
rect 3601 96768 79200 97304
rect 3601 96488 79120 96768
rect 3601 95952 79200 96488
rect 3601 95672 79120 95952
rect 3601 95136 79200 95672
rect 3601 94856 79120 95136
rect 3601 94320 79200 94856
rect 3601 94040 79120 94320
rect 3601 93504 79200 94040
rect 3601 93224 79120 93504
rect 3601 92688 79200 93224
rect 3601 92408 79120 92688
rect 3601 91872 79200 92408
rect 3601 91592 79120 91872
rect 3601 91056 79200 91592
rect 3601 90776 79120 91056
rect 3601 90240 79200 90776
rect 3601 89960 79120 90240
rect 3601 89424 79200 89960
rect 3601 89144 79120 89424
rect 3601 88608 79200 89144
rect 3601 88328 79120 88608
rect 3601 87792 79200 88328
rect 3601 87512 79120 87792
rect 3601 86976 79200 87512
rect 3601 86696 79120 86976
rect 3601 86160 79200 86696
rect 3601 85880 79120 86160
rect 3601 85344 79200 85880
rect 3601 85064 79120 85344
rect 3601 84528 79200 85064
rect 3601 84248 79120 84528
rect 3601 83712 79200 84248
rect 3601 83432 79120 83712
rect 3601 82896 79200 83432
rect 3601 82616 79120 82896
rect 3601 82080 79200 82616
rect 3601 81800 79120 82080
rect 3601 81264 79200 81800
rect 3601 80984 79120 81264
rect 3601 80448 79200 80984
rect 3601 80168 79120 80448
rect 3601 79632 79200 80168
rect 3601 79352 79120 79632
rect 3601 78816 79200 79352
rect 3601 78536 79120 78816
rect 3601 78000 79200 78536
rect 3601 77720 79120 78000
rect 3601 77184 79200 77720
rect 3601 76904 79120 77184
rect 3601 76368 79200 76904
rect 3601 76088 79120 76368
rect 3601 75552 79200 76088
rect 3601 75272 79120 75552
rect 3601 74736 79200 75272
rect 3601 74456 79120 74736
rect 3601 73920 79200 74456
rect 3601 73640 79120 73920
rect 3601 73104 79200 73640
rect 3601 72824 79120 73104
rect 3601 72288 79200 72824
rect 3601 72008 79120 72288
rect 3601 71472 79200 72008
rect 3601 71192 79120 71472
rect 3601 70656 79200 71192
rect 3601 70376 79120 70656
rect 3601 69840 79200 70376
rect 3601 69560 79120 69840
rect 3601 69024 79200 69560
rect 3601 68744 79120 69024
rect 3601 68208 79200 68744
rect 3601 67928 79120 68208
rect 3601 67392 79200 67928
rect 3601 67112 79120 67392
rect 3601 66576 79200 67112
rect 3601 66296 79120 66576
rect 3601 65760 79200 66296
rect 3601 65480 79120 65760
rect 3601 64944 79200 65480
rect 3601 64664 79120 64944
rect 3601 64128 79200 64664
rect 3601 63848 79120 64128
rect 3601 63312 79200 63848
rect 3601 63032 79120 63312
rect 3601 62496 79200 63032
rect 3601 62216 79120 62496
rect 3601 61680 79200 62216
rect 3601 61400 79120 61680
rect 3601 60864 79200 61400
rect 3601 60584 79120 60864
rect 3601 60048 79200 60584
rect 3601 59768 79120 60048
rect 3601 59232 79200 59768
rect 3601 58952 79120 59232
rect 3601 58416 79200 58952
rect 3601 58136 79120 58416
rect 3601 57600 79200 58136
rect 3601 57320 79120 57600
rect 3601 56784 79200 57320
rect 3601 56504 79120 56784
rect 3601 55968 79200 56504
rect 3601 55688 79120 55968
rect 3601 55152 79200 55688
rect 3601 54872 79120 55152
rect 3601 54336 79200 54872
rect 3601 54056 79120 54336
rect 3601 53520 79200 54056
rect 3601 53240 79120 53520
rect 3601 52704 79200 53240
rect 3601 52424 79120 52704
rect 3601 51888 79200 52424
rect 3601 51608 79120 51888
rect 3601 51072 79200 51608
rect 3601 50792 79120 51072
rect 3601 50256 79200 50792
rect 3601 49976 79120 50256
rect 3601 49440 79200 49976
rect 3601 49160 79120 49440
rect 3601 48624 79200 49160
rect 3601 48344 79120 48624
rect 3601 47808 79200 48344
rect 3601 47528 79120 47808
rect 3601 46992 79200 47528
rect 3601 46712 79120 46992
rect 3601 46176 79200 46712
rect 3601 45896 79120 46176
rect 3601 45360 79200 45896
rect 3601 45080 79120 45360
rect 3601 44544 79200 45080
rect 3601 44264 79120 44544
rect 3601 43728 79200 44264
rect 3601 43448 79120 43728
rect 3601 42912 79200 43448
rect 3601 42632 79120 42912
rect 3601 42096 79200 42632
rect 3601 41816 79120 42096
rect 3601 41280 79200 41816
rect 3601 41000 79120 41280
rect 3601 40464 79200 41000
rect 3601 40184 79120 40464
rect 3601 39648 79200 40184
rect 3601 39368 79120 39648
rect 3601 38832 79200 39368
rect 3601 38552 79120 38832
rect 3601 38016 79200 38552
rect 3601 37736 79120 38016
rect 3601 37200 79200 37736
rect 3601 36920 79120 37200
rect 3601 36384 79200 36920
rect 3601 36104 79120 36384
rect 3601 35568 79200 36104
rect 3601 35288 79120 35568
rect 3601 34752 79200 35288
rect 3601 34472 79120 34752
rect 3601 33936 79200 34472
rect 3601 33656 79120 33936
rect 3601 33120 79200 33656
rect 3601 32840 79120 33120
rect 3601 32304 79200 32840
rect 3601 32024 79120 32304
rect 3601 31488 79200 32024
rect 3601 31208 79120 31488
rect 3601 30672 79200 31208
rect 3601 30392 79120 30672
rect 3601 29856 79200 30392
rect 3601 29576 79120 29856
rect 3601 29040 79200 29576
rect 3601 28760 79120 29040
rect 3601 28224 79200 28760
rect 3601 27944 79120 28224
rect 3601 27408 79200 27944
rect 3601 27128 79120 27408
rect 3601 26592 79200 27128
rect 3601 26312 79120 26592
rect 3601 25776 79200 26312
rect 3601 25496 79120 25776
rect 3601 24960 79200 25496
rect 3601 24680 79120 24960
rect 3601 24144 79200 24680
rect 3601 23864 79120 24144
rect 3601 23328 79200 23864
rect 3601 23048 79120 23328
rect 3601 22512 79200 23048
rect 3601 22232 79120 22512
rect 3601 21696 79200 22232
rect 3601 21416 79120 21696
rect 3601 20880 79200 21416
rect 3601 20600 79120 20880
rect 3601 20064 79200 20600
rect 3601 19784 79120 20064
rect 3601 19248 79200 19784
rect 3601 18968 79120 19248
rect 3601 18432 79200 18968
rect 3601 18152 79120 18432
rect 3601 17616 79200 18152
rect 3601 17336 79120 17616
rect 3601 16800 79200 17336
rect 3601 16520 79120 16800
rect 3601 15984 79200 16520
rect 3601 15704 79120 15984
rect 3601 15168 79200 15704
rect 3601 14888 79120 15168
rect 3601 14352 79200 14888
rect 3601 14072 79120 14352
rect 3601 13536 79200 14072
rect 3601 13256 79120 13536
rect 3601 12720 79200 13256
rect 3601 12440 79120 12720
rect 3601 11904 79200 12440
rect 3601 11624 79120 11904
rect 3601 11088 79200 11624
rect 3601 10808 79120 11088
rect 3601 10272 79200 10808
rect 3601 9992 79120 10272
rect 3601 9456 79200 9992
rect 3601 9176 79120 9456
rect 3601 8640 79200 9176
rect 3601 8360 79120 8640
rect 3601 7824 79200 8360
rect 3601 7544 79120 7824
rect 3601 7008 79200 7544
rect 3601 6728 79120 7008
rect 3601 2143 79200 6728
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
<< obsm4 >>
rect 36307 3707 50208 154597
rect 50688 3707 65568 154597
rect 66048 3707 77221 154597
<< labels >>
rlabel metal2 s 754 0 810 800 6 dbg_in[0]
port 1 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 dbg_in[1]
port 2 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 dbg_in[2]
port 3 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 dbg_in[3]
port 4 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 dbg_out[0]
port 5 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 dbg_out[10]
port 6 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 dbg_out[11]
port 7 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 dbg_out[12]
port 8 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 dbg_out[13]
port 9 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 dbg_out[14]
port 10 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 dbg_out[15]
port 11 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 dbg_out[16]
port 12 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 dbg_out[17]
port 13 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 dbg_out[18]
port 14 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 dbg_out[19]
port 15 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 dbg_out[1]
port 16 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 dbg_out[20]
port 17 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 dbg_out[21]
port 18 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 dbg_out[22]
port 19 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 dbg_out[23]
port 20 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 dbg_out[24]
port 21 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 dbg_out[25]
port 22 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 dbg_out[26]
port 23 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 dbg_out[27]
port 24 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 dbg_out[28]
port 25 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 dbg_out[29]
port 26 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 dbg_out[2]
port 27 nsew signal output
rlabel metal2 s 73618 0 73674 800 6 dbg_out[30]
port 28 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 dbg_out[31]
port 29 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 dbg_out[32]
port 30 nsew signal output
rlabel metal2 s 76930 0 76986 800 6 dbg_out[33]
port 31 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 dbg_out[34]
port 32 nsew signal output
rlabel metal2 s 79138 0 79194 800 6 dbg_out[35]
port 33 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 dbg_out[3]
port 34 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 dbg_out[4]
port 35 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 dbg_out[5]
port 36 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 dbg_out[6]
port 37 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 dbg_out[7]
port 38 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 dbg_out[8]
port 39 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 dbg_out[9]
port 40 nsew signal output
rlabel metal2 s 2962 0 3018 800 6 dbg_pc[0]
port 41 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 dbg_pc[10]
port 42 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 dbg_pc[11]
port 43 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 dbg_pc[12]
port 44 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 dbg_pc[13]
port 45 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 dbg_pc[14]
port 46 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 dbg_pc[15]
port 47 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 dbg_pc[1]
port 48 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 dbg_pc[2]
port 49 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 dbg_pc[3]
port 50 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 dbg_pc[4]
port 51 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 dbg_pc[5]
port 52 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 dbg_pc[6]
port 53 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 dbg_pc[7]
port 54 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 dbg_pc[8]
port 55 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 dbg_pc[9]
port 56 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 dbg_r0[0]
port 57 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 dbg_r0[10]
port 58 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 dbg_r0[11]
port 59 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 dbg_r0[12]
port 60 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 dbg_r0[13]
port 61 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 dbg_r0[14]
port 62 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 dbg_r0[15]
port 63 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 dbg_r0[1]
port 64 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 dbg_r0[2]
port 65 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 dbg_r0[3]
port 66 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 dbg_r0[4]
port 67 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 dbg_r0[5]
port 68 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 dbg_r0[6]
port 69 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 dbg_r0[7]
port 70 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 dbg_r0[8]
port 71 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 dbg_r0[9]
port 72 nsew signal output
rlabel metal3 s 79200 6808 80000 6928 6 i_clk
port 73 nsew signal input
rlabel metal3 s 79200 140632 80000 140752 6 i_core_int_sreg[0]
port 74 nsew signal input
rlabel metal3 s 79200 148792 80000 148912 6 i_core_int_sreg[10]
port 75 nsew signal input
rlabel metal3 s 79200 149608 80000 149728 6 i_core_int_sreg[11]
port 76 nsew signal input
rlabel metal3 s 79200 150424 80000 150544 6 i_core_int_sreg[12]
port 77 nsew signal input
rlabel metal3 s 79200 151240 80000 151360 6 i_core_int_sreg[13]
port 78 nsew signal input
rlabel metal3 s 79200 152056 80000 152176 6 i_core_int_sreg[14]
port 79 nsew signal input
rlabel metal3 s 79200 152872 80000 152992 6 i_core_int_sreg[15]
port 80 nsew signal input
rlabel metal3 s 79200 141448 80000 141568 6 i_core_int_sreg[1]
port 81 nsew signal input
rlabel metal3 s 79200 142264 80000 142384 6 i_core_int_sreg[2]
port 82 nsew signal input
rlabel metal3 s 79200 143080 80000 143200 6 i_core_int_sreg[3]
port 83 nsew signal input
rlabel metal3 s 79200 143896 80000 144016 6 i_core_int_sreg[4]
port 84 nsew signal input
rlabel metal3 s 79200 144712 80000 144832 6 i_core_int_sreg[5]
port 85 nsew signal input
rlabel metal3 s 79200 145528 80000 145648 6 i_core_int_sreg[6]
port 86 nsew signal input
rlabel metal3 s 79200 146344 80000 146464 6 i_core_int_sreg[7]
port 87 nsew signal input
rlabel metal3 s 79200 147160 80000 147280 6 i_core_int_sreg[8]
port 88 nsew signal input
rlabel metal3 s 79200 147976 80000 148096 6 i_core_int_sreg[9]
port 89 nsew signal input
rlabel metal3 s 79200 139000 80000 139120 6 i_disable
port 90 nsew signal input
rlabel metal3 s 79200 108808 80000 108928 6 i_irq
port 91 nsew signal input
rlabel metal3 s 79200 139816 80000 139936 6 i_mc_core_int
port 92 nsew signal input
rlabel metal3 s 79200 57400 80000 57520 6 i_mem_ack
port 93 nsew signal input
rlabel metal3 s 79200 28024 80000 28144 6 i_mem_data[0]
port 94 nsew signal input
rlabel metal3 s 79200 44344 80000 44464 6 i_mem_data[10]
port 95 nsew signal input
rlabel metal3 s 79200 45976 80000 46096 6 i_mem_data[11]
port 96 nsew signal input
rlabel metal3 s 79200 47608 80000 47728 6 i_mem_data[12]
port 97 nsew signal input
rlabel metal3 s 79200 49240 80000 49360 6 i_mem_data[13]
port 98 nsew signal input
rlabel metal3 s 79200 50872 80000 50992 6 i_mem_data[14]
port 99 nsew signal input
rlabel metal3 s 79200 52504 80000 52624 6 i_mem_data[15]
port 100 nsew signal input
rlabel metal3 s 79200 29656 80000 29776 6 i_mem_data[1]
port 101 nsew signal input
rlabel metal3 s 79200 31288 80000 31408 6 i_mem_data[2]
port 102 nsew signal input
rlabel metal3 s 79200 32920 80000 33040 6 i_mem_data[3]
port 103 nsew signal input
rlabel metal3 s 79200 34552 80000 34672 6 i_mem_data[4]
port 104 nsew signal input
rlabel metal3 s 79200 36184 80000 36304 6 i_mem_data[5]
port 105 nsew signal input
rlabel metal3 s 79200 37816 80000 37936 6 i_mem_data[6]
port 106 nsew signal input
rlabel metal3 s 79200 39448 80000 39568 6 i_mem_data[7]
port 107 nsew signal input
rlabel metal3 s 79200 41080 80000 41200 6 i_mem_data[8]
port 108 nsew signal input
rlabel metal3 s 79200 42712 80000 42832 6 i_mem_data[9]
port 109 nsew signal input
rlabel metal3 s 79200 58216 80000 58336 6 i_mem_exception
port 110 nsew signal input
rlabel metal3 s 79200 61480 80000 61600 6 i_req_data[0]
port 111 nsew signal input
rlabel metal3 s 79200 77800 80000 77920 6 i_req_data[10]
port 112 nsew signal input
rlabel metal3 s 79200 79432 80000 79552 6 i_req_data[11]
port 113 nsew signal input
rlabel metal3 s 79200 81064 80000 81184 6 i_req_data[12]
port 114 nsew signal input
rlabel metal3 s 79200 82696 80000 82816 6 i_req_data[13]
port 115 nsew signal input
rlabel metal3 s 79200 84328 80000 84448 6 i_req_data[14]
port 116 nsew signal input
rlabel metal3 s 79200 85960 80000 86080 6 i_req_data[15]
port 117 nsew signal input
rlabel metal3 s 79200 87592 80000 87712 6 i_req_data[16]
port 118 nsew signal input
rlabel metal3 s 79200 88408 80000 88528 6 i_req_data[17]
port 119 nsew signal input
rlabel metal3 s 79200 89224 80000 89344 6 i_req_data[18]
port 120 nsew signal input
rlabel metal3 s 79200 90040 80000 90160 6 i_req_data[19]
port 121 nsew signal input
rlabel metal3 s 79200 63112 80000 63232 6 i_req_data[1]
port 122 nsew signal input
rlabel metal3 s 79200 90856 80000 90976 6 i_req_data[20]
port 123 nsew signal input
rlabel metal3 s 79200 91672 80000 91792 6 i_req_data[21]
port 124 nsew signal input
rlabel metal3 s 79200 92488 80000 92608 6 i_req_data[22]
port 125 nsew signal input
rlabel metal3 s 79200 93304 80000 93424 6 i_req_data[23]
port 126 nsew signal input
rlabel metal3 s 79200 94120 80000 94240 6 i_req_data[24]
port 127 nsew signal input
rlabel metal3 s 79200 94936 80000 95056 6 i_req_data[25]
port 128 nsew signal input
rlabel metal3 s 79200 95752 80000 95872 6 i_req_data[26]
port 129 nsew signal input
rlabel metal3 s 79200 96568 80000 96688 6 i_req_data[27]
port 130 nsew signal input
rlabel metal3 s 79200 97384 80000 97504 6 i_req_data[28]
port 131 nsew signal input
rlabel metal3 s 79200 98200 80000 98320 6 i_req_data[29]
port 132 nsew signal input
rlabel metal3 s 79200 64744 80000 64864 6 i_req_data[2]
port 133 nsew signal input
rlabel metal3 s 79200 99016 80000 99136 6 i_req_data[30]
port 134 nsew signal input
rlabel metal3 s 79200 99832 80000 99952 6 i_req_data[31]
port 135 nsew signal input
rlabel metal3 s 79200 66376 80000 66496 6 i_req_data[3]
port 136 nsew signal input
rlabel metal3 s 79200 68008 80000 68128 6 i_req_data[4]
port 137 nsew signal input
rlabel metal3 s 79200 69640 80000 69760 6 i_req_data[5]
port 138 nsew signal input
rlabel metal3 s 79200 71272 80000 71392 6 i_req_data[6]
port 139 nsew signal input
rlabel metal3 s 79200 72904 80000 73024 6 i_req_data[7]
port 140 nsew signal input
rlabel metal3 s 79200 74536 80000 74656 6 i_req_data[8]
port 141 nsew signal input
rlabel metal3 s 79200 76168 80000 76288 6 i_req_data[9]
port 142 nsew signal input
rlabel metal3 s 79200 59032 80000 59152 6 i_req_data_valid
port 143 nsew signal input
rlabel metal3 s 79200 7624 80000 7744 6 i_rst
port 144 nsew signal input
rlabel metal3 s 79200 109624 80000 109744 6 o_c_data_page
port 145 nsew signal output
rlabel metal3 s 79200 100648 80000 100768 6 o_c_instr_long
port 146 nsew signal output
rlabel metal3 s 79200 110440 80000 110560 6 o_c_instr_page
port 147 nsew signal output
rlabel metal3 s 79200 138184 80000 138304 6 o_icache_flush
port 148 nsew signal output
rlabel metal3 s 79200 102280 80000 102400 6 o_instr_long_addr[0]
port 149 nsew signal output
rlabel metal3 s 79200 103096 80000 103216 6 o_instr_long_addr[1]
port 150 nsew signal output
rlabel metal3 s 79200 103912 80000 104032 6 o_instr_long_addr[2]
port 151 nsew signal output
rlabel metal3 s 79200 104728 80000 104848 6 o_instr_long_addr[3]
port 152 nsew signal output
rlabel metal3 s 79200 105544 80000 105664 6 o_instr_long_addr[4]
port 153 nsew signal output
rlabel metal3 s 79200 106360 80000 106480 6 o_instr_long_addr[5]
port 154 nsew signal output
rlabel metal3 s 79200 107176 80000 107296 6 o_instr_long_addr[6]
port 155 nsew signal output
rlabel metal3 s 79200 107992 80000 108112 6 o_instr_long_addr[7]
port 156 nsew signal output
rlabel metal3 s 79200 8440 80000 8560 6 o_mem_addr[0]
port 157 nsew signal output
rlabel metal3 s 79200 23128 80000 23248 6 o_mem_addr[10]
port 158 nsew signal output
rlabel metal3 s 79200 23944 80000 24064 6 o_mem_addr[11]
port 159 nsew signal output
rlabel metal3 s 79200 24760 80000 24880 6 o_mem_addr[12]
port 160 nsew signal output
rlabel metal3 s 79200 25576 80000 25696 6 o_mem_addr[13]
port 161 nsew signal output
rlabel metal3 s 79200 26392 80000 26512 6 o_mem_addr[14]
port 162 nsew signal output
rlabel metal3 s 79200 27208 80000 27328 6 o_mem_addr[15]
port 163 nsew signal output
rlabel metal3 s 79200 10072 80000 10192 6 o_mem_addr[1]
port 164 nsew signal output
rlabel metal3 s 79200 11704 80000 11824 6 o_mem_addr[2]
port 165 nsew signal output
rlabel metal3 s 79200 13336 80000 13456 6 o_mem_addr[3]
port 166 nsew signal output
rlabel metal3 s 79200 14968 80000 15088 6 o_mem_addr[4]
port 167 nsew signal output
rlabel metal3 s 79200 16600 80000 16720 6 o_mem_addr[5]
port 168 nsew signal output
rlabel metal3 s 79200 18232 80000 18352 6 o_mem_addr[6]
port 169 nsew signal output
rlabel metal3 s 79200 19864 80000 19984 6 o_mem_addr[7]
port 170 nsew signal output
rlabel metal3 s 79200 21496 80000 21616 6 o_mem_addr[8]
port 171 nsew signal output
rlabel metal3 s 79200 22312 80000 22432 6 o_mem_addr[9]
port 172 nsew signal output
rlabel metal3 s 79200 9256 80000 9376 6 o_mem_addr_high[0]
port 173 nsew signal output
rlabel metal3 s 79200 10888 80000 11008 6 o_mem_addr_high[1]
port 174 nsew signal output
rlabel metal3 s 79200 12520 80000 12640 6 o_mem_addr_high[2]
port 175 nsew signal output
rlabel metal3 s 79200 14152 80000 14272 6 o_mem_addr_high[3]
port 176 nsew signal output
rlabel metal3 s 79200 15784 80000 15904 6 o_mem_addr_high[4]
port 177 nsew signal output
rlabel metal3 s 79200 17416 80000 17536 6 o_mem_addr_high[5]
port 178 nsew signal output
rlabel metal3 s 79200 19048 80000 19168 6 o_mem_addr_high[6]
port 179 nsew signal output
rlabel metal3 s 79200 20680 80000 20800 6 o_mem_addr_high[7]
port 180 nsew signal output
rlabel metal3 s 79200 28840 80000 28960 6 o_mem_data[0]
port 181 nsew signal output
rlabel metal3 s 79200 45160 80000 45280 6 o_mem_data[10]
port 182 nsew signal output
rlabel metal3 s 79200 46792 80000 46912 6 o_mem_data[11]
port 183 nsew signal output
rlabel metal3 s 79200 48424 80000 48544 6 o_mem_data[12]
port 184 nsew signal output
rlabel metal3 s 79200 50056 80000 50176 6 o_mem_data[13]
port 185 nsew signal output
rlabel metal3 s 79200 51688 80000 51808 6 o_mem_data[14]
port 186 nsew signal output
rlabel metal3 s 79200 53320 80000 53440 6 o_mem_data[15]
port 187 nsew signal output
rlabel metal3 s 79200 30472 80000 30592 6 o_mem_data[1]
port 188 nsew signal output
rlabel metal3 s 79200 32104 80000 32224 6 o_mem_data[2]
port 189 nsew signal output
rlabel metal3 s 79200 33736 80000 33856 6 o_mem_data[3]
port 190 nsew signal output
rlabel metal3 s 79200 35368 80000 35488 6 o_mem_data[4]
port 191 nsew signal output
rlabel metal3 s 79200 37000 80000 37120 6 o_mem_data[5]
port 192 nsew signal output
rlabel metal3 s 79200 38632 80000 38752 6 o_mem_data[6]
port 193 nsew signal output
rlabel metal3 s 79200 40264 80000 40384 6 o_mem_data[7]
port 194 nsew signal output
rlabel metal3 s 79200 41896 80000 42016 6 o_mem_data[8]
port 195 nsew signal output
rlabel metal3 s 79200 43528 80000 43648 6 o_mem_data[9]
port 196 nsew signal output
rlabel metal3 s 79200 101464 80000 101584 6 o_mem_long
port 197 nsew signal output
rlabel metal3 s 79200 54136 80000 54256 6 o_mem_req
port 198 nsew signal output
rlabel metal3 s 79200 55768 80000 55888 6 o_mem_sel[0]
port 199 nsew signal output
rlabel metal3 s 79200 56584 80000 56704 6 o_mem_sel[1]
port 200 nsew signal output
rlabel metal3 s 79200 54952 80000 55072 6 o_mem_we
port 201 nsew signal output
rlabel metal3 s 79200 59848 80000 59968 6 o_req_active
port 202 nsew signal output
rlabel metal3 s 79200 62296 80000 62416 6 o_req_addr[0]
port 203 nsew signal output
rlabel metal3 s 79200 78616 80000 78736 6 o_req_addr[10]
port 204 nsew signal output
rlabel metal3 s 79200 80248 80000 80368 6 o_req_addr[11]
port 205 nsew signal output
rlabel metal3 s 79200 81880 80000 82000 6 o_req_addr[12]
port 206 nsew signal output
rlabel metal3 s 79200 83512 80000 83632 6 o_req_addr[13]
port 207 nsew signal output
rlabel metal3 s 79200 85144 80000 85264 6 o_req_addr[14]
port 208 nsew signal output
rlabel metal3 s 79200 86776 80000 86896 6 o_req_addr[15]
port 209 nsew signal output
rlabel metal3 s 79200 63928 80000 64048 6 o_req_addr[1]
port 210 nsew signal output
rlabel metal3 s 79200 65560 80000 65680 6 o_req_addr[2]
port 211 nsew signal output
rlabel metal3 s 79200 67192 80000 67312 6 o_req_addr[3]
port 212 nsew signal output
rlabel metal3 s 79200 68824 80000 68944 6 o_req_addr[4]
port 213 nsew signal output
rlabel metal3 s 79200 70456 80000 70576 6 o_req_addr[5]
port 214 nsew signal output
rlabel metal3 s 79200 72088 80000 72208 6 o_req_addr[6]
port 215 nsew signal output
rlabel metal3 s 79200 73720 80000 73840 6 o_req_addr[7]
port 216 nsew signal output
rlabel metal3 s 79200 75352 80000 75472 6 o_req_addr[8]
port 217 nsew signal output
rlabel metal3 s 79200 76984 80000 77104 6 o_req_addr[9]
port 218 nsew signal output
rlabel metal3 s 79200 60664 80000 60784 6 o_req_ppl_submit
port 219 nsew signal output
rlabel metal3 s 79200 112072 80000 112192 6 sr_bus_addr[0]
port 220 nsew signal output
rlabel metal3 s 79200 128392 80000 128512 6 sr_bus_addr[10]
port 221 nsew signal output
rlabel metal3 s 79200 130024 80000 130144 6 sr_bus_addr[11]
port 222 nsew signal output
rlabel metal3 s 79200 131656 80000 131776 6 sr_bus_addr[12]
port 223 nsew signal output
rlabel metal3 s 79200 133288 80000 133408 6 sr_bus_addr[13]
port 224 nsew signal output
rlabel metal3 s 79200 134920 80000 135040 6 sr_bus_addr[14]
port 225 nsew signal output
rlabel metal3 s 79200 136552 80000 136672 6 sr_bus_addr[15]
port 226 nsew signal output
rlabel metal3 s 79200 113704 80000 113824 6 sr_bus_addr[1]
port 227 nsew signal output
rlabel metal3 s 79200 115336 80000 115456 6 sr_bus_addr[2]
port 228 nsew signal output
rlabel metal3 s 79200 116968 80000 117088 6 sr_bus_addr[3]
port 229 nsew signal output
rlabel metal3 s 79200 118600 80000 118720 6 sr_bus_addr[4]
port 230 nsew signal output
rlabel metal3 s 79200 120232 80000 120352 6 sr_bus_addr[5]
port 231 nsew signal output
rlabel metal3 s 79200 121864 80000 121984 6 sr_bus_addr[6]
port 232 nsew signal output
rlabel metal3 s 79200 123496 80000 123616 6 sr_bus_addr[7]
port 233 nsew signal output
rlabel metal3 s 79200 125128 80000 125248 6 sr_bus_addr[8]
port 234 nsew signal output
rlabel metal3 s 79200 126760 80000 126880 6 sr_bus_addr[9]
port 235 nsew signal output
rlabel metal3 s 79200 112888 80000 113008 6 sr_bus_data_o[0]
port 236 nsew signal output
rlabel metal3 s 79200 129208 80000 129328 6 sr_bus_data_o[10]
port 237 nsew signal output
rlabel metal3 s 79200 130840 80000 130960 6 sr_bus_data_o[11]
port 238 nsew signal output
rlabel metal3 s 79200 132472 80000 132592 6 sr_bus_data_o[12]
port 239 nsew signal output
rlabel metal3 s 79200 134104 80000 134224 6 sr_bus_data_o[13]
port 240 nsew signal output
rlabel metal3 s 79200 135736 80000 135856 6 sr_bus_data_o[14]
port 241 nsew signal output
rlabel metal3 s 79200 137368 80000 137488 6 sr_bus_data_o[15]
port 242 nsew signal output
rlabel metal3 s 79200 114520 80000 114640 6 sr_bus_data_o[1]
port 243 nsew signal output
rlabel metal3 s 79200 116152 80000 116272 6 sr_bus_data_o[2]
port 244 nsew signal output
rlabel metal3 s 79200 117784 80000 117904 6 sr_bus_data_o[3]
port 245 nsew signal output
rlabel metal3 s 79200 119416 80000 119536 6 sr_bus_data_o[4]
port 246 nsew signal output
rlabel metal3 s 79200 121048 80000 121168 6 sr_bus_data_o[5]
port 247 nsew signal output
rlabel metal3 s 79200 122680 80000 122800 6 sr_bus_data_o[6]
port 248 nsew signal output
rlabel metal3 s 79200 124312 80000 124432 6 sr_bus_data_o[7]
port 249 nsew signal output
rlabel metal3 s 79200 125944 80000 126064 6 sr_bus_data_o[8]
port 250 nsew signal output
rlabel metal3 s 79200 127576 80000 127696 6 sr_bus_data_o[9]
port 251 nsew signal output
rlabel metal3 s 79200 111256 80000 111376 6 sr_bus_we
port 252 nsew signal output
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 253 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 253 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 253 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 254 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 254 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 19491458
string GDS_FILE /home/piotro/caravel_user_project/openlane/core0/runs/22_12_28_20_46/results/signoff/core.magic.gds
string GDS_START 1248270
<< end >>

