magic
tech gf180mcuD
magscale 1 10
timestamp 1700095739
<< nwell >>
rect 1258 175968 534662 176486
rect 1258 175239 67389 175264
rect 1258 174425 534662 175239
rect 1258 174400 61341 174425
rect 1258 173671 60893 173696
rect 1258 172857 534662 173671
rect 1258 172832 109725 172857
rect 1258 172103 75565 172128
rect 1258 171289 534662 172103
rect 1258 171264 57533 171289
rect 1258 170535 57645 170560
rect 1258 169721 534662 170535
rect 1258 169696 65709 169721
rect 1258 168967 75005 168992
rect 1258 168153 534662 168967
rect 1258 168128 87661 168153
rect 1258 167399 57421 167424
rect 1258 166585 534662 167399
rect 1258 166560 56861 166585
rect 1258 165831 78296 165856
rect 1258 165017 534662 165831
rect 1258 164992 57421 165017
rect 1258 164263 65261 164288
rect 1258 163449 534662 164263
rect 1258 163424 57085 163449
rect 1258 162695 96845 162720
rect 1258 161881 534662 162695
rect 1258 161856 94045 161881
rect 1258 161127 65933 161152
rect 1258 160313 534662 161127
rect 1258 160288 41629 160313
rect 1258 159559 29757 159584
rect 1258 158745 534662 159559
rect 1258 158720 29981 158745
rect 1258 157991 36141 158016
rect 1258 157177 534662 157991
rect 1258 157152 47453 157177
rect 1258 156423 29240 156448
rect 1258 155609 534662 156423
rect 1258 155584 48461 155609
rect 1258 154855 30429 154880
rect 1258 154041 534662 154855
rect 1258 154016 65709 154041
rect 1258 153287 36141 153312
rect 1258 152473 534662 153287
rect 1258 152448 57869 152473
rect 1258 151719 26509 151744
rect 1258 150905 534662 151719
rect 1258 150880 26397 150905
rect 1258 150151 26621 150176
rect 1258 149337 534662 150151
rect 1258 149312 31997 149337
rect 1258 148583 20573 148608
rect 1258 147769 534662 148583
rect 1258 147744 39501 147769
rect 1258 147015 20685 147040
rect 1258 146201 534662 147015
rect 1258 146176 46781 146201
rect 1258 145447 20013 145472
rect 1258 144633 534662 145447
rect 1258 144608 24829 144633
rect 1258 143879 20685 143904
rect 1258 143065 534662 143879
rect 1258 143040 41784 143065
rect 1258 142311 30429 142336
rect 1258 141497 534662 142311
rect 1258 141472 16317 141497
rect 1258 140743 14749 140768
rect 1258 139929 534662 140743
rect 1258 139904 8477 139929
rect 1258 139175 26061 139200
rect 1258 138361 534662 139175
rect 1258 138336 16653 138361
rect 1258 137607 6909 137632
rect 1258 136793 534662 137607
rect 1258 136768 25949 136793
rect 1258 136039 13741 136064
rect 1258 135225 534662 136039
rect 1258 135200 7848 135225
rect 1258 134471 28301 134496
rect 1258 133657 534662 134471
rect 1258 133632 8589 133657
rect 1258 132903 20237 132928
rect 1258 132089 534662 132903
rect 1258 132064 39837 132089
rect 1258 131335 50365 131360
rect 1258 130521 534662 131335
rect 1258 130496 15981 130521
rect 1258 129767 10381 129792
rect 1258 128953 534662 129767
rect 1258 128928 10157 128953
rect 1258 128199 19901 128224
rect 1258 127385 534662 128199
rect 1258 127360 15981 127385
rect 1258 126631 33901 126656
rect 1258 125817 534662 126631
rect 1258 125792 10045 125817
rect 1258 125063 10381 125088
rect 1258 124249 534662 125063
rect 1258 124224 15197 124249
rect 1258 123495 27965 123520
rect 1258 122681 534662 123495
rect 1258 122656 23597 122681
rect 1258 121927 27517 121952
rect 1258 121113 534662 121927
rect 1258 121088 10829 121113
rect 1258 120359 19453 120384
rect 1258 119545 534662 120359
rect 1258 119520 9037 119545
rect 1258 118791 11949 118816
rect 1258 117977 534662 118791
rect 1258 117952 26440 117977
rect 1258 117223 38269 117248
rect 1258 116409 534662 117223
rect 1258 116384 31997 116409
rect 1258 115655 85309 115680
rect 1258 114841 534662 115655
rect 1258 114816 8477 114841
rect 1258 114087 14301 114112
rect 1258 113273 534662 114087
rect 1258 113248 9304 113273
rect 1258 112519 27965 112544
rect 1258 111705 534662 112519
rect 1258 111680 22141 111705
rect 1258 110951 10829 110976
rect 1258 110137 534662 110951
rect 1258 110112 7624 110137
rect 1258 109383 13629 109408
rect 1258 108569 534662 109383
rect 1258 108544 30093 108569
rect 1258 107815 10717 107840
rect 1258 107001 534662 107815
rect 1258 106976 22141 107001
rect 1258 106247 10717 106272
rect 1258 105433 534662 106247
rect 1258 105408 63581 105433
rect 1258 104679 18445 104704
rect 1258 103865 534662 104679
rect 1258 103840 10829 103865
rect 1258 103111 10381 103136
rect 1258 102297 534662 103111
rect 1258 102272 17101 102297
rect 1258 101543 20125 101568
rect 1258 100729 534662 101543
rect 1258 100704 18669 100729
rect 1258 99975 27741 100000
rect 1258 99161 534662 99975
rect 1258 99136 26509 99161
rect 1258 98407 77469 98432
rect 1258 97593 534662 98407
rect 1258 97568 18669 97593
rect 1258 96839 19565 96864
rect 1258 96025 534662 96839
rect 1258 96000 16317 96025
rect 1258 95271 12173 95296
rect 1258 94457 534662 95271
rect 1258 94432 73549 94457
rect 1258 93703 12397 93728
rect 1258 92889 534662 93703
rect 1258 92864 19720 92889
rect 1258 92135 26397 92160
rect 1258 91321 534662 92135
rect 1258 91296 23037 91321
rect 1258 90567 13517 90592
rect 1258 89753 534662 90567
rect 1258 89728 8813 89753
rect 1258 88999 10381 89024
rect 1258 88185 534662 88999
rect 1258 88160 8813 88185
rect 1258 87431 20461 87456
rect 1258 86617 534662 87431
rect 1258 86592 32109 86617
rect 1258 85863 67277 85888
rect 1258 85049 534662 85863
rect 1258 85024 6461 85049
rect 1258 84295 5229 84320
rect 1258 83481 534662 84295
rect 1258 83456 22925 83481
rect 1258 82727 6909 82752
rect 1258 81913 534662 82727
rect 1258 81888 6461 81913
rect 1258 81159 14301 81184
rect 1258 80345 534662 81159
rect 1258 80320 48573 80345
rect 1258 79591 4557 79616
rect 1258 78777 534662 79591
rect 1258 78752 7736 78777
rect 1258 78023 5453 78048
rect 1258 77209 534662 78023
rect 1258 77184 15197 77209
rect 1258 76455 20573 76480
rect 1258 75641 534662 76455
rect 1258 75616 7805 75641
rect 1258 74887 5453 74912
rect 1258 74073 534662 74887
rect 1258 74048 25768 74073
rect 1258 73319 4445 73344
rect 1258 72505 534662 73319
rect 1258 72480 14525 72505
rect 1258 71751 4333 71776
rect 1258 70937 534662 71751
rect 1258 70912 24381 70937
rect 1258 70183 4781 70208
rect 1258 69369 534662 70183
rect 1258 69344 45661 69369
rect 1258 68615 5005 68640
rect 1258 67801 534662 68615
rect 1258 67776 23261 67801
rect 1258 67047 5341 67072
rect 1258 66233 534662 67047
rect 1258 66208 45997 66233
rect 1258 65479 30024 65504
rect 1258 64665 534662 65479
rect 1258 64640 25053 64665
rect 1258 63911 5565 63936
rect 1258 63097 534662 63911
rect 1258 63072 147581 63097
rect 1258 62343 5005 62368
rect 1258 61529 534662 62343
rect 1258 61504 41853 61529
rect 1258 60775 5341 60800
rect 1258 59961 534662 60775
rect 1258 59936 22141 59961
rect 1258 59207 5117 59232
rect 1258 58393 534662 59207
rect 1258 58368 41069 58393
rect 1258 57639 5005 57664
rect 1258 56825 534662 57639
rect 1258 56800 10157 56825
rect 1258 56071 4781 56096
rect 1258 55257 534662 56071
rect 1258 55232 9821 55257
rect 1258 54503 4221 54528
rect 1258 53689 534662 54503
rect 1258 53664 22477 53689
rect 1258 52935 3997 52960
rect 1258 52121 534662 52935
rect 1258 52096 14749 52121
rect 1258 51367 33901 51392
rect 1258 50553 534662 51367
rect 1258 50528 8253 50553
rect 1258 49799 10381 49824
rect 1258 48985 534662 49799
rect 1258 48960 8701 48985
rect 1258 48231 14525 48256
rect 1258 47417 534662 48231
rect 1258 47392 25277 47417
rect 1258 46663 22589 46688
rect 1258 45849 534662 46663
rect 1258 45824 32333 45849
rect 1258 45095 15800 45120
rect 1258 44281 534662 45095
rect 1258 44256 42189 44281
rect 1258 43527 12733 43552
rect 1258 42713 534662 43527
rect 1258 42688 53501 42713
rect 1258 41959 61453 41984
rect 1258 41145 534662 41959
rect 1258 41120 15421 41145
rect 1258 40391 19901 40416
rect 1258 39577 534662 40391
rect 1258 39552 10717 39577
rect 1258 38823 5005 38848
rect 1258 38009 534662 38823
rect 1258 37984 15533 38009
rect 1258 37255 4557 37280
rect 1258 36441 534662 37255
rect 1258 36416 45661 36441
rect 1258 35687 6013 35712
rect 1258 34873 534662 35687
rect 1258 34848 6461 34873
rect 1258 34119 5229 34144
rect 1258 33305 534662 34119
rect 1258 33280 101885 33305
rect 1258 32551 45885 32576
rect 1258 31737 534662 32551
rect 1258 31712 8701 31737
rect 1258 30983 14749 31008
rect 1258 30169 534662 30983
rect 1258 30144 8701 30169
rect 1258 29415 22072 29440
rect 1258 28601 534662 29415
rect 1258 28576 101885 28601
rect 1258 27847 35021 27872
rect 1258 27033 534662 27847
rect 1258 27008 24157 27033
rect 1258 26279 43085 26304
rect 1258 25465 534662 26279
rect 1258 25440 6461 25465
rect 1258 24711 4781 24736
rect 1258 23897 534662 24711
rect 1258 23872 10829 23897
rect 1258 23143 4445 23168
rect 1258 22329 534662 23143
rect 1258 22304 26509 22329
rect 1258 21575 18221 21600
rect 1258 20761 534662 21575
rect 1258 20736 6461 20761
rect 1258 20007 5341 20032
rect 1258 19193 534662 20007
rect 1258 19168 18669 19193
rect 1258 18439 5341 18464
rect 1258 17625 534662 18439
rect 1258 17600 31773 17625
rect 1258 16871 26397 16896
rect 1258 16057 534662 16871
rect 1258 16032 25837 16057
rect 1258 15303 5789 15328
rect 1258 14489 534662 15303
rect 1258 14464 7512 14489
rect 1258 13735 58317 13760
rect 1258 12921 534662 13735
rect 1258 12896 24717 12921
rect 1258 12167 27517 12192
rect 1258 11353 534662 12167
rect 1258 11328 8141 11353
rect 1258 10599 10941 10624
rect 1258 9785 534662 10599
rect 1258 9760 40285 9785
rect 1258 9031 14301 9056
rect 1258 8217 534662 9031
rect 1258 8192 40509 8217
rect 1258 7463 66605 7488
rect 1258 6649 534662 7463
rect 1258 6624 65485 6649
rect 1258 5895 73773 5920
rect 1258 5081 534662 5895
rect 1258 5056 73437 5081
rect 1258 4327 82957 4352
rect 1258 3513 534662 4327
rect 1258 3488 203620 3513
<< pwell >>
rect 1258 175264 534662 175968
rect 1258 173696 534662 174400
rect 1258 172128 534662 172832
rect 1258 170560 534662 171264
rect 1258 168992 534662 169696
rect 1258 167424 534662 168128
rect 1258 165856 534662 166560
rect 1258 164288 534662 164992
rect 1258 162720 534662 163424
rect 1258 161152 534662 161856
rect 1258 159584 534662 160288
rect 1258 158016 534662 158720
rect 1258 156448 534662 157152
rect 1258 154880 534662 155584
rect 1258 153312 534662 154016
rect 1258 151744 534662 152448
rect 1258 150176 534662 150880
rect 1258 148608 534662 149312
rect 1258 147040 534662 147744
rect 1258 145472 534662 146176
rect 1258 143904 534662 144608
rect 1258 142336 534662 143040
rect 1258 140768 534662 141472
rect 1258 139200 534662 139904
rect 1258 137632 534662 138336
rect 1258 136064 534662 136768
rect 1258 134496 534662 135200
rect 1258 132928 534662 133632
rect 1258 131360 534662 132064
rect 1258 129792 534662 130496
rect 1258 128224 534662 128928
rect 1258 126656 534662 127360
rect 1258 125088 534662 125792
rect 1258 123520 534662 124224
rect 1258 121952 534662 122656
rect 1258 120384 534662 121088
rect 1258 118816 534662 119520
rect 1258 117248 534662 117952
rect 1258 115680 534662 116384
rect 1258 114112 534662 114816
rect 1258 112544 534662 113248
rect 1258 110976 534662 111680
rect 1258 109408 534662 110112
rect 1258 107840 534662 108544
rect 1258 106272 534662 106976
rect 1258 104704 534662 105408
rect 1258 103136 534662 103840
rect 1258 101568 534662 102272
rect 1258 100000 534662 100704
rect 1258 98432 534662 99136
rect 1258 96864 534662 97568
rect 1258 95296 534662 96000
rect 1258 93728 534662 94432
rect 1258 92160 534662 92864
rect 1258 90592 534662 91296
rect 1258 89024 534662 89728
rect 1258 87456 534662 88160
rect 1258 85888 534662 86592
rect 1258 84320 534662 85024
rect 1258 82752 534662 83456
rect 1258 81184 534662 81888
rect 1258 79616 534662 80320
rect 1258 78048 534662 78752
rect 1258 76480 534662 77184
rect 1258 74912 534662 75616
rect 1258 73344 534662 74048
rect 1258 71776 534662 72480
rect 1258 70208 534662 70912
rect 1258 68640 534662 69344
rect 1258 67072 534662 67776
rect 1258 65504 534662 66208
rect 1258 63936 534662 64640
rect 1258 62368 534662 63072
rect 1258 60800 534662 61504
rect 1258 59232 534662 59936
rect 1258 57664 534662 58368
rect 1258 56096 534662 56800
rect 1258 54528 534662 55232
rect 1258 52960 534662 53664
rect 1258 51392 534662 52096
rect 1258 49824 534662 50528
rect 1258 48256 534662 48960
rect 1258 46688 534662 47392
rect 1258 45120 534662 45824
rect 1258 43552 534662 44256
rect 1258 41984 534662 42688
rect 1258 40416 534662 41120
rect 1258 38848 534662 39552
rect 1258 37280 534662 37984
rect 1258 35712 534662 36416
rect 1258 34144 534662 34848
rect 1258 32576 534662 33280
rect 1258 31008 534662 31712
rect 1258 29440 534662 30144
rect 1258 27872 534662 28576
rect 1258 26304 534662 27008
rect 1258 24736 534662 25440
rect 1258 23168 534662 23872
rect 1258 21600 534662 22304
rect 1258 20032 534662 20736
rect 1258 18464 534662 19168
rect 1258 16896 534662 17600
rect 1258 15328 534662 16032
rect 1258 13760 534662 14464
rect 1258 12192 534662 12896
rect 1258 10624 534662 11328
rect 1258 9056 534662 9760
rect 1258 7488 534662 8192
rect 1258 5920 534662 6624
rect 1258 4352 534662 5056
rect 1258 3050 534662 3488
<< obsm1 >>
rect 1344 3076 534576 176460
<< metal2 >>
rect 9856 0 9968 800
rect 13888 0 14000 800
rect 17920 0 18032 800
rect 21952 0 22064 800
rect 25984 0 26096 800
rect 30016 0 30128 800
rect 34048 0 34160 800
rect 38080 0 38192 800
rect 42112 0 42224 800
rect 46144 0 46256 800
rect 50176 0 50288 800
rect 54208 0 54320 800
rect 58240 0 58352 800
rect 62272 0 62384 800
rect 66304 0 66416 800
rect 70336 0 70448 800
rect 74368 0 74480 800
rect 78400 0 78512 800
rect 82432 0 82544 800
rect 86464 0 86576 800
rect 90496 0 90608 800
rect 94528 0 94640 800
rect 98560 0 98672 800
rect 102592 0 102704 800
rect 106624 0 106736 800
rect 110656 0 110768 800
rect 114688 0 114800 800
rect 118720 0 118832 800
rect 122752 0 122864 800
rect 126784 0 126896 800
rect 130816 0 130928 800
rect 134848 0 134960 800
rect 138880 0 138992 800
rect 142912 0 143024 800
rect 146944 0 147056 800
rect 150976 0 151088 800
rect 155008 0 155120 800
rect 159040 0 159152 800
rect 163072 0 163184 800
rect 167104 0 167216 800
rect 171136 0 171248 800
rect 175168 0 175280 800
rect 179200 0 179312 800
rect 183232 0 183344 800
rect 187264 0 187376 800
rect 191296 0 191408 800
rect 195328 0 195440 800
rect 199360 0 199472 800
rect 203392 0 203504 800
rect 207424 0 207536 800
rect 211456 0 211568 800
rect 215488 0 215600 800
rect 219520 0 219632 800
rect 223552 0 223664 800
rect 227584 0 227696 800
rect 231616 0 231728 800
rect 235648 0 235760 800
rect 239680 0 239792 800
rect 243712 0 243824 800
rect 247744 0 247856 800
rect 251776 0 251888 800
rect 255808 0 255920 800
rect 259840 0 259952 800
rect 263872 0 263984 800
rect 267904 0 268016 800
rect 271936 0 272048 800
rect 275968 0 276080 800
rect 280000 0 280112 800
rect 284032 0 284144 800
rect 288064 0 288176 800
rect 292096 0 292208 800
rect 296128 0 296240 800
rect 300160 0 300272 800
rect 304192 0 304304 800
rect 308224 0 308336 800
rect 312256 0 312368 800
rect 316288 0 316400 800
rect 320320 0 320432 800
rect 324352 0 324464 800
rect 328384 0 328496 800
rect 332416 0 332528 800
rect 336448 0 336560 800
rect 340480 0 340592 800
rect 344512 0 344624 800
rect 348544 0 348656 800
rect 352576 0 352688 800
rect 356608 0 356720 800
rect 360640 0 360752 800
rect 364672 0 364784 800
rect 368704 0 368816 800
rect 372736 0 372848 800
rect 376768 0 376880 800
rect 380800 0 380912 800
rect 384832 0 384944 800
rect 388864 0 388976 800
rect 392896 0 393008 800
rect 396928 0 397040 800
rect 400960 0 401072 800
rect 404992 0 405104 800
rect 409024 0 409136 800
rect 413056 0 413168 800
rect 417088 0 417200 800
rect 421120 0 421232 800
rect 425152 0 425264 800
rect 429184 0 429296 800
rect 433216 0 433328 800
rect 437248 0 437360 800
rect 441280 0 441392 800
rect 445312 0 445424 800
rect 449344 0 449456 800
rect 453376 0 453488 800
rect 457408 0 457520 800
rect 461440 0 461552 800
rect 465472 0 465584 800
rect 469504 0 469616 800
rect 473536 0 473648 800
rect 477568 0 477680 800
rect 481600 0 481712 800
rect 485632 0 485744 800
rect 489664 0 489776 800
rect 493696 0 493808 800
rect 497728 0 497840 800
rect 501760 0 501872 800
rect 505792 0 505904 800
rect 509824 0 509936 800
rect 513856 0 513968 800
rect 517888 0 518000 800
rect 521920 0 522032 800
rect 525952 0 526064 800
<< obsm2 >>
rect 3276 860 533764 178958
rect 3276 466 9796 860
rect 10028 466 13828 860
rect 14060 466 17860 860
rect 18092 466 21892 860
rect 22124 466 25924 860
rect 26156 466 29956 860
rect 30188 466 33988 860
rect 34220 466 38020 860
rect 38252 466 42052 860
rect 42284 466 46084 860
rect 46316 466 50116 860
rect 50348 466 54148 860
rect 54380 466 58180 860
rect 58412 466 62212 860
rect 62444 466 66244 860
rect 66476 466 70276 860
rect 70508 466 74308 860
rect 74540 466 78340 860
rect 78572 466 82372 860
rect 82604 466 86404 860
rect 86636 466 90436 860
rect 90668 466 94468 860
rect 94700 466 98500 860
rect 98732 466 102532 860
rect 102764 466 106564 860
rect 106796 466 110596 860
rect 110828 466 114628 860
rect 114860 466 118660 860
rect 118892 466 122692 860
rect 122924 466 126724 860
rect 126956 466 130756 860
rect 130988 466 134788 860
rect 135020 466 138820 860
rect 139052 466 142852 860
rect 143084 466 146884 860
rect 147116 466 150916 860
rect 151148 466 154948 860
rect 155180 466 158980 860
rect 159212 466 163012 860
rect 163244 466 167044 860
rect 167276 466 171076 860
rect 171308 466 175108 860
rect 175340 466 179140 860
rect 179372 466 183172 860
rect 183404 466 187204 860
rect 187436 466 191236 860
rect 191468 466 195268 860
rect 195500 466 199300 860
rect 199532 466 203332 860
rect 203564 466 207364 860
rect 207596 466 211396 860
rect 211628 466 215428 860
rect 215660 466 219460 860
rect 219692 466 223492 860
rect 223724 466 227524 860
rect 227756 466 231556 860
rect 231788 466 235588 860
rect 235820 466 239620 860
rect 239852 466 243652 860
rect 243884 466 247684 860
rect 247916 466 251716 860
rect 251948 466 255748 860
rect 255980 466 259780 860
rect 260012 466 263812 860
rect 264044 466 267844 860
rect 268076 466 271876 860
rect 272108 466 275908 860
rect 276140 466 279940 860
rect 280172 466 283972 860
rect 284204 466 288004 860
rect 288236 466 292036 860
rect 292268 466 296068 860
rect 296300 466 300100 860
rect 300332 466 304132 860
rect 304364 466 308164 860
rect 308396 466 312196 860
rect 312428 466 316228 860
rect 316460 466 320260 860
rect 320492 466 324292 860
rect 324524 466 328324 860
rect 328556 466 332356 860
rect 332588 466 336388 860
rect 336620 466 340420 860
rect 340652 466 344452 860
rect 344684 466 348484 860
rect 348716 466 352516 860
rect 352748 466 356548 860
rect 356780 466 360580 860
rect 360812 466 364612 860
rect 364844 466 368644 860
rect 368876 466 372676 860
rect 372908 466 376708 860
rect 376940 466 380740 860
rect 380972 466 384772 860
rect 385004 466 388804 860
rect 389036 466 392836 860
rect 393068 466 396868 860
rect 397100 466 400900 860
rect 401132 466 404932 860
rect 405164 466 408964 860
rect 409196 466 412996 860
rect 413228 466 417028 860
rect 417260 466 421060 860
rect 421292 466 425092 860
rect 425324 466 429124 860
rect 429356 466 433156 860
rect 433388 466 437188 860
rect 437420 466 441220 860
rect 441452 466 445252 860
rect 445484 466 449284 860
rect 449516 466 453316 860
rect 453548 466 457348 860
rect 457580 466 461380 860
rect 461612 466 465412 860
rect 465644 466 469444 860
rect 469676 466 473476 860
rect 473708 466 477508 860
rect 477740 466 481540 860
rect 481772 466 485572 860
rect 485804 466 489604 860
rect 489836 466 493636 860
rect 493868 466 497668 860
rect 497900 466 501700 860
rect 501932 466 505732 860
rect 505964 466 509764 860
rect 509996 466 513796 860
rect 514028 466 517828 860
rect 518060 466 521860 860
rect 522092 466 525892 860
rect 526124 466 533764 860
<< obsm3 >>
rect 3378 364 533774 178948
<< metal4 >>
rect 4448 3076 4768 176460
rect 19808 3076 20128 176460
rect 35168 3076 35488 176460
rect 50528 3076 50848 176460
rect 65888 3076 66208 176460
rect 81248 3076 81568 176460
rect 96608 3076 96928 176460
rect 111968 3076 112288 176460
rect 127328 3076 127648 176460
rect 142688 3076 143008 176460
rect 158048 3076 158368 176460
rect 173408 3076 173728 176460
rect 188768 3076 189088 176460
rect 204128 3076 204448 176460
rect 219488 3076 219808 176460
rect 234848 3076 235168 176460
rect 250208 3076 250528 176460
rect 265568 3076 265888 176460
rect 280928 3076 281248 176460
rect 296288 3076 296608 176460
rect 311648 3076 311968 176460
rect 327008 3076 327328 176460
rect 342368 3076 342688 176460
rect 357728 3076 358048 176460
rect 373088 3076 373408 176460
rect 388448 3076 388768 176460
rect 403808 3076 404128 176460
rect 419168 3076 419488 176460
rect 434528 3076 434848 176460
rect 449888 3076 450208 176460
rect 465248 3076 465568 176460
rect 480608 3076 480928 176460
rect 495968 3076 496288 176460
rect 511328 3076 511648 176460
rect 526688 3076 527008 176460
<< obsm4 >>
rect 11676 176520 529172 178734
rect 11676 3016 19748 176520
rect 20188 3016 35108 176520
rect 35548 3016 50468 176520
rect 50908 3016 65828 176520
rect 66268 3016 81188 176520
rect 81628 3016 96548 176520
rect 96988 3016 111908 176520
rect 112348 3016 127268 176520
rect 127708 3016 142628 176520
rect 143068 3016 157988 176520
rect 158428 3016 173348 176520
rect 173788 3016 188708 176520
rect 189148 3016 204068 176520
rect 204508 3016 219428 176520
rect 219868 3016 234788 176520
rect 235228 3016 250148 176520
rect 250588 3016 265508 176520
rect 265948 3016 280868 176520
rect 281308 3016 296228 176520
rect 296668 3016 311588 176520
rect 312028 3016 326948 176520
rect 327388 3016 342308 176520
rect 342748 3016 357668 176520
rect 358108 3016 373028 176520
rect 373468 3016 388388 176520
rect 388828 3016 403748 176520
rect 404188 3016 419108 176520
rect 419548 3016 434468 176520
rect 434908 3016 449828 176520
rect 450268 3016 465188 176520
rect 465628 3016 480548 176520
rect 480988 3016 495908 176520
rect 496348 3016 511268 176520
rect 511708 3016 526628 176520
rect 527068 3016 529172 176520
rect 11676 354 529172 3016
<< labels >>
rlabel metal2 s 9856 0 9968 800 6 i_clk
port 1 nsew signal input
rlabel metal2 s 13888 0 14000 800 6 i_rst
port 2 nsew signal input
rlabel metal2 s 17920 0 18032 800 6 mem_ack
port 3 nsew signal output
rlabel metal2 s 62272 0 62384 800 6 mem_addr[0]
port 4 nsew signal input
rlabel metal2 s 320320 0 320432 800 6 mem_addr[10]
port 5 nsew signal input
rlabel metal2 s 344512 0 344624 800 6 mem_addr[11]
port 6 nsew signal input
rlabel metal2 s 368704 0 368816 800 6 mem_addr[12]
port 7 nsew signal input
rlabel metal2 s 392896 0 393008 800 6 mem_addr[13]
port 8 nsew signal input
rlabel metal2 s 417088 0 417200 800 6 mem_addr[14]
port 9 nsew signal input
rlabel metal2 s 441280 0 441392 800 6 mem_addr[15]
port 10 nsew signal input
rlabel metal2 s 465472 0 465584 800 6 mem_addr[16]
port 11 nsew signal input
rlabel metal2 s 473536 0 473648 800 6 mem_addr[17]
port 12 nsew signal input
rlabel metal2 s 481600 0 481712 800 6 mem_addr[18]
port 13 nsew signal input
rlabel metal2 s 489664 0 489776 800 6 mem_addr[19]
port 14 nsew signal input
rlabel metal2 s 94528 0 94640 800 6 mem_addr[1]
port 15 nsew signal input
rlabel metal2 s 497728 0 497840 800 6 mem_addr[20]
port 16 nsew signal input
rlabel metal2 s 505792 0 505904 800 6 mem_addr[21]
port 17 nsew signal input
rlabel metal2 s 513856 0 513968 800 6 mem_addr[22]
port 18 nsew signal input
rlabel metal2 s 521920 0 522032 800 6 mem_addr[23]
port 19 nsew signal input
rlabel metal2 s 126784 0 126896 800 6 mem_addr[2]
port 20 nsew signal input
rlabel metal2 s 150976 0 151088 800 6 mem_addr[3]
port 21 nsew signal input
rlabel metal2 s 175168 0 175280 800 6 mem_addr[4]
port 22 nsew signal input
rlabel metal2 s 199360 0 199472 800 6 mem_addr[5]
port 23 nsew signal input
rlabel metal2 s 223552 0 223664 800 6 mem_addr[6]
port 24 nsew signal input
rlabel metal2 s 247744 0 247856 800 6 mem_addr[7]
port 25 nsew signal input
rlabel metal2 s 271936 0 272048 800 6 mem_addr[8]
port 26 nsew signal input
rlabel metal2 s 296128 0 296240 800 6 mem_addr[9]
port 27 nsew signal input
rlabel metal2 s 21952 0 22064 800 6 mem_cache_enable
port 28 nsew signal input
rlabel metal2 s 25984 0 26096 800 6 mem_exception
port 29 nsew signal output
rlabel metal2 s 66304 0 66416 800 6 mem_i_data[0]
port 30 nsew signal input
rlabel metal2 s 324352 0 324464 800 6 mem_i_data[10]
port 31 nsew signal input
rlabel metal2 s 348544 0 348656 800 6 mem_i_data[11]
port 32 nsew signal input
rlabel metal2 s 372736 0 372848 800 6 mem_i_data[12]
port 33 nsew signal input
rlabel metal2 s 396928 0 397040 800 6 mem_i_data[13]
port 34 nsew signal input
rlabel metal2 s 421120 0 421232 800 6 mem_i_data[14]
port 35 nsew signal input
rlabel metal2 s 445312 0 445424 800 6 mem_i_data[15]
port 36 nsew signal input
rlabel metal2 s 98560 0 98672 800 6 mem_i_data[1]
port 37 nsew signal input
rlabel metal2 s 130816 0 130928 800 6 mem_i_data[2]
port 38 nsew signal input
rlabel metal2 s 155008 0 155120 800 6 mem_i_data[3]
port 39 nsew signal input
rlabel metal2 s 179200 0 179312 800 6 mem_i_data[4]
port 40 nsew signal input
rlabel metal2 s 203392 0 203504 800 6 mem_i_data[5]
port 41 nsew signal input
rlabel metal2 s 227584 0 227696 800 6 mem_i_data[6]
port 42 nsew signal input
rlabel metal2 s 251776 0 251888 800 6 mem_i_data[7]
port 43 nsew signal input
rlabel metal2 s 275968 0 276080 800 6 mem_i_data[8]
port 44 nsew signal input
rlabel metal2 s 300160 0 300272 800 6 mem_i_data[9]
port 45 nsew signal input
rlabel metal2 s 70336 0 70448 800 6 mem_o_data[0]
port 46 nsew signal output
rlabel metal2 s 328384 0 328496 800 6 mem_o_data[10]
port 47 nsew signal output
rlabel metal2 s 352576 0 352688 800 6 mem_o_data[11]
port 48 nsew signal output
rlabel metal2 s 376768 0 376880 800 6 mem_o_data[12]
port 49 nsew signal output
rlabel metal2 s 400960 0 401072 800 6 mem_o_data[13]
port 50 nsew signal output
rlabel metal2 s 425152 0 425264 800 6 mem_o_data[14]
port 51 nsew signal output
rlabel metal2 s 449344 0 449456 800 6 mem_o_data[15]
port 52 nsew signal output
rlabel metal2 s 102592 0 102704 800 6 mem_o_data[1]
port 53 nsew signal output
rlabel metal2 s 134848 0 134960 800 6 mem_o_data[2]
port 54 nsew signal output
rlabel metal2 s 159040 0 159152 800 6 mem_o_data[3]
port 55 nsew signal output
rlabel metal2 s 183232 0 183344 800 6 mem_o_data[4]
port 56 nsew signal output
rlabel metal2 s 207424 0 207536 800 6 mem_o_data[5]
port 57 nsew signal output
rlabel metal2 s 231616 0 231728 800 6 mem_o_data[6]
port 58 nsew signal output
rlabel metal2 s 255808 0 255920 800 6 mem_o_data[7]
port 59 nsew signal output
rlabel metal2 s 280000 0 280112 800 6 mem_o_data[8]
port 60 nsew signal output
rlabel metal2 s 304192 0 304304 800 6 mem_o_data[9]
port 61 nsew signal output
rlabel metal2 s 30016 0 30128 800 6 mem_req
port 62 nsew signal input
rlabel metal2 s 74368 0 74480 800 6 mem_sel[0]
port 63 nsew signal input
rlabel metal2 s 106624 0 106736 800 6 mem_sel[1]
port 64 nsew signal input
rlabel metal2 s 34048 0 34160 800 6 mem_we
port 65 nsew signal input
rlabel metal4 s 4448 3076 4768 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 219488 3076 219808 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 250208 3076 250528 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 280928 3076 281248 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 311648 3076 311968 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 342368 3076 342688 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 373088 3076 373408 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 403808 3076 404128 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 434528 3076 434848 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 465248 3076 465568 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 495968 3076 496288 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 526688 3076 527008 176460 6 vccd1
port 66 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 234848 3076 235168 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 265568 3076 265888 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 296288 3076 296608 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 327008 3076 327328 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 357728 3076 358048 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 388448 3076 388768 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 419168 3076 419488 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 449888 3076 450208 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 480608 3076 480928 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal4 s 511328 3076 511648 176460 6 vssd1
port 67 nsew ground bidirectional
rlabel metal2 s 38080 0 38192 800 6 wb_4_burst
port 68 nsew signal output
rlabel metal2 s 42112 0 42224 800 6 wb_ack
port 69 nsew signal input
rlabel metal2 s 78400 0 78512 800 6 wb_adr[0]
port 70 nsew signal output
rlabel metal2 s 332416 0 332528 800 6 wb_adr[10]
port 71 nsew signal output
rlabel metal2 s 356608 0 356720 800 6 wb_adr[11]
port 72 nsew signal output
rlabel metal2 s 380800 0 380912 800 6 wb_adr[12]
port 73 nsew signal output
rlabel metal2 s 404992 0 405104 800 6 wb_adr[13]
port 74 nsew signal output
rlabel metal2 s 429184 0 429296 800 6 wb_adr[14]
port 75 nsew signal output
rlabel metal2 s 453376 0 453488 800 6 wb_adr[15]
port 76 nsew signal output
rlabel metal2 s 469504 0 469616 800 6 wb_adr[16]
port 77 nsew signal output
rlabel metal2 s 477568 0 477680 800 6 wb_adr[17]
port 78 nsew signal output
rlabel metal2 s 485632 0 485744 800 6 wb_adr[18]
port 79 nsew signal output
rlabel metal2 s 493696 0 493808 800 6 wb_adr[19]
port 80 nsew signal output
rlabel metal2 s 110656 0 110768 800 6 wb_adr[1]
port 81 nsew signal output
rlabel metal2 s 501760 0 501872 800 6 wb_adr[20]
port 82 nsew signal output
rlabel metal2 s 509824 0 509936 800 6 wb_adr[21]
port 83 nsew signal output
rlabel metal2 s 517888 0 518000 800 6 wb_adr[22]
port 84 nsew signal output
rlabel metal2 s 525952 0 526064 800 6 wb_adr[23]
port 85 nsew signal output
rlabel metal2 s 138880 0 138992 800 6 wb_adr[2]
port 86 nsew signal output
rlabel metal2 s 163072 0 163184 800 6 wb_adr[3]
port 87 nsew signal output
rlabel metal2 s 187264 0 187376 800 6 wb_adr[4]
port 88 nsew signal output
rlabel metal2 s 211456 0 211568 800 6 wb_adr[5]
port 89 nsew signal output
rlabel metal2 s 235648 0 235760 800 6 wb_adr[6]
port 90 nsew signal output
rlabel metal2 s 259840 0 259952 800 6 wb_adr[7]
port 91 nsew signal output
rlabel metal2 s 284032 0 284144 800 6 wb_adr[8]
port 92 nsew signal output
rlabel metal2 s 308224 0 308336 800 6 wb_adr[9]
port 93 nsew signal output
rlabel metal2 s 46144 0 46256 800 6 wb_cyc
port 94 nsew signal output
rlabel metal2 s 50176 0 50288 800 6 wb_err
port 95 nsew signal input
rlabel metal2 s 82432 0 82544 800 6 wb_i_dat[0]
port 96 nsew signal input
rlabel metal2 s 336448 0 336560 800 6 wb_i_dat[10]
port 97 nsew signal input
rlabel metal2 s 360640 0 360752 800 6 wb_i_dat[11]
port 98 nsew signal input
rlabel metal2 s 384832 0 384944 800 6 wb_i_dat[12]
port 99 nsew signal input
rlabel metal2 s 409024 0 409136 800 6 wb_i_dat[13]
port 100 nsew signal input
rlabel metal2 s 433216 0 433328 800 6 wb_i_dat[14]
port 101 nsew signal input
rlabel metal2 s 457408 0 457520 800 6 wb_i_dat[15]
port 102 nsew signal input
rlabel metal2 s 114688 0 114800 800 6 wb_i_dat[1]
port 103 nsew signal input
rlabel metal2 s 142912 0 143024 800 6 wb_i_dat[2]
port 104 nsew signal input
rlabel metal2 s 167104 0 167216 800 6 wb_i_dat[3]
port 105 nsew signal input
rlabel metal2 s 191296 0 191408 800 6 wb_i_dat[4]
port 106 nsew signal input
rlabel metal2 s 215488 0 215600 800 6 wb_i_dat[5]
port 107 nsew signal input
rlabel metal2 s 239680 0 239792 800 6 wb_i_dat[6]
port 108 nsew signal input
rlabel metal2 s 263872 0 263984 800 6 wb_i_dat[7]
port 109 nsew signal input
rlabel metal2 s 288064 0 288176 800 6 wb_i_dat[8]
port 110 nsew signal input
rlabel metal2 s 312256 0 312368 800 6 wb_i_dat[9]
port 111 nsew signal input
rlabel metal2 s 86464 0 86576 800 6 wb_o_dat[0]
port 112 nsew signal output
rlabel metal2 s 340480 0 340592 800 6 wb_o_dat[10]
port 113 nsew signal output
rlabel metal2 s 364672 0 364784 800 6 wb_o_dat[11]
port 114 nsew signal output
rlabel metal2 s 388864 0 388976 800 6 wb_o_dat[12]
port 115 nsew signal output
rlabel metal2 s 413056 0 413168 800 6 wb_o_dat[13]
port 116 nsew signal output
rlabel metal2 s 437248 0 437360 800 6 wb_o_dat[14]
port 117 nsew signal output
rlabel metal2 s 461440 0 461552 800 6 wb_o_dat[15]
port 118 nsew signal output
rlabel metal2 s 118720 0 118832 800 6 wb_o_dat[1]
port 119 nsew signal output
rlabel metal2 s 146944 0 147056 800 6 wb_o_dat[2]
port 120 nsew signal output
rlabel metal2 s 171136 0 171248 800 6 wb_o_dat[3]
port 121 nsew signal output
rlabel metal2 s 195328 0 195440 800 6 wb_o_dat[4]
port 122 nsew signal output
rlabel metal2 s 219520 0 219632 800 6 wb_o_dat[5]
port 123 nsew signal output
rlabel metal2 s 243712 0 243824 800 6 wb_o_dat[6]
port 124 nsew signal output
rlabel metal2 s 267904 0 268016 800 6 wb_o_dat[7]
port 125 nsew signal output
rlabel metal2 s 292096 0 292208 800 6 wb_o_dat[8]
port 126 nsew signal output
rlabel metal2 s 316288 0 316400 800 6 wb_o_dat[9]
port 127 nsew signal output
rlabel metal2 s 90496 0 90608 800 6 wb_sel[0]
port 128 nsew signal output
rlabel metal2 s 122752 0 122864 800 6 wb_sel[1]
port 129 nsew signal output
rlabel metal2 s 54208 0 54320 800 6 wb_stb
port 130 nsew signal output
rlabel metal2 s 58240 0 58352 800 6 wb_we
port 131 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 536000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 66294626
string GDS_FILE /home/piotro/caravel_user_project/openlane/dcache/runs/23_11_16_01_38/results/signoff/dcache.magic.gds
string GDS_START 469046
<< end >>

