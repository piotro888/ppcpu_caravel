magic
tech sky130B
magscale 1 2
timestamp 1663051489
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 14 2128 29702 27792
<< metal2 >>
rect 18 29200 74 30000
rect 662 29200 718 30000
rect 1306 29200 1362 30000
rect 1950 29200 2006 30000
rect 2594 29200 2650 30000
rect 3238 29200 3294 30000
rect 3882 29200 3938 30000
rect 4526 29200 4582 30000
rect 5170 29200 5226 30000
rect 5814 29200 5870 30000
rect 6458 29200 6514 30000
rect 7102 29200 7158 30000
rect 7746 29200 7802 30000
rect 8390 29200 8446 30000
rect 9034 29200 9090 30000
rect 9678 29200 9734 30000
rect 10966 29200 11022 30000
rect 11610 29200 11666 30000
rect 12254 29200 12310 30000
rect 12898 29200 12954 30000
rect 13542 29200 13598 30000
rect 14186 29200 14242 30000
rect 14830 29200 14886 30000
rect 15474 29200 15530 30000
rect 16118 29200 16174 30000
rect 16762 29200 16818 30000
rect 17406 29200 17462 30000
rect 18050 29200 18106 30000
rect 18694 29200 18750 30000
rect 19338 29200 19394 30000
rect 19982 29200 20038 30000
rect 20626 29200 20682 30000
rect 21270 29200 21326 30000
rect 21914 29200 21970 30000
rect 22558 29200 22614 30000
rect 23202 29200 23258 30000
rect 23846 29200 23902 30000
rect 24490 29200 24546 30000
rect 25134 29200 25190 30000
rect 25778 29200 25834 30000
rect 26422 29200 26478 30000
rect 27066 29200 27122 30000
rect 27710 29200 27766 30000
rect 28354 29200 28410 30000
rect 28998 29200 29054 30000
rect 29642 29200 29698 30000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
<< obsm2 >>
rect 130 29144 606 29345
rect 774 29144 1250 29345
rect 1418 29144 1894 29345
rect 2062 29144 2538 29345
rect 2706 29144 3182 29345
rect 3350 29144 3826 29345
rect 3994 29144 4470 29345
rect 4638 29144 5114 29345
rect 5282 29144 5758 29345
rect 5926 29144 6402 29345
rect 6570 29144 7046 29345
rect 7214 29144 7690 29345
rect 7858 29144 8334 29345
rect 8502 29144 8978 29345
rect 9146 29144 9622 29345
rect 9790 29144 10910 29345
rect 11078 29144 11554 29345
rect 11722 29144 12198 29345
rect 12366 29144 12842 29345
rect 13010 29144 13486 29345
rect 13654 29144 14130 29345
rect 14298 29144 14774 29345
rect 14942 29144 15418 29345
rect 15586 29144 16062 29345
rect 16230 29144 16706 29345
rect 16874 29144 17350 29345
rect 17518 29144 17994 29345
rect 18162 29144 18638 29345
rect 18806 29144 19282 29345
rect 19450 29144 19926 29345
rect 20094 29144 20570 29345
rect 20738 29144 21214 29345
rect 21382 29144 21858 29345
rect 22026 29144 22502 29345
rect 22670 29144 23146 29345
rect 23314 29144 23790 29345
rect 23958 29144 24434 29345
rect 24602 29144 25078 29345
rect 25246 29144 25722 29345
rect 25890 29144 26366 29345
rect 26534 29144 27010 29345
rect 27178 29144 27654 29345
rect 27822 29144 28298 29345
rect 28466 29144 28942 29345
rect 29110 29144 29586 29345
rect 20 856 29696 29144
rect 130 31 606 856
rect 774 31 1250 856
rect 1418 31 1894 856
rect 2062 31 2538 856
rect 2706 31 3182 856
rect 3350 31 3826 856
rect 3994 31 4470 856
rect 4638 31 5114 856
rect 5282 31 5758 856
rect 5926 31 6402 856
rect 6570 31 7046 856
rect 7214 31 7690 856
rect 7858 31 8334 856
rect 8502 31 8978 856
rect 9146 31 9622 856
rect 9790 31 10266 856
rect 10434 31 10910 856
rect 11078 31 11554 856
rect 11722 31 12198 856
rect 12366 31 12842 856
rect 13010 31 13486 856
rect 13654 31 14130 856
rect 14298 31 14774 856
rect 14942 31 15418 856
rect 15586 31 16062 856
rect 16230 31 16706 856
rect 16874 31 17350 856
rect 17518 31 17994 856
rect 18162 31 18638 856
rect 18806 31 19282 856
rect 19450 31 19926 856
rect 20094 31 20570 856
rect 20738 31 21214 856
rect 21382 31 21858 856
rect 22026 31 22502 856
rect 22670 31 23146 856
rect 23314 31 23790 856
rect 23958 31 24434 856
rect 24602 31 25078 856
rect 25246 31 25722 856
rect 25890 31 26366 856
rect 26534 31 27010 856
rect 27178 31 27654 856
rect 27822 31 28298 856
rect 28466 31 28942 856
rect 29110 31 29586 856
<< metal3 >>
rect 0 29248 800 29368
rect 29200 29248 30000 29368
rect 0 28568 800 28688
rect 29200 28568 30000 28688
rect 0 27888 800 28008
rect 29200 27888 30000 28008
rect 0 27208 800 27328
rect 29200 27208 30000 27328
rect 0 26528 800 26648
rect 29200 26528 30000 26648
rect 0 25848 800 25968
rect 29200 25848 30000 25968
rect 0 25168 800 25288
rect 29200 25168 30000 25288
rect 0 24488 800 24608
rect 29200 24488 30000 24608
rect 0 23808 800 23928
rect 29200 23808 30000 23928
rect 0 23128 800 23248
rect 29200 23128 30000 23248
rect 0 22448 800 22568
rect 29200 22448 30000 22568
rect 0 21768 800 21888
rect 29200 21768 30000 21888
rect 0 21088 800 21208
rect 29200 21088 30000 21208
rect 0 20408 800 20528
rect 29200 20408 30000 20528
rect 0 19728 800 19848
rect 29200 19728 30000 19848
rect 0 19048 800 19168
rect 29200 19048 30000 19168
rect 0 18368 800 18488
rect 29200 18368 30000 18488
rect 0 17688 800 17808
rect 29200 17688 30000 17808
rect 0 17008 800 17128
rect 29200 17008 30000 17128
rect 0 16328 800 16448
rect 29200 16328 30000 16448
rect 0 15648 800 15768
rect 29200 15648 30000 15768
rect 0 14968 800 15088
rect 29200 14968 30000 15088
rect 0 14288 800 14408
rect 29200 14288 30000 14408
rect 0 13608 800 13728
rect 29200 13608 30000 13728
rect 0 12928 800 13048
rect 29200 12928 30000 13048
rect 0 12248 800 12368
rect 29200 12248 30000 12368
rect 0 11568 800 11688
rect 29200 11568 30000 11688
rect 0 10888 800 11008
rect 29200 10888 30000 11008
rect 0 10208 800 10328
rect 29200 10208 30000 10328
rect 0 9528 800 9648
rect 29200 9528 30000 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 29200 8168 30000 8288
rect 0 7488 800 7608
rect 29200 7488 30000 7608
rect 0 6808 800 6928
rect 29200 6808 30000 6928
rect 0 6128 800 6248
rect 29200 6128 30000 6248
rect 0 5448 800 5568
rect 29200 5448 30000 5568
rect 0 4768 800 4888
rect 29200 4768 30000 4888
rect 0 4088 800 4208
rect 29200 4088 30000 4208
rect 0 3408 800 3528
rect 29200 3408 30000 3528
rect 0 2728 800 2848
rect 29200 2728 30000 2848
rect 0 2048 800 2168
rect 29200 2048 30000 2168
rect 0 1368 800 1488
rect 29200 1368 30000 1488
rect 0 688 800 808
rect 29200 688 30000 808
rect 29200 8 30000 128
<< obsm3 >>
rect 880 29168 29120 29341
rect 800 28768 29200 29168
rect 880 28488 29120 28768
rect 800 28088 29200 28488
rect 880 27808 29120 28088
rect 800 27408 29200 27808
rect 880 27128 29120 27408
rect 800 26728 29200 27128
rect 880 26448 29120 26728
rect 800 26048 29200 26448
rect 880 25768 29120 26048
rect 800 25368 29200 25768
rect 880 25088 29120 25368
rect 800 24688 29200 25088
rect 880 24408 29120 24688
rect 800 24008 29200 24408
rect 880 23728 29120 24008
rect 800 23328 29200 23728
rect 880 23048 29120 23328
rect 800 22648 29200 23048
rect 880 22368 29120 22648
rect 800 21968 29200 22368
rect 880 21688 29120 21968
rect 800 21288 29200 21688
rect 880 21008 29120 21288
rect 800 20608 29200 21008
rect 880 20328 29120 20608
rect 800 19928 29200 20328
rect 880 19648 29120 19928
rect 800 19248 29200 19648
rect 880 18968 29120 19248
rect 800 18568 29200 18968
rect 880 18288 29120 18568
rect 800 17888 29200 18288
rect 880 17608 29120 17888
rect 800 17208 29200 17608
rect 880 16928 29120 17208
rect 800 16528 29200 16928
rect 880 16248 29120 16528
rect 800 15848 29200 16248
rect 880 15568 29120 15848
rect 800 15168 29200 15568
rect 880 14888 29120 15168
rect 800 14488 29200 14888
rect 880 14208 29120 14488
rect 800 13808 29200 14208
rect 880 13528 29120 13808
rect 800 13128 29200 13528
rect 880 12848 29120 13128
rect 800 12448 29200 12848
rect 880 12168 29120 12448
rect 800 11768 29200 12168
rect 880 11488 29120 11768
rect 800 11088 29200 11488
rect 880 10808 29120 11088
rect 800 10408 29200 10808
rect 880 10128 29120 10408
rect 800 9728 29200 10128
rect 880 9448 29120 9728
rect 800 9048 29200 9448
rect 880 8768 29200 9048
rect 800 8368 29200 8768
rect 880 8088 29120 8368
rect 800 7688 29200 8088
rect 880 7408 29120 7688
rect 800 7008 29200 7408
rect 880 6728 29120 7008
rect 800 6328 29200 6728
rect 880 6048 29120 6328
rect 800 5648 29200 6048
rect 880 5368 29120 5648
rect 800 4968 29200 5368
rect 880 4688 29120 4968
rect 800 4288 29200 4688
rect 880 4008 29120 4288
rect 800 3608 29200 4008
rect 880 3328 29120 3608
rect 800 2928 29200 3328
rect 880 2648 29120 2928
rect 800 2248 29200 2648
rect 880 1968 29120 2248
rect 800 1568 29200 1968
rect 880 1288 29120 1568
rect 800 888 29200 1288
rect 880 608 29120 888
rect 800 208 29200 608
rect 800 35 29120 208
<< metal4 >>
rect 4418 2128 4738 27792
rect 7892 2128 8212 27792
rect 11366 2128 11686 27792
rect 14840 2128 15160 27792
rect 18314 2128 18634 27792
rect 21788 2128 22108 27792
rect 25262 2128 25582 27792
<< labels >>
rlabel metal2 s 7102 29200 7158 30000 6 b0_drv[0]
port 1 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 b0_drv[10]
port 2 nsew signal output
rlabel metal2 s 29642 29200 29698 30000 6 b0_drv[11]
port 3 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 b0_drv[12]
port 4 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 b0_drv[13]
port 5 nsew signal output
rlabel metal3 s 29200 9528 30000 9648 6 b0_drv[14]
port 6 nsew signal output
rlabel metal3 s 29200 25168 30000 25288 6 b0_drv[15]
port 7 nsew signal output
rlabel metal3 s 29200 17008 30000 17128 6 b0_drv[16]
port 8 nsew signal output
rlabel metal2 s 19338 29200 19394 30000 6 b0_drv[17]
port 9 nsew signal output
rlabel metal3 s 29200 4088 30000 4208 6 b0_drv[18]
port 10 nsew signal output
rlabel metal3 s 29200 19048 30000 19168 6 b0_drv[19]
port 11 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 b0_drv[1]
port 12 nsew signal output
rlabel metal2 s 23846 29200 23902 30000 6 b0_drv[20]
port 13 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 b0_drv[21]
port 14 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 b0_drv[22]
port 15 nsew signal output
rlabel metal2 s 28354 29200 28410 30000 6 b0_drv[23]
port 16 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 b0_drv[24]
port 17 nsew signal output
rlabel metal2 s 5814 29200 5870 30000 6 b0_drv[25]
port 18 nsew signal output
rlabel metal2 s 662 29200 718 30000 6 b0_drv[26]
port 19 nsew signal output
rlabel metal2 s 13542 29200 13598 30000 6 b0_drv[27]
port 20 nsew signal output
rlabel metal3 s 29200 10888 30000 11008 6 b0_drv[28]
port 21 nsew signal output
rlabel metal3 s 29200 2728 30000 2848 6 b0_drv[29]
port 22 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 b0_drv[2]
port 23 nsew signal output
rlabel metal3 s 29200 27208 30000 27328 6 b0_drv[30]
port 24 nsew signal output
rlabel metal2 s 16118 29200 16174 30000 6 b0_drv[31]
port 25 nsew signal output
rlabel metal2 s 11610 29200 11666 30000 6 b0_drv[32]
port 26 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 b0_drv[33]
port 27 nsew signal output
rlabel metal2 s 18050 29200 18106 30000 6 b0_drv[34]
port 28 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 b0_drv[35]
port 29 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 b0_drv[36]
port 30 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 b0_drv[37]
port 31 nsew signal output
rlabel metal3 s 29200 23808 30000 23928 6 b0_drv[38]
port 32 nsew signal output
rlabel metal2 s 25778 29200 25834 30000 6 b0_drv[39]
port 33 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 b0_drv[3]
port 34 nsew signal output
rlabel metal2 s 16762 29200 16818 30000 6 b0_drv[40]
port 35 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 b0_drv[41]
port 36 nsew signal output
rlabel metal3 s 29200 6808 30000 6928 6 b0_drv[42]
port 37 nsew signal output
rlabel metal2 s 7746 29200 7802 30000 6 b0_drv[43]
port 38 nsew signal output
rlabel metal3 s 29200 1368 30000 1488 6 b0_drv[44]
port 39 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 b0_drv[45]
port 40 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 b0_drv[46]
port 41 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 b0_drv[47]
port 42 nsew signal output
rlabel metal2 s 27066 29200 27122 30000 6 b0_drv[48]
port 43 nsew signal output
rlabel metal2 s 14186 29200 14242 30000 6 b0_drv[49]
port 44 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 b0_drv[4]
port 45 nsew signal output
rlabel metal3 s 29200 8 30000 128 6 b0_drv[50]
port 46 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 b0_drv[51]
port 47 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 b0_drv[52]
port 48 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 b0_drv[53]
port 49 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 b0_drv[54]
port 50 nsew signal output
rlabel metal2 s 12254 29200 12310 30000 6 b0_drv[55]
port 51 nsew signal output
rlabel metal2 s 17406 29200 17462 30000 6 b0_drv[56]
port 52 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 b0_drv[57]
port 53 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 b0_drv[58]
port 54 nsew signal output
rlabel metal3 s 29200 24488 30000 24608 6 b0_drv[59]
port 55 nsew signal output
rlabel metal2 s 2594 29200 2650 30000 6 b0_drv[5]
port 56 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 b0_drv[60]
port 57 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 b0_drv[61]
port 58 nsew signal output
rlabel metal3 s 0 688 800 808 6 b0_drv[62]
port 59 nsew signal output
rlabel metal3 s 29200 15648 30000 15768 6 b0_drv[63]
port 60 nsew signal output
rlabel metal2 s 12898 29200 12954 30000 6 b0_drv[64]
port 61 nsew signal output
rlabel metal3 s 29200 21768 30000 21888 6 b0_drv[65]
port 62 nsew signal output
rlabel metal2 s 26422 29200 26478 30000 6 b0_drv[66]
port 63 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 b0_drv[67]
port 64 nsew signal output
rlabel metal2 s 24490 29200 24546 30000 6 b0_drv[68]
port 65 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 b0_drv[69]
port 66 nsew signal output
rlabel metal2 s 9678 29200 9734 30000 6 b0_drv[6]
port 67 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 b0_drv[70]
port 68 nsew signal output
rlabel metal3 s 29200 11568 30000 11688 6 b0_drv[71]
port 69 nsew signal output
rlabel metal3 s 29200 2048 30000 2168 6 b0_drv[72]
port 70 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 b0_drv[73]
port 71 nsew signal output
rlabel metal3 s 29200 27888 30000 28008 6 b0_drv[74]
port 72 nsew signal output
rlabel metal3 s 29200 21088 30000 21208 6 b0_drv[75]
port 73 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 b0_drv[76]
port 74 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 b0_drv[77]
port 75 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 b0_drv[78]
port 76 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 b0_drv[79]
port 77 nsew signal output
rlabel metal3 s 29200 12928 30000 13048 6 b0_drv[7]
port 78 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 b0_drv[80]
port 79 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 b0_drv[81]
port 80 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 b0_drv[82]
port 81 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 b0_drv[8]
port 82 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 b0_drv[9]
port 83 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 cw_clk_i
port 84 nsew signal input
rlabel metal2 s 23202 29200 23258 30000 6 cw_clk_o
port 85 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 cw_dir
port 86 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 cw_dir_b_o
port 87 nsew signal input
rlabel metal3 s 29200 13608 30000 13728 6 cw_dir_b_oo
port 88 nsew signal output
rlabel metal3 s 29200 7488 30000 7608 6 cw_dir_o
port 89 nsew signal output
rlabel metal2 s 27710 29200 27766 30000 6 cw_req_i
port 90 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 cw_req_o
port 91 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 cw_rst_i
port 92 nsew signal input
rlabel metal3 s 29200 25848 30000 25968 6 cw_rst_o
port 93 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 io_oeb_15_0[0]
port 94 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_oeb_15_0[10]
port 95 nsew signal output
rlabel metal2 s 5170 29200 5226 30000 6 io_oeb_15_0[11]
port 96 nsew signal output
rlabel metal2 s 6458 29200 6514 30000 6 io_oeb_15_0[12]
port 97 nsew signal output
rlabel metal2 s 1306 29200 1362 30000 6 io_oeb_15_0[13]
port 98 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 io_oeb_15_0[14]
port 99 nsew signal output
rlabel metal3 s 29200 14968 30000 15088 6 io_oeb_15_0[15]
port 100 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 io_oeb_15_0[1]
port 101 nsew signal output
rlabel metal2 s 10966 29200 11022 30000 6 io_oeb_15_0[2]
port 102 nsew signal output
rlabel metal3 s 29200 16328 30000 16448 6 io_oeb_15_0[3]
port 103 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 io_oeb_15_0[4]
port 104 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 io_oeb_15_0[5]
port 105 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 io_oeb_15_0[6]
port 106 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 io_oeb_15_0[7]
port 107 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 io_oeb_15_0[8]
port 108 nsew signal output
rlabel metal3 s 29200 28568 30000 28688 6 io_oeb_15_0[9]
port 109 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 io_oeb_18_16[0]
port 110 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_oeb_18_16[1]
port 111 nsew signal output
rlabel metal2 s 19982 29200 20038 30000 6 io_oeb_18_16[2]
port 112 nsew signal output
rlabel metal2 s 18694 29200 18750 30000 6 io_oeb_20_19[0]
port 113 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_oeb_20_19[1]
port 114 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 io_oeb_21
port 115 nsew signal output
rlabel metal3 s 29200 3408 30000 3528 6 io_oeb_22
port 116 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 io_out[0]
port 117 nsew signal output
rlabel metal3 s 29200 23128 30000 23248 6 io_out[10]
port 118 nsew signal output
rlabel metal2 s 8390 29200 8446 30000 6 io_out[11]
port 119 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 io_out[12]
port 120 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 io_out[13]
port 121 nsew signal output
rlabel metal3 s 29200 6128 30000 6248 6 io_out[14]
port 122 nsew signal output
rlabel metal3 s 29200 17688 30000 17808 6 io_out[1]
port 123 nsew signal output
rlabel metal2 s 9034 29200 9090 30000 6 io_out[2]
port 124 nsew signal output
rlabel metal3 s 29200 12248 30000 12368 6 io_out[3]
port 125 nsew signal output
rlabel metal2 s 1950 29200 2006 30000 6 io_out[4]
port 126 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 io_out[5]
port 127 nsew signal output
rlabel metal3 s 29200 22448 30000 22568 6 io_out[6]
port 128 nsew signal output
rlabel metal2 s 22558 29200 22614 30000 6 io_out[7]
port 129 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 io_out[8]
port 130 nsew signal output
rlabel metal3 s 29200 8168 30000 8288 6 io_out[9]
port 131 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 io_out_20_19[0]
port 132 nsew signal output
rlabel metal3 s 29200 688 30000 808 6 io_out_20_19[1]
port 133 nsew signal output
rlabel metal2 s 3238 29200 3294 30000 6 io_out_22
port 134 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 la_data_out_16_17[0]
port 135 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 la_data_out_16_17[1]
port 136 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 la_data_out_21
port 137 nsew signal output
rlabel metal3 s 29200 5448 30000 5568 6 la_data_out_37_36[0]
port 138 nsew signal output
rlabel metal3 s 29200 26528 30000 26648 6 la_data_out_37_36[1]
port 139 nsew signal output
rlabel metal3 s 29200 18368 30000 18488 6 la_data_out_77_62[0]
port 140 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 la_data_out_77_62[10]
port 141 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 la_data_out_77_62[11]
port 142 nsew signal output
rlabel metal3 s 29200 10208 30000 10328 6 la_data_out_77_62[12]
port 143 nsew signal output
rlabel metal2 s 662 0 718 800 6 la_data_out_77_62[13]
port 144 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 la_data_out_77_62[14]
port 145 nsew signal output
rlabel metal3 s 29200 29248 30000 29368 6 la_data_out_77_62[15]
port 146 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 la_data_out_77_62[1]
port 147 nsew signal output
rlabel metal2 s 28998 29200 29054 30000 6 la_data_out_77_62[2]
port 148 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out_77_62[3]
port 149 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 la_data_out_77_62[4]
port 150 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 la_data_out_77_62[5]
port 151 nsew signal output
rlabel metal2 s 18 0 74 800 6 la_data_out_77_62[6]
port 152 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 la_data_out_77_62[7]
port 153 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 la_data_out_77_62[8]
port 154 nsew signal output
rlabel metal2 s 3882 29200 3938 30000 6 la_data_out_77_62[9]
port 155 nsew signal output
rlabel metal2 s 15474 29200 15530 30000 6 la_data_out_97_95[0]
port 156 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 la_data_out_97_95[1]
port 157 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 la_data_out_97_95[2]
port 158 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 la_datb_i[0]
port 159 nsew signal input
rlabel metal2 s 20626 29200 20682 30000 6 la_datb_i[1]
port 160 nsew signal input
rlabel metal2 s 14830 29200 14886 30000 6 la_datb_i[2]
port 161 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 la_datb_o[0]
port 162 nsew signal output
rlabel metal2 s 25134 29200 25190 30000 6 la_datb_o[1]
port 163 nsew signal output
rlabel metal3 s 29200 4768 30000 4888 6 la_datb_o[2]
port 164 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 oeb_out[0]
port 165 nsew signal output
rlabel metal3 s 29200 20408 30000 20528 6 oeb_out[10]
port 166 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 oeb_out[11]
port 167 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 oeb_out[12]
port 168 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 oeb_out[13]
port 169 nsew signal output
rlabel metal3 s 29200 19728 30000 19848 6 oeb_out[14]
port 170 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 oeb_out[1]
port 171 nsew signal output
rlabel metal2 s 21914 29200 21970 30000 6 oeb_out[2]
port 172 nsew signal output
rlabel metal2 s 21270 29200 21326 30000 6 oeb_out[3]
port 173 nsew signal output
rlabel metal2 s 18 29200 74 30000 6 oeb_out[4]
port 174 nsew signal output
rlabel metal2 s 4526 29200 4582 30000 6 oeb_out[5]
port 175 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 oeb_out[6]
port 176 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 oeb_out[7]
port 177 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 oeb_out[8]
port 178 nsew signal output
rlabel metal3 s 29200 14288 30000 14408 6 oeb_out[9]
port 179 nsew signal output
rlabel metal4 s 4418 2128 4738 27792 6 vccd1
port 180 nsew power bidirectional
rlabel metal4 s 11366 2128 11686 27792 6 vccd1
port 180 nsew power bidirectional
rlabel metal4 s 18314 2128 18634 27792 6 vccd1
port 180 nsew power bidirectional
rlabel metal4 s 25262 2128 25582 27792 6 vccd1
port 180 nsew power bidirectional
rlabel metal4 s 7892 2128 8212 27792 6 vssd1
port 181 nsew ground bidirectional
rlabel metal4 s 14840 2128 15160 27792 6 vssd1
port 181 nsew ground bidirectional
rlabel metal4 s 21788 2128 22108 27792 6 vssd1
port 181 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 602484
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/uprj_w_const/runs/22_09_13_08_43/results/signoff/uprj_w_const.magic.gds
string GDS_START 50412
<< end >>

