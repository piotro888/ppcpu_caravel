VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO interconnect_inner
  CLASS BLOCK ;
  FOREIGN interconnect_inner ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 800.000 ;
  PIN c0_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END c0_clk
  PIN c0_dbg_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END c0_dbg_pc[0]
  PIN c0_dbg_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END c0_dbg_pc[10]
  PIN c0_dbg_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END c0_dbg_pc[11]
  PIN c0_dbg_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END c0_dbg_pc[12]
  PIN c0_dbg_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END c0_dbg_pc[13]
  PIN c0_dbg_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END c0_dbg_pc[14]
  PIN c0_dbg_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END c0_dbg_pc[15]
  PIN c0_dbg_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END c0_dbg_pc[1]
  PIN c0_dbg_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END c0_dbg_pc[2]
  PIN c0_dbg_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END c0_dbg_pc[3]
  PIN c0_dbg_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END c0_dbg_pc[4]
  PIN c0_dbg_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END c0_dbg_pc[5]
  PIN c0_dbg_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END c0_dbg_pc[6]
  PIN c0_dbg_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END c0_dbg_pc[7]
  PIN c0_dbg_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END c0_dbg_pc[8]
  PIN c0_dbg_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END c0_dbg_pc[9]
  PIN c0_dbg_r0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END c0_dbg_r0[0]
  PIN c0_dbg_r0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END c0_dbg_r0[10]
  PIN c0_dbg_r0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END c0_dbg_r0[11]
  PIN c0_dbg_r0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END c0_dbg_r0[12]
  PIN c0_dbg_r0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END c0_dbg_r0[13]
  PIN c0_dbg_r0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END c0_dbg_r0[14]
  PIN c0_dbg_r0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END c0_dbg_r0[15]
  PIN c0_dbg_r0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END c0_dbg_r0[1]
  PIN c0_dbg_r0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END c0_dbg_r0[2]
  PIN c0_dbg_r0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END c0_dbg_r0[3]
  PIN c0_dbg_r0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END c0_dbg_r0[4]
  PIN c0_dbg_r0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END c0_dbg_r0[5]
  PIN c0_dbg_r0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END c0_dbg_r0[6]
  PIN c0_dbg_r0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END c0_dbg_r0[7]
  PIN c0_dbg_r0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END c0_dbg_r0[8]
  PIN c0_dbg_r0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END c0_dbg_r0[9]
  PIN c0_disable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END c0_disable
  PIN c0_i_core_int_sreg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END c0_i_core_int_sreg[0]
  PIN c0_i_core_int_sreg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END c0_i_core_int_sreg[10]
  PIN c0_i_core_int_sreg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END c0_i_core_int_sreg[11]
  PIN c0_i_core_int_sreg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END c0_i_core_int_sreg[12]
  PIN c0_i_core_int_sreg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END c0_i_core_int_sreg[13]
  PIN c0_i_core_int_sreg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END c0_i_core_int_sreg[14]
  PIN c0_i_core_int_sreg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END c0_i_core_int_sreg[15]
  PIN c0_i_core_int_sreg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END c0_i_core_int_sreg[1]
  PIN c0_i_core_int_sreg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END c0_i_core_int_sreg[2]
  PIN c0_i_core_int_sreg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END c0_i_core_int_sreg[3]
  PIN c0_i_core_int_sreg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END c0_i_core_int_sreg[4]
  PIN c0_i_core_int_sreg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END c0_i_core_int_sreg[5]
  PIN c0_i_core_int_sreg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END c0_i_core_int_sreg[6]
  PIN c0_i_core_int_sreg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END c0_i_core_int_sreg[7]
  PIN c0_i_core_int_sreg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END c0_i_core_int_sreg[8]
  PIN c0_i_core_int_sreg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END c0_i_core_int_sreg[9]
  PIN c0_i_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END c0_i_irq
  PIN c0_i_mc_core_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END c0_i_mc_core_int
  PIN c0_i_mem_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END c0_i_mem_ack
  PIN c0_i_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END c0_i_mem_data[0]
  PIN c0_i_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END c0_i_mem_data[10]
  PIN c0_i_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END c0_i_mem_data[11]
  PIN c0_i_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END c0_i_mem_data[12]
  PIN c0_i_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END c0_i_mem_data[13]
  PIN c0_i_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END c0_i_mem_data[14]
  PIN c0_i_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END c0_i_mem_data[15]
  PIN c0_i_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END c0_i_mem_data[1]
  PIN c0_i_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END c0_i_mem_data[2]
  PIN c0_i_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END c0_i_mem_data[3]
  PIN c0_i_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END c0_i_mem_data[4]
  PIN c0_i_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END c0_i_mem_data[5]
  PIN c0_i_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END c0_i_mem_data[6]
  PIN c0_i_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END c0_i_mem_data[7]
  PIN c0_i_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END c0_i_mem_data[8]
  PIN c0_i_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END c0_i_mem_data[9]
  PIN c0_i_mem_exception
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END c0_i_mem_exception
  PIN c0_i_req_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END c0_i_req_data[0]
  PIN c0_i_req_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END c0_i_req_data[10]
  PIN c0_i_req_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END c0_i_req_data[11]
  PIN c0_i_req_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END c0_i_req_data[12]
  PIN c0_i_req_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END c0_i_req_data[13]
  PIN c0_i_req_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END c0_i_req_data[14]
  PIN c0_i_req_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END c0_i_req_data[15]
  PIN c0_i_req_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END c0_i_req_data[16]
  PIN c0_i_req_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END c0_i_req_data[17]
  PIN c0_i_req_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END c0_i_req_data[18]
  PIN c0_i_req_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END c0_i_req_data[19]
  PIN c0_i_req_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END c0_i_req_data[1]
  PIN c0_i_req_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END c0_i_req_data[20]
  PIN c0_i_req_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END c0_i_req_data[21]
  PIN c0_i_req_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END c0_i_req_data[22]
  PIN c0_i_req_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END c0_i_req_data[23]
  PIN c0_i_req_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END c0_i_req_data[24]
  PIN c0_i_req_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END c0_i_req_data[25]
  PIN c0_i_req_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END c0_i_req_data[26]
  PIN c0_i_req_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END c0_i_req_data[27]
  PIN c0_i_req_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END c0_i_req_data[28]
  PIN c0_i_req_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END c0_i_req_data[29]
  PIN c0_i_req_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END c0_i_req_data[2]
  PIN c0_i_req_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END c0_i_req_data[30]
  PIN c0_i_req_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END c0_i_req_data[31]
  PIN c0_i_req_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END c0_i_req_data[3]
  PIN c0_i_req_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END c0_i_req_data[4]
  PIN c0_i_req_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END c0_i_req_data[5]
  PIN c0_i_req_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END c0_i_req_data[6]
  PIN c0_i_req_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END c0_i_req_data[7]
  PIN c0_i_req_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END c0_i_req_data[8]
  PIN c0_i_req_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END c0_i_req_data[9]
  PIN c0_i_req_data_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END c0_i_req_data_valid
  PIN c0_o_c_data_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END c0_o_c_data_page
  PIN c0_o_c_instr_long
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END c0_o_c_instr_long
  PIN c0_o_c_instr_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END c0_o_c_instr_page
  PIN c0_o_icache_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END c0_o_icache_flush
  PIN c0_o_instr_long_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END c0_o_instr_long_addr[0]
  PIN c0_o_instr_long_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END c0_o_instr_long_addr[1]
  PIN c0_o_instr_long_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END c0_o_instr_long_addr[2]
  PIN c0_o_instr_long_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END c0_o_instr_long_addr[3]
  PIN c0_o_instr_long_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END c0_o_instr_long_addr[4]
  PIN c0_o_instr_long_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END c0_o_instr_long_addr[5]
  PIN c0_o_instr_long_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END c0_o_instr_long_addr[6]
  PIN c0_o_instr_long_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END c0_o_instr_long_addr[7]
  PIN c0_o_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END c0_o_mem_addr[0]
  PIN c0_o_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END c0_o_mem_addr[10]
  PIN c0_o_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END c0_o_mem_addr[11]
  PIN c0_o_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END c0_o_mem_addr[12]
  PIN c0_o_mem_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END c0_o_mem_addr[13]
  PIN c0_o_mem_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END c0_o_mem_addr[14]
  PIN c0_o_mem_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END c0_o_mem_addr[15]
  PIN c0_o_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END c0_o_mem_addr[1]
  PIN c0_o_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END c0_o_mem_addr[2]
  PIN c0_o_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END c0_o_mem_addr[3]
  PIN c0_o_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END c0_o_mem_addr[4]
  PIN c0_o_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END c0_o_mem_addr[5]
  PIN c0_o_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END c0_o_mem_addr[6]
  PIN c0_o_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END c0_o_mem_addr[7]
  PIN c0_o_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END c0_o_mem_addr[8]
  PIN c0_o_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END c0_o_mem_addr[9]
  PIN c0_o_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END c0_o_mem_data[0]
  PIN c0_o_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END c0_o_mem_data[10]
  PIN c0_o_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END c0_o_mem_data[11]
  PIN c0_o_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END c0_o_mem_data[12]
  PIN c0_o_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END c0_o_mem_data[13]
  PIN c0_o_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END c0_o_mem_data[14]
  PIN c0_o_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END c0_o_mem_data[15]
  PIN c0_o_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END c0_o_mem_data[1]
  PIN c0_o_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END c0_o_mem_data[2]
  PIN c0_o_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END c0_o_mem_data[3]
  PIN c0_o_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END c0_o_mem_data[4]
  PIN c0_o_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END c0_o_mem_data[5]
  PIN c0_o_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END c0_o_mem_data[6]
  PIN c0_o_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END c0_o_mem_data[7]
  PIN c0_o_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END c0_o_mem_data[8]
  PIN c0_o_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END c0_o_mem_data[9]
  PIN c0_o_mem_high_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END c0_o_mem_high_addr[0]
  PIN c0_o_mem_high_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END c0_o_mem_high_addr[1]
  PIN c0_o_mem_high_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END c0_o_mem_high_addr[2]
  PIN c0_o_mem_high_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END c0_o_mem_high_addr[3]
  PIN c0_o_mem_high_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END c0_o_mem_high_addr[4]
  PIN c0_o_mem_high_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END c0_o_mem_high_addr[5]
  PIN c0_o_mem_high_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END c0_o_mem_high_addr[6]
  PIN c0_o_mem_high_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END c0_o_mem_high_addr[7]
  PIN c0_o_mem_long_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END c0_o_mem_long_mode
  PIN c0_o_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END c0_o_mem_req
  PIN c0_o_mem_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END c0_o_mem_sel[0]
  PIN c0_o_mem_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END c0_o_mem_sel[1]
  PIN c0_o_mem_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END c0_o_mem_we
  PIN c0_o_req_active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END c0_o_req_active
  PIN c0_o_req_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END c0_o_req_addr[0]
  PIN c0_o_req_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END c0_o_req_addr[10]
  PIN c0_o_req_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END c0_o_req_addr[11]
  PIN c0_o_req_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END c0_o_req_addr[12]
  PIN c0_o_req_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END c0_o_req_addr[13]
  PIN c0_o_req_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END c0_o_req_addr[14]
  PIN c0_o_req_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END c0_o_req_addr[15]
  PIN c0_o_req_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END c0_o_req_addr[1]
  PIN c0_o_req_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END c0_o_req_addr[2]
  PIN c0_o_req_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END c0_o_req_addr[3]
  PIN c0_o_req_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END c0_o_req_addr[4]
  PIN c0_o_req_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END c0_o_req_addr[5]
  PIN c0_o_req_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END c0_o_req_addr[6]
  PIN c0_o_req_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END c0_o_req_addr[7]
  PIN c0_o_req_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END c0_o_req_addr[8]
  PIN c0_o_req_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END c0_o_req_addr[9]
  PIN c0_o_req_ppl_submit
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END c0_o_req_ppl_submit
  PIN c0_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END c0_rst
  PIN c0_sr_bus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END c0_sr_bus_addr[0]
  PIN c0_sr_bus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END c0_sr_bus_addr[10]
  PIN c0_sr_bus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END c0_sr_bus_addr[11]
  PIN c0_sr_bus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END c0_sr_bus_addr[12]
  PIN c0_sr_bus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END c0_sr_bus_addr[13]
  PIN c0_sr_bus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END c0_sr_bus_addr[14]
  PIN c0_sr_bus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END c0_sr_bus_addr[15]
  PIN c0_sr_bus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END c0_sr_bus_addr[1]
  PIN c0_sr_bus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END c0_sr_bus_addr[2]
  PIN c0_sr_bus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END c0_sr_bus_addr[3]
  PIN c0_sr_bus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END c0_sr_bus_addr[4]
  PIN c0_sr_bus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END c0_sr_bus_addr[5]
  PIN c0_sr_bus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END c0_sr_bus_addr[6]
  PIN c0_sr_bus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END c0_sr_bus_addr[7]
  PIN c0_sr_bus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END c0_sr_bus_addr[8]
  PIN c0_sr_bus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END c0_sr_bus_addr[9]
  PIN c0_sr_bus_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END c0_sr_bus_data_o[0]
  PIN c0_sr_bus_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END c0_sr_bus_data_o[10]
  PIN c0_sr_bus_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END c0_sr_bus_data_o[11]
  PIN c0_sr_bus_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END c0_sr_bus_data_o[12]
  PIN c0_sr_bus_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END c0_sr_bus_data_o[13]
  PIN c0_sr_bus_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END c0_sr_bus_data_o[14]
  PIN c0_sr_bus_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END c0_sr_bus_data_o[15]
  PIN c0_sr_bus_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END c0_sr_bus_data_o[1]
  PIN c0_sr_bus_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END c0_sr_bus_data_o[2]
  PIN c0_sr_bus_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END c0_sr_bus_data_o[3]
  PIN c0_sr_bus_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END c0_sr_bus_data_o[4]
  PIN c0_sr_bus_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END c0_sr_bus_data_o[5]
  PIN c0_sr_bus_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END c0_sr_bus_data_o[6]
  PIN c0_sr_bus_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END c0_sr_bus_data_o[7]
  PIN c0_sr_bus_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END c0_sr_bus_data_o[8]
  PIN c0_sr_bus_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END c0_sr_bus_data_o[9]
  PIN c0_sr_bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END c0_sr_bus_we
  PIN c1_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END c1_clk
  PIN c1_dbg_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END c1_dbg_pc[0]
  PIN c1_dbg_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END c1_dbg_pc[10]
  PIN c1_dbg_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END c1_dbg_pc[11]
  PIN c1_dbg_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END c1_dbg_pc[12]
  PIN c1_dbg_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END c1_dbg_pc[13]
  PIN c1_dbg_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END c1_dbg_pc[14]
  PIN c1_dbg_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END c1_dbg_pc[15]
  PIN c1_dbg_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END c1_dbg_pc[1]
  PIN c1_dbg_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END c1_dbg_pc[2]
  PIN c1_dbg_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END c1_dbg_pc[3]
  PIN c1_dbg_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END c1_dbg_pc[4]
  PIN c1_dbg_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END c1_dbg_pc[5]
  PIN c1_dbg_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END c1_dbg_pc[6]
  PIN c1_dbg_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END c1_dbg_pc[7]
  PIN c1_dbg_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END c1_dbg_pc[8]
  PIN c1_dbg_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END c1_dbg_pc[9]
  PIN c1_dbg_r0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END c1_dbg_r0[0]
  PIN c1_dbg_r0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END c1_dbg_r0[10]
  PIN c1_dbg_r0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END c1_dbg_r0[11]
  PIN c1_dbg_r0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END c1_dbg_r0[12]
  PIN c1_dbg_r0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END c1_dbg_r0[13]
  PIN c1_dbg_r0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END c1_dbg_r0[14]
  PIN c1_dbg_r0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END c1_dbg_r0[15]
  PIN c1_dbg_r0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END c1_dbg_r0[1]
  PIN c1_dbg_r0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END c1_dbg_r0[2]
  PIN c1_dbg_r0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END c1_dbg_r0[3]
  PIN c1_dbg_r0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END c1_dbg_r0[4]
  PIN c1_dbg_r0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END c1_dbg_r0[5]
  PIN c1_dbg_r0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END c1_dbg_r0[6]
  PIN c1_dbg_r0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END c1_dbg_r0[7]
  PIN c1_dbg_r0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END c1_dbg_r0[8]
  PIN c1_dbg_r0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END c1_dbg_r0[9]
  PIN c1_disable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END c1_disable
  PIN c1_i_core_int_sreg[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END c1_i_core_int_sreg[0]
  PIN c1_i_core_int_sreg[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END c1_i_core_int_sreg[10]
  PIN c1_i_core_int_sreg[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END c1_i_core_int_sreg[11]
  PIN c1_i_core_int_sreg[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END c1_i_core_int_sreg[12]
  PIN c1_i_core_int_sreg[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END c1_i_core_int_sreg[13]
  PIN c1_i_core_int_sreg[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END c1_i_core_int_sreg[14]
  PIN c1_i_core_int_sreg[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END c1_i_core_int_sreg[15]
  PIN c1_i_core_int_sreg[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END c1_i_core_int_sreg[1]
  PIN c1_i_core_int_sreg[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END c1_i_core_int_sreg[2]
  PIN c1_i_core_int_sreg[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END c1_i_core_int_sreg[3]
  PIN c1_i_core_int_sreg[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END c1_i_core_int_sreg[4]
  PIN c1_i_core_int_sreg[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END c1_i_core_int_sreg[5]
  PIN c1_i_core_int_sreg[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END c1_i_core_int_sreg[6]
  PIN c1_i_core_int_sreg[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END c1_i_core_int_sreg[7]
  PIN c1_i_core_int_sreg[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END c1_i_core_int_sreg[8]
  PIN c1_i_core_int_sreg[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END c1_i_core_int_sreg[9]
  PIN c1_i_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END c1_i_irq
  PIN c1_i_mc_core_int
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END c1_i_mc_core_int
  PIN c1_i_mem_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END c1_i_mem_ack
  PIN c1_i_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END c1_i_mem_data[0]
  PIN c1_i_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END c1_i_mem_data[10]
  PIN c1_i_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END c1_i_mem_data[11]
  PIN c1_i_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END c1_i_mem_data[12]
  PIN c1_i_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END c1_i_mem_data[13]
  PIN c1_i_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END c1_i_mem_data[14]
  PIN c1_i_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END c1_i_mem_data[15]
  PIN c1_i_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END c1_i_mem_data[1]
  PIN c1_i_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END c1_i_mem_data[2]
  PIN c1_i_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END c1_i_mem_data[3]
  PIN c1_i_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END c1_i_mem_data[4]
  PIN c1_i_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END c1_i_mem_data[5]
  PIN c1_i_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END c1_i_mem_data[6]
  PIN c1_i_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END c1_i_mem_data[7]
  PIN c1_i_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END c1_i_mem_data[8]
  PIN c1_i_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END c1_i_mem_data[9]
  PIN c1_i_mem_exception
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END c1_i_mem_exception
  PIN c1_i_req_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END c1_i_req_data[0]
  PIN c1_i_req_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END c1_i_req_data[10]
  PIN c1_i_req_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.880 4.000 604.480 ;
    END
  END c1_i_req_data[11]
  PIN c1_i_req_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END c1_i_req_data[12]
  PIN c1_i_req_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END c1_i_req_data[13]
  PIN c1_i_req_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END c1_i_req_data[14]
  PIN c1_i_req_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END c1_i_req_data[15]
  PIN c1_i_req_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END c1_i_req_data[16]
  PIN c1_i_req_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END c1_i_req_data[17]
  PIN c1_i_req_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END c1_i_req_data[18]
  PIN c1_i_req_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END c1_i_req_data[19]
  PIN c1_i_req_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END c1_i_req_data[1]
  PIN c1_i_req_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END c1_i_req_data[20]
  PIN c1_i_req_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END c1_i_req_data[21]
  PIN c1_i_req_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END c1_i_req_data[22]
  PIN c1_i_req_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END c1_i_req_data[23]
  PIN c1_i_req_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END c1_i_req_data[24]
  PIN c1_i_req_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END c1_i_req_data[25]
  PIN c1_i_req_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END c1_i_req_data[26]
  PIN c1_i_req_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END c1_i_req_data[27]
  PIN c1_i_req_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END c1_i_req_data[28]
  PIN c1_i_req_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END c1_i_req_data[29]
  PIN c1_i_req_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END c1_i_req_data[2]
  PIN c1_i_req_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END c1_i_req_data[30]
  PIN c1_i_req_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END c1_i_req_data[31]
  PIN c1_i_req_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END c1_i_req_data[3]
  PIN c1_i_req_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END c1_i_req_data[4]
  PIN c1_i_req_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END c1_i_req_data[5]
  PIN c1_i_req_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END c1_i_req_data[6]
  PIN c1_i_req_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END c1_i_req_data[7]
  PIN c1_i_req_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END c1_i_req_data[8]
  PIN c1_i_req_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END c1_i_req_data[9]
  PIN c1_i_req_data_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END c1_i_req_data_valid
  PIN c1_o_c_data_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END c1_o_c_data_page
  PIN c1_o_c_instr_long
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END c1_o_c_instr_long
  PIN c1_o_c_instr_page
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END c1_o_c_instr_page
  PIN c1_o_icache_flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END c1_o_icache_flush
  PIN c1_o_instr_long_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END c1_o_instr_long_addr[0]
  PIN c1_o_instr_long_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END c1_o_instr_long_addr[1]
  PIN c1_o_instr_long_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END c1_o_instr_long_addr[2]
  PIN c1_o_instr_long_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END c1_o_instr_long_addr[3]
  PIN c1_o_instr_long_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END c1_o_instr_long_addr[4]
  PIN c1_o_instr_long_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END c1_o_instr_long_addr[5]
  PIN c1_o_instr_long_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END c1_o_instr_long_addr[6]
  PIN c1_o_instr_long_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END c1_o_instr_long_addr[7]
  PIN c1_o_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END c1_o_mem_addr[0]
  PIN c1_o_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END c1_o_mem_addr[10]
  PIN c1_o_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END c1_o_mem_addr[11]
  PIN c1_o_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END c1_o_mem_addr[12]
  PIN c1_o_mem_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END c1_o_mem_addr[13]
  PIN c1_o_mem_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END c1_o_mem_addr[14]
  PIN c1_o_mem_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END c1_o_mem_addr[15]
  PIN c1_o_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END c1_o_mem_addr[1]
  PIN c1_o_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END c1_o_mem_addr[2]
  PIN c1_o_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END c1_o_mem_addr[3]
  PIN c1_o_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END c1_o_mem_addr[4]
  PIN c1_o_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END c1_o_mem_addr[5]
  PIN c1_o_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END c1_o_mem_addr[6]
  PIN c1_o_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END c1_o_mem_addr[7]
  PIN c1_o_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END c1_o_mem_addr[8]
  PIN c1_o_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END c1_o_mem_addr[9]
  PIN c1_o_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END c1_o_mem_data[0]
  PIN c1_o_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END c1_o_mem_data[10]
  PIN c1_o_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END c1_o_mem_data[11]
  PIN c1_o_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END c1_o_mem_data[12]
  PIN c1_o_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END c1_o_mem_data[13]
  PIN c1_o_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END c1_o_mem_data[14]
  PIN c1_o_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END c1_o_mem_data[15]
  PIN c1_o_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END c1_o_mem_data[1]
  PIN c1_o_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END c1_o_mem_data[2]
  PIN c1_o_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END c1_o_mem_data[3]
  PIN c1_o_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END c1_o_mem_data[4]
  PIN c1_o_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END c1_o_mem_data[5]
  PIN c1_o_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END c1_o_mem_data[6]
  PIN c1_o_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END c1_o_mem_data[7]
  PIN c1_o_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END c1_o_mem_data[8]
  PIN c1_o_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END c1_o_mem_data[9]
  PIN c1_o_mem_high_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END c1_o_mem_high_addr[0]
  PIN c1_o_mem_high_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END c1_o_mem_high_addr[1]
  PIN c1_o_mem_high_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END c1_o_mem_high_addr[2]
  PIN c1_o_mem_high_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END c1_o_mem_high_addr[3]
  PIN c1_o_mem_high_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END c1_o_mem_high_addr[4]
  PIN c1_o_mem_high_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END c1_o_mem_high_addr[5]
  PIN c1_o_mem_high_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END c1_o_mem_high_addr[6]
  PIN c1_o_mem_high_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END c1_o_mem_high_addr[7]
  PIN c1_o_mem_long_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END c1_o_mem_long_mode
  PIN c1_o_mem_req
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END c1_o_mem_req
  PIN c1_o_mem_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END c1_o_mem_sel[0]
  PIN c1_o_mem_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END c1_o_mem_sel[1]
  PIN c1_o_mem_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END c1_o_mem_we
  PIN c1_o_req_active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END c1_o_req_active
  PIN c1_o_req_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END c1_o_req_addr[0]
  PIN c1_o_req_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END c1_o_req_addr[10]
  PIN c1_o_req_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END c1_o_req_addr[11]
  PIN c1_o_req_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END c1_o_req_addr[12]
  PIN c1_o_req_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END c1_o_req_addr[13]
  PIN c1_o_req_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END c1_o_req_addr[14]
  PIN c1_o_req_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END c1_o_req_addr[15]
  PIN c1_o_req_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END c1_o_req_addr[1]
  PIN c1_o_req_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END c1_o_req_addr[2]
  PIN c1_o_req_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END c1_o_req_addr[3]
  PIN c1_o_req_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END c1_o_req_addr[4]
  PIN c1_o_req_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END c1_o_req_addr[5]
  PIN c1_o_req_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END c1_o_req_addr[6]
  PIN c1_o_req_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END c1_o_req_addr[7]
  PIN c1_o_req_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END c1_o_req_addr[8]
  PIN c1_o_req_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END c1_o_req_addr[9]
  PIN c1_o_req_ppl_submit
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END c1_o_req_ppl_submit
  PIN c1_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END c1_rst
  PIN c1_sr_bus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END c1_sr_bus_addr[0]
  PIN c1_sr_bus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END c1_sr_bus_addr[10]
  PIN c1_sr_bus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END c1_sr_bus_addr[11]
  PIN c1_sr_bus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END c1_sr_bus_addr[12]
  PIN c1_sr_bus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END c1_sr_bus_addr[13]
  PIN c1_sr_bus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END c1_sr_bus_addr[14]
  PIN c1_sr_bus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END c1_sr_bus_addr[15]
  PIN c1_sr_bus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END c1_sr_bus_addr[1]
  PIN c1_sr_bus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END c1_sr_bus_addr[2]
  PIN c1_sr_bus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END c1_sr_bus_addr[3]
  PIN c1_sr_bus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END c1_sr_bus_addr[4]
  PIN c1_sr_bus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END c1_sr_bus_addr[5]
  PIN c1_sr_bus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END c1_sr_bus_addr[6]
  PIN c1_sr_bus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END c1_sr_bus_addr[7]
  PIN c1_sr_bus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END c1_sr_bus_addr[8]
  PIN c1_sr_bus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END c1_sr_bus_addr[9]
  PIN c1_sr_bus_data_o[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END c1_sr_bus_data_o[0]
  PIN c1_sr_bus_data_o[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END c1_sr_bus_data_o[10]
  PIN c1_sr_bus_data_o[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END c1_sr_bus_data_o[11]
  PIN c1_sr_bus_data_o[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END c1_sr_bus_data_o[12]
  PIN c1_sr_bus_data_o[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END c1_sr_bus_data_o[13]
  PIN c1_sr_bus_data_o[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END c1_sr_bus_data_o[14]
  PIN c1_sr_bus_data_o[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END c1_sr_bus_data_o[15]
  PIN c1_sr_bus_data_o[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END c1_sr_bus_data_o[1]
  PIN c1_sr_bus_data_o[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END c1_sr_bus_data_o[2]
  PIN c1_sr_bus_data_o[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END c1_sr_bus_data_o[3]
  PIN c1_sr_bus_data_o[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END c1_sr_bus_data_o[4]
  PIN c1_sr_bus_data_o[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END c1_sr_bus_data_o[5]
  PIN c1_sr_bus_data_o[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END c1_sr_bus_data_o[6]
  PIN c1_sr_bus_data_o[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END c1_sr_bus_data_o[7]
  PIN c1_sr_bus_data_o[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END c1_sr_bus_data_o[8]
  PIN c1_sr_bus_data_o[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END c1_sr_bus_data_o[9]
  PIN c1_sr_bus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END c1_sr_bus_we
  PIN core_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 796.000 7.270 800.000 ;
    END
  END core_clock
  PIN core_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 796.000 11.410 800.000 ;
    END
  END core_reset
  PIN dcache_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END dcache_clk
  PIN dcache_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END dcache_mem_ack
  PIN dcache_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END dcache_mem_addr[0]
  PIN dcache_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END dcache_mem_addr[10]
  PIN dcache_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END dcache_mem_addr[11]
  PIN dcache_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END dcache_mem_addr[12]
  PIN dcache_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END dcache_mem_addr[13]
  PIN dcache_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END dcache_mem_addr[14]
  PIN dcache_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END dcache_mem_addr[15]
  PIN dcache_mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END dcache_mem_addr[16]
  PIN dcache_mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END dcache_mem_addr[17]
  PIN dcache_mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END dcache_mem_addr[18]
  PIN dcache_mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END dcache_mem_addr[19]
  PIN dcache_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END dcache_mem_addr[1]
  PIN dcache_mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END dcache_mem_addr[20]
  PIN dcache_mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END dcache_mem_addr[21]
  PIN dcache_mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END dcache_mem_addr[22]
  PIN dcache_mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END dcache_mem_addr[23]
  PIN dcache_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END dcache_mem_addr[2]
  PIN dcache_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END dcache_mem_addr[3]
  PIN dcache_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END dcache_mem_addr[4]
  PIN dcache_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END dcache_mem_addr[5]
  PIN dcache_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END dcache_mem_addr[6]
  PIN dcache_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END dcache_mem_addr[7]
  PIN dcache_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END dcache_mem_addr[8]
  PIN dcache_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END dcache_mem_addr[9]
  PIN dcache_mem_cache_enable
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END dcache_mem_cache_enable
  PIN dcache_mem_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END dcache_mem_exception
  PIN dcache_mem_i_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END dcache_mem_i_data[0]
  PIN dcache_mem_i_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END dcache_mem_i_data[10]
  PIN dcache_mem_i_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END dcache_mem_i_data[11]
  PIN dcache_mem_i_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END dcache_mem_i_data[12]
  PIN dcache_mem_i_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END dcache_mem_i_data[13]
  PIN dcache_mem_i_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END dcache_mem_i_data[14]
  PIN dcache_mem_i_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END dcache_mem_i_data[15]
  PIN dcache_mem_i_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END dcache_mem_i_data[1]
  PIN dcache_mem_i_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END dcache_mem_i_data[2]
  PIN dcache_mem_i_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END dcache_mem_i_data[3]
  PIN dcache_mem_i_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END dcache_mem_i_data[4]
  PIN dcache_mem_i_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END dcache_mem_i_data[5]
  PIN dcache_mem_i_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END dcache_mem_i_data[6]
  PIN dcache_mem_i_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END dcache_mem_i_data[7]
  PIN dcache_mem_i_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END dcache_mem_i_data[8]
  PIN dcache_mem_i_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END dcache_mem_i_data[9]
  PIN dcache_mem_o_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END dcache_mem_o_data[0]
  PIN dcache_mem_o_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END dcache_mem_o_data[10]
  PIN dcache_mem_o_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END dcache_mem_o_data[11]
  PIN dcache_mem_o_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END dcache_mem_o_data[12]
  PIN dcache_mem_o_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END dcache_mem_o_data[13]
  PIN dcache_mem_o_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END dcache_mem_o_data[14]
  PIN dcache_mem_o_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END dcache_mem_o_data[15]
  PIN dcache_mem_o_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END dcache_mem_o_data[1]
  PIN dcache_mem_o_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END dcache_mem_o_data[2]
  PIN dcache_mem_o_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END dcache_mem_o_data[3]
  PIN dcache_mem_o_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END dcache_mem_o_data[4]
  PIN dcache_mem_o_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END dcache_mem_o_data[5]
  PIN dcache_mem_o_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END dcache_mem_o_data[6]
  PIN dcache_mem_o_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END dcache_mem_o_data[7]
  PIN dcache_mem_o_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END dcache_mem_o_data[8]
  PIN dcache_mem_o_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END dcache_mem_o_data[9]
  PIN dcache_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END dcache_mem_req
  PIN dcache_mem_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END dcache_mem_sel[0]
  PIN dcache_mem_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END dcache_mem_sel[1]
  PIN dcache_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END dcache_mem_we
  PIN dcache_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END dcache_rst
  PIN dcache_wb_4_burst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END dcache_wb_4_burst
  PIN dcache_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END dcache_wb_ack
  PIN dcache_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END dcache_wb_adr[0]
  PIN dcache_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END dcache_wb_adr[10]
  PIN dcache_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END dcache_wb_adr[11]
  PIN dcache_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END dcache_wb_adr[12]
  PIN dcache_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END dcache_wb_adr[13]
  PIN dcache_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END dcache_wb_adr[14]
  PIN dcache_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END dcache_wb_adr[15]
  PIN dcache_wb_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END dcache_wb_adr[16]
  PIN dcache_wb_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END dcache_wb_adr[17]
  PIN dcache_wb_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END dcache_wb_adr[18]
  PIN dcache_wb_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END dcache_wb_adr[19]
  PIN dcache_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END dcache_wb_adr[1]
  PIN dcache_wb_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END dcache_wb_adr[20]
  PIN dcache_wb_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END dcache_wb_adr[21]
  PIN dcache_wb_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END dcache_wb_adr[22]
  PIN dcache_wb_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END dcache_wb_adr[23]
  PIN dcache_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END dcache_wb_adr[2]
  PIN dcache_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END dcache_wb_adr[3]
  PIN dcache_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END dcache_wb_adr[4]
  PIN dcache_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END dcache_wb_adr[5]
  PIN dcache_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END dcache_wb_adr[6]
  PIN dcache_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END dcache_wb_adr[7]
  PIN dcache_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END dcache_wb_adr[8]
  PIN dcache_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END dcache_wb_adr[9]
  PIN dcache_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END dcache_wb_cyc
  PIN dcache_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END dcache_wb_err
  PIN dcache_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END dcache_wb_i_dat[0]
  PIN dcache_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END dcache_wb_i_dat[10]
  PIN dcache_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END dcache_wb_i_dat[11]
  PIN dcache_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END dcache_wb_i_dat[12]
  PIN dcache_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END dcache_wb_i_dat[13]
  PIN dcache_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END dcache_wb_i_dat[14]
  PIN dcache_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END dcache_wb_i_dat[15]
  PIN dcache_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END dcache_wb_i_dat[1]
  PIN dcache_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END dcache_wb_i_dat[2]
  PIN dcache_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END dcache_wb_i_dat[3]
  PIN dcache_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END dcache_wb_i_dat[4]
  PIN dcache_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END dcache_wb_i_dat[5]
  PIN dcache_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END dcache_wb_i_dat[6]
  PIN dcache_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END dcache_wb_i_dat[7]
  PIN dcache_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END dcache_wb_i_dat[8]
  PIN dcache_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END dcache_wb_i_dat[9]
  PIN dcache_wb_o_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END dcache_wb_o_dat[0]
  PIN dcache_wb_o_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END dcache_wb_o_dat[10]
  PIN dcache_wb_o_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END dcache_wb_o_dat[11]
  PIN dcache_wb_o_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END dcache_wb_o_dat[12]
  PIN dcache_wb_o_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END dcache_wb_o_dat[13]
  PIN dcache_wb_o_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END dcache_wb_o_dat[14]
  PIN dcache_wb_o_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END dcache_wb_o_dat[15]
  PIN dcache_wb_o_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END dcache_wb_o_dat[1]
  PIN dcache_wb_o_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END dcache_wb_o_dat[2]
  PIN dcache_wb_o_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END dcache_wb_o_dat[3]
  PIN dcache_wb_o_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END dcache_wb_o_dat[4]
  PIN dcache_wb_o_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END dcache_wb_o_dat[5]
  PIN dcache_wb_o_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END dcache_wb_o_dat[6]
  PIN dcache_wb_o_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END dcache_wb_o_dat[7]
  PIN dcache_wb_o_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END dcache_wb_o_dat[8]
  PIN dcache_wb_o_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END dcache_wb_o_dat[9]
  PIN dcache_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END dcache_wb_sel[0]
  PIN dcache_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END dcache_wb_sel[1]
  PIN dcache_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END dcache_wb_stb
  PIN dcache_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END dcache_wb_we
  PIN ic0_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.800 300.000 22.400 ;
    END
  END ic0_clk
  PIN ic0_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 25.880 300.000 26.480 ;
    END
  END ic0_mem_ack
  PIN ic0_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 66.680 300.000 67.280 ;
    END
  END ic0_mem_addr[0]
  PIN ic0_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 238.040 300.000 238.640 ;
    END
  END ic0_mem_addr[10]
  PIN ic0_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.360 300.000 254.960 ;
    END
  END ic0_mem_addr[11]
  PIN ic0_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.680 300.000 271.280 ;
    END
  END ic0_mem_addr[12]
  PIN ic0_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 287.000 300.000 287.600 ;
    END
  END ic0_mem_addr[13]
  PIN ic0_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 303.320 300.000 303.920 ;
    END
  END ic0_mem_addr[14]
  PIN ic0_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 319.640 300.000 320.240 ;
    END
  END ic0_mem_addr[15]
  PIN ic0_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.080 300.000 87.680 ;
    END
  END ic0_mem_addr[1]
  PIN ic0_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.480 300.000 108.080 ;
    END
  END ic0_mem_addr[2]
  PIN ic0_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.800 300.000 124.400 ;
    END
  END ic0_mem_addr[3]
  PIN ic0_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 140.120 300.000 140.720 ;
    END
  END ic0_mem_addr[4]
  PIN ic0_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.440 300.000 157.040 ;
    END
  END ic0_mem_addr[5]
  PIN ic0_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.760 300.000 173.360 ;
    END
  END ic0_mem_addr[6]
  PIN ic0_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 189.080 300.000 189.680 ;
    END
  END ic0_mem_addr[7]
  PIN ic0_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.400 300.000 206.000 ;
    END
  END ic0_mem_addr[8]
  PIN ic0_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.720 300.000 222.320 ;
    END
  END ic0_mem_addr[9]
  PIN ic0_mem_cache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.960 300.000 30.560 ;
    END
  END ic0_mem_cache_flush
  PIN ic0_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.760 300.000 71.360 ;
    END
  END ic0_mem_data[0]
  PIN ic0_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.120 300.000 242.720 ;
    END
  END ic0_mem_data[10]
  PIN ic0_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END ic0_mem_data[11]
  PIN ic0_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.760 300.000 275.360 ;
    END
  END ic0_mem_data[12]
  PIN ic0_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 291.080 300.000 291.680 ;
    END
  END ic0_mem_data[13]
  PIN ic0_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 307.400 300.000 308.000 ;
    END
  END ic0_mem_data[14]
  PIN ic0_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 323.720 300.000 324.320 ;
    END
  END ic0_mem_data[15]
  PIN ic0_mem_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 335.960 300.000 336.560 ;
    END
  END ic0_mem_data[16]
  PIN ic0_mem_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 340.040 300.000 340.640 ;
    END
  END ic0_mem_data[17]
  PIN ic0_mem_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 344.120 300.000 344.720 ;
    END
  END ic0_mem_data[18]
  PIN ic0_mem_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 348.200 300.000 348.800 ;
    END
  END ic0_mem_data[19]
  PIN ic0_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.160 300.000 91.760 ;
    END
  END ic0_mem_data[1]
  PIN ic0_mem_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 352.280 300.000 352.880 ;
    END
  END ic0_mem_data[20]
  PIN ic0_mem_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 356.360 300.000 356.960 ;
    END
  END ic0_mem_data[21]
  PIN ic0_mem_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 360.440 300.000 361.040 ;
    END
  END ic0_mem_data[22]
  PIN ic0_mem_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 364.520 300.000 365.120 ;
    END
  END ic0_mem_data[23]
  PIN ic0_mem_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 368.600 300.000 369.200 ;
    END
  END ic0_mem_data[24]
  PIN ic0_mem_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 372.680 300.000 373.280 ;
    END
  END ic0_mem_data[25]
  PIN ic0_mem_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 376.760 300.000 377.360 ;
    END
  END ic0_mem_data[26]
  PIN ic0_mem_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 380.840 300.000 381.440 ;
    END
  END ic0_mem_data[27]
  PIN ic0_mem_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 384.920 300.000 385.520 ;
    END
  END ic0_mem_data[28]
  PIN ic0_mem_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 389.000 300.000 389.600 ;
    END
  END ic0_mem_data[29]
  PIN ic0_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.560 300.000 112.160 ;
    END
  END ic0_mem_data[2]
  PIN ic0_mem_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 393.080 300.000 393.680 ;
    END
  END ic0_mem_data[30]
  PIN ic0_mem_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 397.160 300.000 397.760 ;
    END
  END ic0_mem_data[31]
  PIN ic0_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.880 300.000 128.480 ;
    END
  END ic0_mem_data[3]
  PIN ic0_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.200 300.000 144.800 ;
    END
  END ic0_mem_data[4]
  PIN ic0_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.520 300.000 161.120 ;
    END
  END ic0_mem_data[5]
  PIN ic0_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END ic0_mem_data[6]
  PIN ic0_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.160 300.000 193.760 ;
    END
  END ic0_mem_data[7]
  PIN ic0_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.480 300.000 210.080 ;
    END
  END ic0_mem_data[8]
  PIN ic0_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.800 300.000 226.400 ;
    END
  END ic0_mem_data[9]
  PIN ic0_mem_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.040 300.000 34.640 ;
    END
  END ic0_mem_ppl_submit
  PIN ic0_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 38.120 300.000 38.720 ;
    END
  END ic0_mem_req
  PIN ic0_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.200 300.000 42.800 ;
    END
  END ic0_rst
  PIN ic0_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 46.280 300.000 46.880 ;
    END
  END ic0_wb_ack
  PIN ic0_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.840 300.000 75.440 ;
    END
  END ic0_wb_adr[0]
  PIN ic0_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 246.200 300.000 246.800 ;
    END
  END ic0_wb_adr[10]
  PIN ic0_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.520 300.000 263.120 ;
    END
  END ic0_wb_adr[11]
  PIN ic0_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 278.840 300.000 279.440 ;
    END
  END ic0_wb_adr[12]
  PIN ic0_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.160 300.000 295.760 ;
    END
  END ic0_wb_adr[13]
  PIN ic0_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 311.480 300.000 312.080 ;
    END
  END ic0_wb_adr[14]
  PIN ic0_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 327.800 300.000 328.400 ;
    END
  END ic0_wb_adr[15]
  PIN ic0_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END ic0_wb_adr[1]
  PIN ic0_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.640 300.000 116.240 ;
    END
  END ic0_wb_adr[2]
  PIN ic0_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 131.960 300.000 132.560 ;
    END
  END ic0_wb_adr[3]
  PIN ic0_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.280 300.000 148.880 ;
    END
  END ic0_wb_adr[4]
  PIN ic0_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.600 300.000 165.200 ;
    END
  END ic0_wb_adr[5]
  PIN ic0_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.920 300.000 181.520 ;
    END
  END ic0_wb_adr[6]
  PIN ic0_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 197.240 300.000 197.840 ;
    END
  END ic0_wb_adr[7]
  PIN ic0_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.560 300.000 214.160 ;
    END
  END ic0_wb_adr[8]
  PIN ic0_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.880 300.000 230.480 ;
    END
  END ic0_wb_adr[9]
  PIN ic0_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.360 300.000 50.960 ;
    END
  END ic0_wb_cyc
  PIN ic0_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.440 300.000 55.040 ;
    END
  END ic0_wb_err
  PIN ic0_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.920 300.000 79.520 ;
    END
  END ic0_wb_i_dat[0]
  PIN ic0_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.280 300.000 250.880 ;
    END
  END ic0_wb_i_dat[10]
  PIN ic0_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.600 300.000 267.200 ;
    END
  END ic0_wb_i_dat[11]
  PIN ic0_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.920 300.000 283.520 ;
    END
  END ic0_wb_i_dat[12]
  PIN ic0_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 299.240 300.000 299.840 ;
    END
  END ic0_wb_i_dat[13]
  PIN ic0_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 315.560 300.000 316.160 ;
    END
  END ic0_wb_i_dat[14]
  PIN ic0_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 331.880 300.000 332.480 ;
    END
  END ic0_wb_i_dat[15]
  PIN ic0_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.320 300.000 99.920 ;
    END
  END ic0_wb_i_dat[1]
  PIN ic0_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.720 300.000 120.320 ;
    END
  END ic0_wb_i_dat[2]
  PIN ic0_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END ic0_wb_i_dat[3]
  PIN ic0_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.360 300.000 152.960 ;
    END
  END ic0_wb_i_dat[4]
  PIN ic0_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.680 300.000 169.280 ;
    END
  END ic0_wb_i_dat[5]
  PIN ic0_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.000 300.000 185.600 ;
    END
  END ic0_wb_i_dat[6]
  PIN ic0_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END ic0_wb_i_dat[7]
  PIN ic0_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 217.640 300.000 218.240 ;
    END
  END ic0_wb_i_dat[8]
  PIN ic0_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 233.960 300.000 234.560 ;
    END
  END ic0_wb_i_dat[9]
  PIN ic0_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.000 300.000 83.600 ;
    END
  END ic0_wb_sel[0]
  PIN ic0_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 103.400 300.000 104.000 ;
    END
  END ic0_wb_sel[1]
  PIN ic0_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 58.520 300.000 59.120 ;
    END
  END ic0_wb_stb
  PIN ic0_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.600 300.000 63.200 ;
    END
  END ic0_wb_we
  PIN ic1_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 401.240 300.000 401.840 ;
    END
  END ic1_clk
  PIN ic1_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 405.320 300.000 405.920 ;
    END
  END ic1_mem_ack
  PIN ic1_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 446.120 300.000 446.720 ;
    END
  END ic1_mem_addr[0]
  PIN ic1_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 617.480 300.000 618.080 ;
    END
  END ic1_mem_addr[10]
  PIN ic1_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 633.800 300.000 634.400 ;
    END
  END ic1_mem_addr[11]
  PIN ic1_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 650.120 300.000 650.720 ;
    END
  END ic1_mem_addr[12]
  PIN ic1_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 666.440 300.000 667.040 ;
    END
  END ic1_mem_addr[13]
  PIN ic1_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 682.760 300.000 683.360 ;
    END
  END ic1_mem_addr[14]
  PIN ic1_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 699.080 300.000 699.680 ;
    END
  END ic1_mem_addr[15]
  PIN ic1_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 466.520 300.000 467.120 ;
    END
  END ic1_mem_addr[1]
  PIN ic1_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 486.920 300.000 487.520 ;
    END
  END ic1_mem_addr[2]
  PIN ic1_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 503.240 300.000 503.840 ;
    END
  END ic1_mem_addr[3]
  PIN ic1_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 519.560 300.000 520.160 ;
    END
  END ic1_mem_addr[4]
  PIN ic1_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 535.880 300.000 536.480 ;
    END
  END ic1_mem_addr[5]
  PIN ic1_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 552.200 300.000 552.800 ;
    END
  END ic1_mem_addr[6]
  PIN ic1_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 568.520 300.000 569.120 ;
    END
  END ic1_mem_addr[7]
  PIN ic1_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 584.840 300.000 585.440 ;
    END
  END ic1_mem_addr[8]
  PIN ic1_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 601.160 300.000 601.760 ;
    END
  END ic1_mem_addr[9]
  PIN ic1_mem_cache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 409.400 300.000 410.000 ;
    END
  END ic1_mem_cache_flush
  PIN ic1_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 450.200 300.000 450.800 ;
    END
  END ic1_mem_data[0]
  PIN ic1_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 621.560 300.000 622.160 ;
    END
  END ic1_mem_data[10]
  PIN ic1_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 637.880 300.000 638.480 ;
    END
  END ic1_mem_data[11]
  PIN ic1_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 654.200 300.000 654.800 ;
    END
  END ic1_mem_data[12]
  PIN ic1_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 670.520 300.000 671.120 ;
    END
  END ic1_mem_data[13]
  PIN ic1_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 686.840 300.000 687.440 ;
    END
  END ic1_mem_data[14]
  PIN ic1_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 703.160 300.000 703.760 ;
    END
  END ic1_mem_data[15]
  PIN ic1_mem_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 715.400 300.000 716.000 ;
    END
  END ic1_mem_data[16]
  PIN ic1_mem_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 719.480 300.000 720.080 ;
    END
  END ic1_mem_data[17]
  PIN ic1_mem_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 723.560 300.000 724.160 ;
    END
  END ic1_mem_data[18]
  PIN ic1_mem_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 727.640 300.000 728.240 ;
    END
  END ic1_mem_data[19]
  PIN ic1_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 470.600 300.000 471.200 ;
    END
  END ic1_mem_data[1]
  PIN ic1_mem_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 731.720 300.000 732.320 ;
    END
  END ic1_mem_data[20]
  PIN ic1_mem_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 735.800 300.000 736.400 ;
    END
  END ic1_mem_data[21]
  PIN ic1_mem_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 739.880 300.000 740.480 ;
    END
  END ic1_mem_data[22]
  PIN ic1_mem_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 743.960 300.000 744.560 ;
    END
  END ic1_mem_data[23]
  PIN ic1_mem_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 748.040 300.000 748.640 ;
    END
  END ic1_mem_data[24]
  PIN ic1_mem_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 752.120 300.000 752.720 ;
    END
  END ic1_mem_data[25]
  PIN ic1_mem_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 756.200 300.000 756.800 ;
    END
  END ic1_mem_data[26]
  PIN ic1_mem_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 760.280 300.000 760.880 ;
    END
  END ic1_mem_data[27]
  PIN ic1_mem_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 764.360 300.000 764.960 ;
    END
  END ic1_mem_data[28]
  PIN ic1_mem_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 768.440 300.000 769.040 ;
    END
  END ic1_mem_data[29]
  PIN ic1_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 491.000 300.000 491.600 ;
    END
  END ic1_mem_data[2]
  PIN ic1_mem_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 772.520 300.000 773.120 ;
    END
  END ic1_mem_data[30]
  PIN ic1_mem_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 776.600 300.000 777.200 ;
    END
  END ic1_mem_data[31]
  PIN ic1_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 507.320 300.000 507.920 ;
    END
  END ic1_mem_data[3]
  PIN ic1_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 523.640 300.000 524.240 ;
    END
  END ic1_mem_data[4]
  PIN ic1_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 539.960 300.000 540.560 ;
    END
  END ic1_mem_data[5]
  PIN ic1_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 556.280 300.000 556.880 ;
    END
  END ic1_mem_data[6]
  PIN ic1_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 572.600 300.000 573.200 ;
    END
  END ic1_mem_data[7]
  PIN ic1_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 588.920 300.000 589.520 ;
    END
  END ic1_mem_data[8]
  PIN ic1_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 605.240 300.000 605.840 ;
    END
  END ic1_mem_data[9]
  PIN ic1_mem_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 413.480 300.000 414.080 ;
    END
  END ic1_mem_ppl_submit
  PIN ic1_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 417.560 300.000 418.160 ;
    END
  END ic1_mem_req
  PIN ic1_rst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 421.640 300.000 422.240 ;
    END
  END ic1_rst
  PIN ic1_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 425.720 300.000 426.320 ;
    END
  END ic1_wb_ack
  PIN ic1_wb_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 454.280 300.000 454.880 ;
    END
  END ic1_wb_adr[0]
  PIN ic1_wb_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 625.640 300.000 626.240 ;
    END
  END ic1_wb_adr[10]
  PIN ic1_wb_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 641.960 300.000 642.560 ;
    END
  END ic1_wb_adr[11]
  PIN ic1_wb_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 658.280 300.000 658.880 ;
    END
  END ic1_wb_adr[12]
  PIN ic1_wb_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 674.600 300.000 675.200 ;
    END
  END ic1_wb_adr[13]
  PIN ic1_wb_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 690.920 300.000 691.520 ;
    END
  END ic1_wb_adr[14]
  PIN ic1_wb_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 707.240 300.000 707.840 ;
    END
  END ic1_wb_adr[15]
  PIN ic1_wb_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 474.680 300.000 475.280 ;
    END
  END ic1_wb_adr[1]
  PIN ic1_wb_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 495.080 300.000 495.680 ;
    END
  END ic1_wb_adr[2]
  PIN ic1_wb_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 511.400 300.000 512.000 ;
    END
  END ic1_wb_adr[3]
  PIN ic1_wb_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 527.720 300.000 528.320 ;
    END
  END ic1_wb_adr[4]
  PIN ic1_wb_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 544.040 300.000 544.640 ;
    END
  END ic1_wb_adr[5]
  PIN ic1_wb_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 560.360 300.000 560.960 ;
    END
  END ic1_wb_adr[6]
  PIN ic1_wb_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 576.680 300.000 577.280 ;
    END
  END ic1_wb_adr[7]
  PIN ic1_wb_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 593.000 300.000 593.600 ;
    END
  END ic1_wb_adr[8]
  PIN ic1_wb_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 609.320 300.000 609.920 ;
    END
  END ic1_wb_adr[9]
  PIN ic1_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 429.800 300.000 430.400 ;
    END
  END ic1_wb_cyc
  PIN ic1_wb_err
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 433.880 300.000 434.480 ;
    END
  END ic1_wb_err
  PIN ic1_wb_i_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 458.360 300.000 458.960 ;
    END
  END ic1_wb_i_dat[0]
  PIN ic1_wb_i_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 629.720 300.000 630.320 ;
    END
  END ic1_wb_i_dat[10]
  PIN ic1_wb_i_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 646.040 300.000 646.640 ;
    END
  END ic1_wb_i_dat[11]
  PIN ic1_wb_i_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 662.360 300.000 662.960 ;
    END
  END ic1_wb_i_dat[12]
  PIN ic1_wb_i_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 678.680 300.000 679.280 ;
    END
  END ic1_wb_i_dat[13]
  PIN ic1_wb_i_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 695.000 300.000 695.600 ;
    END
  END ic1_wb_i_dat[14]
  PIN ic1_wb_i_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 711.320 300.000 711.920 ;
    END
  END ic1_wb_i_dat[15]
  PIN ic1_wb_i_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 478.760 300.000 479.360 ;
    END
  END ic1_wb_i_dat[1]
  PIN ic1_wb_i_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 499.160 300.000 499.760 ;
    END
  END ic1_wb_i_dat[2]
  PIN ic1_wb_i_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 515.480 300.000 516.080 ;
    END
  END ic1_wb_i_dat[3]
  PIN ic1_wb_i_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 531.800 300.000 532.400 ;
    END
  END ic1_wb_i_dat[4]
  PIN ic1_wb_i_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 548.120 300.000 548.720 ;
    END
  END ic1_wb_i_dat[5]
  PIN ic1_wb_i_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 564.440 300.000 565.040 ;
    END
  END ic1_wb_i_dat[6]
  PIN ic1_wb_i_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 580.760 300.000 581.360 ;
    END
  END ic1_wb_i_dat[7]
  PIN ic1_wb_i_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 597.080 300.000 597.680 ;
    END
  END ic1_wb_i_dat[8]
  PIN ic1_wb_i_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 613.400 300.000 614.000 ;
    END
  END ic1_wb_i_dat[9]
  PIN ic1_wb_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 462.440 300.000 463.040 ;
    END
  END ic1_wb_sel[0]
  PIN ic1_wb_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 482.840 300.000 483.440 ;
    END
  END ic1_wb_sel[1]
  PIN ic1_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 437.960 300.000 438.560 ;
    END
  END ic1_wb_stb
  PIN ic1_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 442.040 300.000 442.640 ;
    END
  END ic1_wb_we
  PIN inner_disable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 796.000 15.550 800.000 ;
    END
  END inner_disable
  PIN inner_embed_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 796.000 19.690 800.000 ;
    END
  END inner_embed_mode
  PIN inner_ext_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 796.000 23.830 800.000 ;
    END
  END inner_ext_irq
  PIN inner_wb_4_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 796.000 27.970 800.000 ;
    END
  END inner_wb_4_burst
  PIN inner_wb_8_burst
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 796.000 32.110 800.000 ;
    END
  END inner_wb_8_burst
  PIN inner_wb_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 796.000 36.250 800.000 ;
    END
  END inner_wb_ack
  PIN inner_wb_adr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 796.000 56.950 800.000 ;
    END
  END inner_wb_adr[0]
  PIN inner_wb_adr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 796.000 189.430 800.000 ;
    END
  END inner_wb_adr[10]
  PIN inner_wb_adr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 796.000 201.850 800.000 ;
    END
  END inner_wb_adr[11]
  PIN inner_wb_adr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 796.000 214.270 800.000 ;
    END
  END inner_wb_adr[12]
  PIN inner_wb_adr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 796.000 226.690 800.000 ;
    END
  END inner_wb_adr[13]
  PIN inner_wb_adr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 796.000 239.110 800.000 ;
    END
  END inner_wb_adr[14]
  PIN inner_wb_adr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 796.000 251.530 800.000 ;
    END
  END inner_wb_adr[15]
  PIN inner_wb_adr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 796.000 263.950 800.000 ;
    END
  END inner_wb_adr[16]
  PIN inner_wb_adr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 796.000 268.090 800.000 ;
    END
  END inner_wb_adr[17]
  PIN inner_wb_adr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 796.000 272.230 800.000 ;
    END
  END inner_wb_adr[18]
  PIN inner_wb_adr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 796.000 276.370 800.000 ;
    END
  END inner_wb_adr[19]
  PIN inner_wb_adr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 796.000 73.510 800.000 ;
    END
  END inner_wb_adr[1]
  PIN inner_wb_adr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 796.000 280.510 800.000 ;
    END
  END inner_wb_adr[20]
  PIN inner_wb_adr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 796.000 284.650 800.000 ;
    END
  END inner_wb_adr[21]
  PIN inner_wb_adr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 796.000 288.790 800.000 ;
    END
  END inner_wb_adr[22]
  PIN inner_wb_adr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 796.000 292.930 800.000 ;
    END
  END inner_wb_adr[23]
  PIN inner_wb_adr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 796.000 90.070 800.000 ;
    END
  END inner_wb_adr[2]
  PIN inner_wb_adr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 796.000 102.490 800.000 ;
    END
  END inner_wb_adr[3]
  PIN inner_wb_adr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 796.000 114.910 800.000 ;
    END
  END inner_wb_adr[4]
  PIN inner_wb_adr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 796.000 127.330 800.000 ;
    END
  END inner_wb_adr[5]
  PIN inner_wb_adr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 796.000 139.750 800.000 ;
    END
  END inner_wb_adr[6]
  PIN inner_wb_adr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 796.000 152.170 800.000 ;
    END
  END inner_wb_adr[7]
  PIN inner_wb_adr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 796.000 164.590 800.000 ;
    END
  END inner_wb_adr[8]
  PIN inner_wb_adr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 796.000 177.010 800.000 ;
    END
  END inner_wb_adr[9]
  PIN inner_wb_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 796.000 40.390 800.000 ;
    END
  END inner_wb_cyc
  PIN inner_wb_err
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 796.000 44.530 800.000 ;
    END
  END inner_wb_err
  PIN inner_wb_i_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 796.000 61.090 800.000 ;
    END
  END inner_wb_i_dat[0]
  PIN inner_wb_i_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 796.000 193.570 800.000 ;
    END
  END inner_wb_i_dat[10]
  PIN inner_wb_i_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 796.000 205.990 800.000 ;
    END
  END inner_wb_i_dat[11]
  PIN inner_wb_i_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 796.000 218.410 800.000 ;
    END
  END inner_wb_i_dat[12]
  PIN inner_wb_i_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 796.000 230.830 800.000 ;
    END
  END inner_wb_i_dat[13]
  PIN inner_wb_i_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 796.000 243.250 800.000 ;
    END
  END inner_wb_i_dat[14]
  PIN inner_wb_i_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 796.000 255.670 800.000 ;
    END
  END inner_wb_i_dat[15]
  PIN inner_wb_i_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 796.000 77.650 800.000 ;
    END
  END inner_wb_i_dat[1]
  PIN inner_wb_i_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 796.000 94.210 800.000 ;
    END
  END inner_wb_i_dat[2]
  PIN inner_wb_i_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 796.000 106.630 800.000 ;
    END
  END inner_wb_i_dat[3]
  PIN inner_wb_i_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 796.000 119.050 800.000 ;
    END
  END inner_wb_i_dat[4]
  PIN inner_wb_i_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 796.000 131.470 800.000 ;
    END
  END inner_wb_i_dat[5]
  PIN inner_wb_i_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 796.000 143.890 800.000 ;
    END
  END inner_wb_i_dat[6]
  PIN inner_wb_i_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 796.000 156.310 800.000 ;
    END
  END inner_wb_i_dat[7]
  PIN inner_wb_i_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 796.000 168.730 800.000 ;
    END
  END inner_wb_i_dat[8]
  PIN inner_wb_i_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 796.000 181.150 800.000 ;
    END
  END inner_wb_i_dat[9]
  PIN inner_wb_o_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 796.000 65.230 800.000 ;
    END
  END inner_wb_o_dat[0]
  PIN inner_wb_o_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 796.000 197.710 800.000 ;
    END
  END inner_wb_o_dat[10]
  PIN inner_wb_o_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 796.000 210.130 800.000 ;
    END
  END inner_wb_o_dat[11]
  PIN inner_wb_o_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 796.000 222.550 800.000 ;
    END
  END inner_wb_o_dat[12]
  PIN inner_wb_o_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 796.000 234.970 800.000 ;
    END
  END inner_wb_o_dat[13]
  PIN inner_wb_o_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 796.000 247.390 800.000 ;
    END
  END inner_wb_o_dat[14]
  PIN inner_wb_o_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 796.000 259.810 800.000 ;
    END
  END inner_wb_o_dat[15]
  PIN inner_wb_o_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 796.000 81.790 800.000 ;
    END
  END inner_wb_o_dat[1]
  PIN inner_wb_o_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 796.000 98.350 800.000 ;
    END
  END inner_wb_o_dat[2]
  PIN inner_wb_o_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 796.000 110.770 800.000 ;
    END
  END inner_wb_o_dat[3]
  PIN inner_wb_o_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 796.000 123.190 800.000 ;
    END
  END inner_wb_o_dat[4]
  PIN inner_wb_o_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 796.000 135.610 800.000 ;
    END
  END inner_wb_o_dat[5]
  PIN inner_wb_o_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 796.000 148.030 800.000 ;
    END
  END inner_wb_o_dat[6]
  PIN inner_wb_o_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 796.000 160.450 800.000 ;
    END
  END inner_wb_o_dat[7]
  PIN inner_wb_o_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 796.000 172.870 800.000 ;
    END
  END inner_wb_o_dat[8]
  PIN inner_wb_o_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 796.000 185.290 800.000 ;
    END
  END inner_wb_o_dat[9]
  PIN inner_wb_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 796.000 69.370 800.000 ;
    END
  END inner_wb_sel[0]
  PIN inner_wb_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 796.000 85.930 800.000 ;
    END
  END inner_wb_sel[1]
  PIN inner_wb_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 796.000 48.670 800.000 ;
    END
  END inner_wb_stb
  PIN inner_wb_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 796.000 52.810 800.000 ;
    END
  END inner_wb_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 788.885 ;
      LAYER met1 ;
        RECT 1.450 10.240 299.850 793.180 ;
      LAYER met2 ;
        RECT 1.480 795.720 6.710 796.690 ;
        RECT 7.550 795.720 10.850 796.690 ;
        RECT 11.690 795.720 14.990 796.690 ;
        RECT 15.830 795.720 19.130 796.690 ;
        RECT 19.970 795.720 23.270 796.690 ;
        RECT 24.110 795.720 27.410 796.690 ;
        RECT 28.250 795.720 31.550 796.690 ;
        RECT 32.390 795.720 35.690 796.690 ;
        RECT 36.530 795.720 39.830 796.690 ;
        RECT 40.670 795.720 43.970 796.690 ;
        RECT 44.810 795.720 48.110 796.690 ;
        RECT 48.950 795.720 52.250 796.690 ;
        RECT 53.090 795.720 56.390 796.690 ;
        RECT 57.230 795.720 60.530 796.690 ;
        RECT 61.370 795.720 64.670 796.690 ;
        RECT 65.510 795.720 68.810 796.690 ;
        RECT 69.650 795.720 72.950 796.690 ;
        RECT 73.790 795.720 77.090 796.690 ;
        RECT 77.930 795.720 81.230 796.690 ;
        RECT 82.070 795.720 85.370 796.690 ;
        RECT 86.210 795.720 89.510 796.690 ;
        RECT 90.350 795.720 93.650 796.690 ;
        RECT 94.490 795.720 97.790 796.690 ;
        RECT 98.630 795.720 101.930 796.690 ;
        RECT 102.770 795.720 106.070 796.690 ;
        RECT 106.910 795.720 110.210 796.690 ;
        RECT 111.050 795.720 114.350 796.690 ;
        RECT 115.190 795.720 118.490 796.690 ;
        RECT 119.330 795.720 122.630 796.690 ;
        RECT 123.470 795.720 126.770 796.690 ;
        RECT 127.610 795.720 130.910 796.690 ;
        RECT 131.750 795.720 135.050 796.690 ;
        RECT 135.890 795.720 139.190 796.690 ;
        RECT 140.030 795.720 143.330 796.690 ;
        RECT 144.170 795.720 147.470 796.690 ;
        RECT 148.310 795.720 151.610 796.690 ;
        RECT 152.450 795.720 155.750 796.690 ;
        RECT 156.590 795.720 159.890 796.690 ;
        RECT 160.730 795.720 164.030 796.690 ;
        RECT 164.870 795.720 168.170 796.690 ;
        RECT 169.010 795.720 172.310 796.690 ;
        RECT 173.150 795.720 176.450 796.690 ;
        RECT 177.290 795.720 180.590 796.690 ;
        RECT 181.430 795.720 184.730 796.690 ;
        RECT 185.570 795.720 188.870 796.690 ;
        RECT 189.710 795.720 193.010 796.690 ;
        RECT 193.850 795.720 197.150 796.690 ;
        RECT 197.990 795.720 201.290 796.690 ;
        RECT 202.130 795.720 205.430 796.690 ;
        RECT 206.270 795.720 209.570 796.690 ;
        RECT 210.410 795.720 213.710 796.690 ;
        RECT 214.550 795.720 217.850 796.690 ;
        RECT 218.690 795.720 221.990 796.690 ;
        RECT 222.830 795.720 226.130 796.690 ;
        RECT 226.970 795.720 230.270 796.690 ;
        RECT 231.110 795.720 234.410 796.690 ;
        RECT 235.250 795.720 238.550 796.690 ;
        RECT 239.390 795.720 242.690 796.690 ;
        RECT 243.530 795.720 246.830 796.690 ;
        RECT 247.670 795.720 250.970 796.690 ;
        RECT 251.810 795.720 255.110 796.690 ;
        RECT 255.950 795.720 259.250 796.690 ;
        RECT 260.090 795.720 263.390 796.690 ;
        RECT 264.230 795.720 267.530 796.690 ;
        RECT 268.370 795.720 271.670 796.690 ;
        RECT 272.510 795.720 275.810 796.690 ;
        RECT 276.650 795.720 279.950 796.690 ;
        RECT 280.790 795.720 284.090 796.690 ;
        RECT 284.930 795.720 288.230 796.690 ;
        RECT 289.070 795.720 292.370 796.690 ;
        RECT 293.210 795.720 299.820 796.690 ;
        RECT 1.480 4.280 299.820 795.720 ;
        RECT 1.480 3.670 2.110 4.280 ;
        RECT 2.950 3.670 4.410 4.280 ;
        RECT 5.250 3.670 6.710 4.280 ;
        RECT 7.550 3.670 9.010 4.280 ;
        RECT 9.850 3.670 11.310 4.280 ;
        RECT 12.150 3.670 13.610 4.280 ;
        RECT 14.450 3.670 15.910 4.280 ;
        RECT 16.750 3.670 18.210 4.280 ;
        RECT 19.050 3.670 20.510 4.280 ;
        RECT 21.350 3.670 22.810 4.280 ;
        RECT 23.650 3.670 25.110 4.280 ;
        RECT 25.950 3.670 27.410 4.280 ;
        RECT 28.250 3.670 29.710 4.280 ;
        RECT 30.550 3.670 32.010 4.280 ;
        RECT 32.850 3.670 34.310 4.280 ;
        RECT 35.150 3.670 36.610 4.280 ;
        RECT 37.450 3.670 38.910 4.280 ;
        RECT 39.750 3.670 41.210 4.280 ;
        RECT 42.050 3.670 43.510 4.280 ;
        RECT 44.350 3.670 45.810 4.280 ;
        RECT 46.650 3.670 48.110 4.280 ;
        RECT 48.950 3.670 50.410 4.280 ;
        RECT 51.250 3.670 52.710 4.280 ;
        RECT 53.550 3.670 55.010 4.280 ;
        RECT 55.850 3.670 57.310 4.280 ;
        RECT 58.150 3.670 59.610 4.280 ;
        RECT 60.450 3.670 61.910 4.280 ;
        RECT 62.750 3.670 64.210 4.280 ;
        RECT 65.050 3.670 66.510 4.280 ;
        RECT 67.350 3.670 68.810 4.280 ;
        RECT 69.650 3.670 71.110 4.280 ;
        RECT 71.950 3.670 73.410 4.280 ;
        RECT 74.250 3.670 75.710 4.280 ;
        RECT 76.550 3.670 78.010 4.280 ;
        RECT 78.850 3.670 80.310 4.280 ;
        RECT 81.150 3.670 82.610 4.280 ;
        RECT 83.450 3.670 84.910 4.280 ;
        RECT 85.750 3.670 87.210 4.280 ;
        RECT 88.050 3.670 89.510 4.280 ;
        RECT 90.350 3.670 91.810 4.280 ;
        RECT 92.650 3.670 94.110 4.280 ;
        RECT 94.950 3.670 96.410 4.280 ;
        RECT 97.250 3.670 98.710 4.280 ;
        RECT 99.550 3.670 101.010 4.280 ;
        RECT 101.850 3.670 103.310 4.280 ;
        RECT 104.150 3.670 105.610 4.280 ;
        RECT 106.450 3.670 107.910 4.280 ;
        RECT 108.750 3.670 110.210 4.280 ;
        RECT 111.050 3.670 112.510 4.280 ;
        RECT 113.350 3.670 114.810 4.280 ;
        RECT 115.650 3.670 117.110 4.280 ;
        RECT 117.950 3.670 119.410 4.280 ;
        RECT 120.250 3.670 121.710 4.280 ;
        RECT 122.550 3.670 124.010 4.280 ;
        RECT 124.850 3.670 126.310 4.280 ;
        RECT 127.150 3.670 128.610 4.280 ;
        RECT 129.450 3.670 130.910 4.280 ;
        RECT 131.750 3.670 133.210 4.280 ;
        RECT 134.050 3.670 135.510 4.280 ;
        RECT 136.350 3.670 137.810 4.280 ;
        RECT 138.650 3.670 140.110 4.280 ;
        RECT 140.950 3.670 142.410 4.280 ;
        RECT 143.250 3.670 144.710 4.280 ;
        RECT 145.550 3.670 147.010 4.280 ;
        RECT 147.850 3.670 149.310 4.280 ;
        RECT 150.150 3.670 151.610 4.280 ;
        RECT 152.450 3.670 153.910 4.280 ;
        RECT 154.750 3.670 156.210 4.280 ;
        RECT 157.050 3.670 158.510 4.280 ;
        RECT 159.350 3.670 160.810 4.280 ;
        RECT 161.650 3.670 163.110 4.280 ;
        RECT 163.950 3.670 165.410 4.280 ;
        RECT 166.250 3.670 167.710 4.280 ;
        RECT 168.550 3.670 170.010 4.280 ;
        RECT 170.850 3.670 172.310 4.280 ;
        RECT 173.150 3.670 174.610 4.280 ;
        RECT 175.450 3.670 176.910 4.280 ;
        RECT 177.750 3.670 179.210 4.280 ;
        RECT 180.050 3.670 181.510 4.280 ;
        RECT 182.350 3.670 183.810 4.280 ;
        RECT 184.650 3.670 186.110 4.280 ;
        RECT 186.950 3.670 188.410 4.280 ;
        RECT 189.250 3.670 190.710 4.280 ;
        RECT 191.550 3.670 193.010 4.280 ;
        RECT 193.850 3.670 195.310 4.280 ;
        RECT 196.150 3.670 197.610 4.280 ;
        RECT 198.450 3.670 199.910 4.280 ;
        RECT 200.750 3.670 202.210 4.280 ;
        RECT 203.050 3.670 204.510 4.280 ;
        RECT 205.350 3.670 206.810 4.280 ;
        RECT 207.650 3.670 209.110 4.280 ;
        RECT 209.950 3.670 211.410 4.280 ;
        RECT 212.250 3.670 213.710 4.280 ;
        RECT 214.550 3.670 216.010 4.280 ;
        RECT 216.850 3.670 218.310 4.280 ;
        RECT 219.150 3.670 220.610 4.280 ;
        RECT 221.450 3.670 222.910 4.280 ;
        RECT 223.750 3.670 225.210 4.280 ;
        RECT 226.050 3.670 227.510 4.280 ;
        RECT 228.350 3.670 229.810 4.280 ;
        RECT 230.650 3.670 232.110 4.280 ;
        RECT 232.950 3.670 234.410 4.280 ;
        RECT 235.250 3.670 236.710 4.280 ;
        RECT 237.550 3.670 239.010 4.280 ;
        RECT 239.850 3.670 241.310 4.280 ;
        RECT 242.150 3.670 243.610 4.280 ;
        RECT 244.450 3.670 245.910 4.280 ;
        RECT 246.750 3.670 248.210 4.280 ;
        RECT 249.050 3.670 250.510 4.280 ;
        RECT 251.350 3.670 252.810 4.280 ;
        RECT 253.650 3.670 255.110 4.280 ;
        RECT 255.950 3.670 257.410 4.280 ;
        RECT 258.250 3.670 259.710 4.280 ;
        RECT 260.550 3.670 262.010 4.280 ;
        RECT 262.850 3.670 264.310 4.280 ;
        RECT 265.150 3.670 266.610 4.280 ;
        RECT 267.450 3.670 268.910 4.280 ;
        RECT 269.750 3.670 271.210 4.280 ;
        RECT 272.050 3.670 273.510 4.280 ;
        RECT 274.350 3.670 275.810 4.280 ;
        RECT 276.650 3.670 278.110 4.280 ;
        RECT 278.950 3.670 280.410 4.280 ;
        RECT 281.250 3.670 282.710 4.280 ;
        RECT 283.550 3.670 285.010 4.280 ;
        RECT 285.850 3.670 287.310 4.280 ;
        RECT 288.150 3.670 289.610 4.280 ;
        RECT 290.450 3.670 291.910 4.280 ;
        RECT 292.750 3.670 294.210 4.280 ;
        RECT 295.050 3.670 296.510 4.280 ;
        RECT 297.350 3.670 299.820 4.280 ;
      LAYER met3 ;
        RECT 3.030 777.600 296.000 788.965 ;
        RECT 3.030 776.200 295.600 777.600 ;
        RECT 3.030 773.520 296.000 776.200 ;
        RECT 3.030 772.120 295.600 773.520 ;
        RECT 3.030 769.440 296.000 772.120 ;
        RECT 3.030 768.040 295.600 769.440 ;
        RECT 3.030 765.360 296.000 768.040 ;
        RECT 3.030 763.960 295.600 765.360 ;
        RECT 3.030 761.280 296.000 763.960 ;
        RECT 3.030 759.880 295.600 761.280 ;
        RECT 3.030 757.200 296.000 759.880 ;
        RECT 3.030 755.800 295.600 757.200 ;
        RECT 3.030 753.120 296.000 755.800 ;
        RECT 3.030 751.720 295.600 753.120 ;
        RECT 3.030 749.040 296.000 751.720 ;
        RECT 3.030 747.640 295.600 749.040 ;
        RECT 3.030 744.960 296.000 747.640 ;
        RECT 3.030 743.560 295.600 744.960 ;
        RECT 3.030 740.880 296.000 743.560 ;
        RECT 3.030 739.480 295.600 740.880 ;
        RECT 3.030 736.800 296.000 739.480 ;
        RECT 3.030 735.400 295.600 736.800 ;
        RECT 3.030 732.720 296.000 735.400 ;
        RECT 3.030 731.320 295.600 732.720 ;
        RECT 3.030 728.640 296.000 731.320 ;
        RECT 3.030 727.240 295.600 728.640 ;
        RECT 3.030 724.560 296.000 727.240 ;
        RECT 3.030 723.160 295.600 724.560 ;
        RECT 3.030 720.480 296.000 723.160 ;
        RECT 3.030 719.080 295.600 720.480 ;
        RECT 3.030 716.400 296.000 719.080 ;
        RECT 3.030 715.000 295.600 716.400 ;
        RECT 3.030 712.320 296.000 715.000 ;
        RECT 3.030 710.920 295.600 712.320 ;
        RECT 3.030 708.240 296.000 710.920 ;
        RECT 3.030 706.840 295.600 708.240 ;
        RECT 3.030 704.160 296.000 706.840 ;
        RECT 3.030 702.760 295.600 704.160 ;
        RECT 3.030 700.080 296.000 702.760 ;
        RECT 3.030 698.680 295.600 700.080 ;
        RECT 3.030 696.000 296.000 698.680 ;
        RECT 3.030 694.600 295.600 696.000 ;
        RECT 3.030 691.920 296.000 694.600 ;
        RECT 3.030 690.520 295.600 691.920 ;
        RECT 3.030 687.840 296.000 690.520 ;
        RECT 4.400 686.440 295.600 687.840 ;
        RECT 4.400 683.760 296.000 686.440 ;
        RECT 4.400 682.360 295.600 683.760 ;
        RECT 4.400 679.680 296.000 682.360 ;
        RECT 4.400 678.280 295.600 679.680 ;
        RECT 4.400 675.600 296.000 678.280 ;
        RECT 4.400 674.200 295.600 675.600 ;
        RECT 4.400 671.520 296.000 674.200 ;
        RECT 4.400 670.120 295.600 671.520 ;
        RECT 4.400 667.440 296.000 670.120 ;
        RECT 4.400 666.040 295.600 667.440 ;
        RECT 4.400 663.360 296.000 666.040 ;
        RECT 4.400 661.960 295.600 663.360 ;
        RECT 4.400 659.280 296.000 661.960 ;
        RECT 4.400 657.880 295.600 659.280 ;
        RECT 4.400 655.200 296.000 657.880 ;
        RECT 4.400 653.800 295.600 655.200 ;
        RECT 4.400 651.120 296.000 653.800 ;
        RECT 4.400 649.720 295.600 651.120 ;
        RECT 4.400 647.040 296.000 649.720 ;
        RECT 4.400 645.640 295.600 647.040 ;
        RECT 4.400 642.960 296.000 645.640 ;
        RECT 4.400 641.560 295.600 642.960 ;
        RECT 4.400 638.880 296.000 641.560 ;
        RECT 4.400 637.480 295.600 638.880 ;
        RECT 4.400 634.800 296.000 637.480 ;
        RECT 4.400 633.400 295.600 634.800 ;
        RECT 4.400 630.720 296.000 633.400 ;
        RECT 4.400 629.320 295.600 630.720 ;
        RECT 4.400 626.640 296.000 629.320 ;
        RECT 4.400 625.240 295.600 626.640 ;
        RECT 4.400 622.560 296.000 625.240 ;
        RECT 4.400 621.160 295.600 622.560 ;
        RECT 4.400 618.480 296.000 621.160 ;
        RECT 4.400 617.080 295.600 618.480 ;
        RECT 4.400 614.400 296.000 617.080 ;
        RECT 4.400 613.000 295.600 614.400 ;
        RECT 4.400 610.320 296.000 613.000 ;
        RECT 4.400 608.920 295.600 610.320 ;
        RECT 4.400 606.240 296.000 608.920 ;
        RECT 4.400 604.840 295.600 606.240 ;
        RECT 4.400 602.160 296.000 604.840 ;
        RECT 4.400 600.760 295.600 602.160 ;
        RECT 4.400 598.080 296.000 600.760 ;
        RECT 4.400 596.680 295.600 598.080 ;
        RECT 4.400 594.000 296.000 596.680 ;
        RECT 4.400 592.600 295.600 594.000 ;
        RECT 4.400 589.920 296.000 592.600 ;
        RECT 4.400 588.520 295.600 589.920 ;
        RECT 4.400 585.840 296.000 588.520 ;
        RECT 4.400 584.440 295.600 585.840 ;
        RECT 4.400 581.760 296.000 584.440 ;
        RECT 4.400 580.360 295.600 581.760 ;
        RECT 4.400 577.680 296.000 580.360 ;
        RECT 4.400 576.280 295.600 577.680 ;
        RECT 4.400 573.600 296.000 576.280 ;
        RECT 4.400 572.200 295.600 573.600 ;
        RECT 4.400 569.520 296.000 572.200 ;
        RECT 4.400 568.120 295.600 569.520 ;
        RECT 4.400 565.440 296.000 568.120 ;
        RECT 4.400 564.040 295.600 565.440 ;
        RECT 4.400 561.360 296.000 564.040 ;
        RECT 4.400 559.960 295.600 561.360 ;
        RECT 4.400 557.280 296.000 559.960 ;
        RECT 4.400 555.880 295.600 557.280 ;
        RECT 4.400 553.200 296.000 555.880 ;
        RECT 4.400 551.800 295.600 553.200 ;
        RECT 4.400 549.120 296.000 551.800 ;
        RECT 4.400 547.720 295.600 549.120 ;
        RECT 4.400 545.040 296.000 547.720 ;
        RECT 4.400 543.640 295.600 545.040 ;
        RECT 4.400 540.960 296.000 543.640 ;
        RECT 4.400 539.560 295.600 540.960 ;
        RECT 4.400 536.880 296.000 539.560 ;
        RECT 4.400 535.480 295.600 536.880 ;
        RECT 4.400 532.800 296.000 535.480 ;
        RECT 4.400 531.400 295.600 532.800 ;
        RECT 4.400 528.720 296.000 531.400 ;
        RECT 4.400 527.320 295.600 528.720 ;
        RECT 4.400 524.640 296.000 527.320 ;
        RECT 4.400 523.240 295.600 524.640 ;
        RECT 4.400 520.560 296.000 523.240 ;
        RECT 4.400 519.160 295.600 520.560 ;
        RECT 4.400 516.480 296.000 519.160 ;
        RECT 4.400 515.080 295.600 516.480 ;
        RECT 4.400 512.400 296.000 515.080 ;
        RECT 4.400 511.000 295.600 512.400 ;
        RECT 4.400 508.320 296.000 511.000 ;
        RECT 4.400 506.920 295.600 508.320 ;
        RECT 4.400 504.240 296.000 506.920 ;
        RECT 4.400 502.840 295.600 504.240 ;
        RECT 4.400 500.160 296.000 502.840 ;
        RECT 4.400 498.760 295.600 500.160 ;
        RECT 4.400 496.080 296.000 498.760 ;
        RECT 4.400 494.680 295.600 496.080 ;
        RECT 4.400 492.000 296.000 494.680 ;
        RECT 4.400 490.600 295.600 492.000 ;
        RECT 4.400 487.920 296.000 490.600 ;
        RECT 4.400 486.520 295.600 487.920 ;
        RECT 4.400 483.840 296.000 486.520 ;
        RECT 4.400 482.440 295.600 483.840 ;
        RECT 4.400 479.760 296.000 482.440 ;
        RECT 4.400 478.360 295.600 479.760 ;
        RECT 4.400 475.680 296.000 478.360 ;
        RECT 4.400 474.280 295.600 475.680 ;
        RECT 4.400 471.600 296.000 474.280 ;
        RECT 4.400 470.200 295.600 471.600 ;
        RECT 4.400 467.520 296.000 470.200 ;
        RECT 4.400 466.120 295.600 467.520 ;
        RECT 4.400 463.440 296.000 466.120 ;
        RECT 4.400 462.040 295.600 463.440 ;
        RECT 4.400 459.360 296.000 462.040 ;
        RECT 4.400 457.960 295.600 459.360 ;
        RECT 4.400 455.280 296.000 457.960 ;
        RECT 4.400 453.880 295.600 455.280 ;
        RECT 4.400 451.200 296.000 453.880 ;
        RECT 4.400 449.800 295.600 451.200 ;
        RECT 4.400 447.120 296.000 449.800 ;
        RECT 4.400 445.720 295.600 447.120 ;
        RECT 4.400 443.040 296.000 445.720 ;
        RECT 4.400 441.640 295.600 443.040 ;
        RECT 4.400 438.960 296.000 441.640 ;
        RECT 4.400 437.560 295.600 438.960 ;
        RECT 4.400 434.880 296.000 437.560 ;
        RECT 4.400 433.480 295.600 434.880 ;
        RECT 4.400 430.800 296.000 433.480 ;
        RECT 4.400 429.400 295.600 430.800 ;
        RECT 4.400 426.720 296.000 429.400 ;
        RECT 4.400 425.320 295.600 426.720 ;
        RECT 4.400 422.640 296.000 425.320 ;
        RECT 4.400 421.240 295.600 422.640 ;
        RECT 4.400 418.560 296.000 421.240 ;
        RECT 4.400 417.160 295.600 418.560 ;
        RECT 4.400 414.480 296.000 417.160 ;
        RECT 4.400 413.080 295.600 414.480 ;
        RECT 4.400 410.400 296.000 413.080 ;
        RECT 4.400 409.000 295.600 410.400 ;
        RECT 4.400 406.320 296.000 409.000 ;
        RECT 4.400 404.920 295.600 406.320 ;
        RECT 4.400 402.240 296.000 404.920 ;
        RECT 4.400 400.840 295.600 402.240 ;
        RECT 4.400 398.160 296.000 400.840 ;
        RECT 4.400 396.760 295.600 398.160 ;
        RECT 4.400 394.080 296.000 396.760 ;
        RECT 4.400 392.680 295.600 394.080 ;
        RECT 4.400 390.000 296.000 392.680 ;
        RECT 4.400 388.600 295.600 390.000 ;
        RECT 4.400 385.920 296.000 388.600 ;
        RECT 4.400 384.520 295.600 385.920 ;
        RECT 4.400 381.840 296.000 384.520 ;
        RECT 4.400 380.440 295.600 381.840 ;
        RECT 4.400 377.760 296.000 380.440 ;
        RECT 4.400 376.360 295.600 377.760 ;
        RECT 4.400 373.680 296.000 376.360 ;
        RECT 4.400 372.280 295.600 373.680 ;
        RECT 4.400 369.600 296.000 372.280 ;
        RECT 4.400 368.200 295.600 369.600 ;
        RECT 4.400 365.520 296.000 368.200 ;
        RECT 4.400 364.120 295.600 365.520 ;
        RECT 4.400 361.440 296.000 364.120 ;
        RECT 4.400 360.040 295.600 361.440 ;
        RECT 4.400 357.360 296.000 360.040 ;
        RECT 4.400 355.960 295.600 357.360 ;
        RECT 4.400 353.280 296.000 355.960 ;
        RECT 4.400 351.880 295.600 353.280 ;
        RECT 4.400 349.200 296.000 351.880 ;
        RECT 4.400 347.800 295.600 349.200 ;
        RECT 4.400 345.120 296.000 347.800 ;
        RECT 4.400 343.720 295.600 345.120 ;
        RECT 4.400 341.040 296.000 343.720 ;
        RECT 4.400 339.640 295.600 341.040 ;
        RECT 4.400 336.960 296.000 339.640 ;
        RECT 4.400 335.560 295.600 336.960 ;
        RECT 4.400 332.880 296.000 335.560 ;
        RECT 4.400 331.480 295.600 332.880 ;
        RECT 4.400 328.800 296.000 331.480 ;
        RECT 4.400 327.400 295.600 328.800 ;
        RECT 4.400 324.720 296.000 327.400 ;
        RECT 4.400 323.320 295.600 324.720 ;
        RECT 4.400 320.640 296.000 323.320 ;
        RECT 4.400 319.240 295.600 320.640 ;
        RECT 4.400 316.560 296.000 319.240 ;
        RECT 4.400 315.160 295.600 316.560 ;
        RECT 4.400 312.480 296.000 315.160 ;
        RECT 4.400 311.080 295.600 312.480 ;
        RECT 4.400 308.400 296.000 311.080 ;
        RECT 4.400 307.000 295.600 308.400 ;
        RECT 4.400 304.320 296.000 307.000 ;
        RECT 4.400 302.920 295.600 304.320 ;
        RECT 4.400 300.240 296.000 302.920 ;
        RECT 4.400 298.840 295.600 300.240 ;
        RECT 4.400 296.160 296.000 298.840 ;
        RECT 4.400 294.760 295.600 296.160 ;
        RECT 4.400 292.080 296.000 294.760 ;
        RECT 4.400 290.680 295.600 292.080 ;
        RECT 4.400 288.000 296.000 290.680 ;
        RECT 4.400 286.600 295.600 288.000 ;
        RECT 4.400 283.920 296.000 286.600 ;
        RECT 4.400 282.520 295.600 283.920 ;
        RECT 4.400 279.840 296.000 282.520 ;
        RECT 4.400 278.440 295.600 279.840 ;
        RECT 4.400 275.760 296.000 278.440 ;
        RECT 4.400 274.360 295.600 275.760 ;
        RECT 4.400 271.680 296.000 274.360 ;
        RECT 4.400 270.280 295.600 271.680 ;
        RECT 4.400 267.600 296.000 270.280 ;
        RECT 4.400 266.200 295.600 267.600 ;
        RECT 4.400 263.520 296.000 266.200 ;
        RECT 4.400 262.120 295.600 263.520 ;
        RECT 4.400 259.440 296.000 262.120 ;
        RECT 4.400 258.040 295.600 259.440 ;
        RECT 4.400 255.360 296.000 258.040 ;
        RECT 4.400 253.960 295.600 255.360 ;
        RECT 4.400 251.280 296.000 253.960 ;
        RECT 4.400 249.880 295.600 251.280 ;
        RECT 4.400 247.200 296.000 249.880 ;
        RECT 4.400 245.800 295.600 247.200 ;
        RECT 4.400 243.120 296.000 245.800 ;
        RECT 4.400 241.720 295.600 243.120 ;
        RECT 4.400 239.040 296.000 241.720 ;
        RECT 4.400 237.640 295.600 239.040 ;
        RECT 4.400 234.960 296.000 237.640 ;
        RECT 4.400 233.560 295.600 234.960 ;
        RECT 4.400 230.880 296.000 233.560 ;
        RECT 4.400 229.480 295.600 230.880 ;
        RECT 4.400 226.800 296.000 229.480 ;
        RECT 4.400 225.400 295.600 226.800 ;
        RECT 4.400 222.720 296.000 225.400 ;
        RECT 4.400 221.320 295.600 222.720 ;
        RECT 4.400 218.640 296.000 221.320 ;
        RECT 4.400 217.240 295.600 218.640 ;
        RECT 4.400 214.560 296.000 217.240 ;
        RECT 4.400 213.160 295.600 214.560 ;
        RECT 4.400 210.480 296.000 213.160 ;
        RECT 4.400 209.080 295.600 210.480 ;
        RECT 4.400 206.400 296.000 209.080 ;
        RECT 4.400 205.000 295.600 206.400 ;
        RECT 4.400 202.320 296.000 205.000 ;
        RECT 4.400 200.920 295.600 202.320 ;
        RECT 4.400 198.240 296.000 200.920 ;
        RECT 4.400 196.840 295.600 198.240 ;
        RECT 4.400 194.160 296.000 196.840 ;
        RECT 4.400 192.760 295.600 194.160 ;
        RECT 4.400 190.080 296.000 192.760 ;
        RECT 4.400 188.680 295.600 190.080 ;
        RECT 4.400 186.000 296.000 188.680 ;
        RECT 4.400 184.600 295.600 186.000 ;
        RECT 4.400 181.920 296.000 184.600 ;
        RECT 4.400 180.520 295.600 181.920 ;
        RECT 4.400 177.840 296.000 180.520 ;
        RECT 4.400 176.440 295.600 177.840 ;
        RECT 4.400 173.760 296.000 176.440 ;
        RECT 4.400 172.360 295.600 173.760 ;
        RECT 4.400 169.680 296.000 172.360 ;
        RECT 4.400 168.280 295.600 169.680 ;
        RECT 4.400 165.600 296.000 168.280 ;
        RECT 4.400 164.200 295.600 165.600 ;
        RECT 4.400 161.520 296.000 164.200 ;
        RECT 4.400 160.120 295.600 161.520 ;
        RECT 4.400 157.440 296.000 160.120 ;
        RECT 4.400 156.040 295.600 157.440 ;
        RECT 4.400 153.360 296.000 156.040 ;
        RECT 4.400 151.960 295.600 153.360 ;
        RECT 4.400 149.280 296.000 151.960 ;
        RECT 4.400 147.880 295.600 149.280 ;
        RECT 4.400 145.200 296.000 147.880 ;
        RECT 4.400 143.800 295.600 145.200 ;
        RECT 4.400 141.120 296.000 143.800 ;
        RECT 4.400 139.720 295.600 141.120 ;
        RECT 4.400 137.040 296.000 139.720 ;
        RECT 4.400 135.640 295.600 137.040 ;
        RECT 4.400 132.960 296.000 135.640 ;
        RECT 4.400 131.560 295.600 132.960 ;
        RECT 4.400 128.880 296.000 131.560 ;
        RECT 4.400 127.480 295.600 128.880 ;
        RECT 4.400 124.800 296.000 127.480 ;
        RECT 4.400 123.400 295.600 124.800 ;
        RECT 4.400 120.720 296.000 123.400 ;
        RECT 4.400 119.320 295.600 120.720 ;
        RECT 4.400 116.640 296.000 119.320 ;
        RECT 4.400 115.240 295.600 116.640 ;
        RECT 4.400 112.560 296.000 115.240 ;
        RECT 4.400 111.160 295.600 112.560 ;
        RECT 3.030 108.480 296.000 111.160 ;
        RECT 3.030 107.080 295.600 108.480 ;
        RECT 3.030 104.400 296.000 107.080 ;
        RECT 3.030 103.000 295.600 104.400 ;
        RECT 3.030 100.320 296.000 103.000 ;
        RECT 3.030 98.920 295.600 100.320 ;
        RECT 3.030 96.240 296.000 98.920 ;
        RECT 3.030 94.840 295.600 96.240 ;
        RECT 3.030 92.160 296.000 94.840 ;
        RECT 3.030 90.760 295.600 92.160 ;
        RECT 3.030 88.080 296.000 90.760 ;
        RECT 3.030 86.680 295.600 88.080 ;
        RECT 3.030 84.000 296.000 86.680 ;
        RECT 3.030 82.600 295.600 84.000 ;
        RECT 3.030 79.920 296.000 82.600 ;
        RECT 3.030 78.520 295.600 79.920 ;
        RECT 3.030 75.840 296.000 78.520 ;
        RECT 3.030 74.440 295.600 75.840 ;
        RECT 3.030 71.760 296.000 74.440 ;
        RECT 3.030 70.360 295.600 71.760 ;
        RECT 3.030 67.680 296.000 70.360 ;
        RECT 3.030 66.280 295.600 67.680 ;
        RECT 3.030 63.600 296.000 66.280 ;
        RECT 3.030 62.200 295.600 63.600 ;
        RECT 3.030 59.520 296.000 62.200 ;
        RECT 3.030 58.120 295.600 59.520 ;
        RECT 3.030 55.440 296.000 58.120 ;
        RECT 3.030 54.040 295.600 55.440 ;
        RECT 3.030 51.360 296.000 54.040 ;
        RECT 3.030 49.960 295.600 51.360 ;
        RECT 3.030 47.280 296.000 49.960 ;
        RECT 3.030 45.880 295.600 47.280 ;
        RECT 3.030 43.200 296.000 45.880 ;
        RECT 3.030 41.800 295.600 43.200 ;
        RECT 3.030 39.120 296.000 41.800 ;
        RECT 3.030 37.720 295.600 39.120 ;
        RECT 3.030 35.040 296.000 37.720 ;
        RECT 3.030 33.640 295.600 35.040 ;
        RECT 3.030 30.960 296.000 33.640 ;
        RECT 3.030 29.560 295.600 30.960 ;
        RECT 3.030 26.880 296.000 29.560 ;
        RECT 3.030 25.480 295.600 26.880 ;
        RECT 3.030 22.800 296.000 25.480 ;
        RECT 3.030 21.400 295.600 22.800 ;
        RECT 3.030 10.715 296.000 21.400 ;
      LAYER met4 ;
        RECT 0.310 11.735 20.640 787.265 ;
        RECT 23.040 11.735 97.440 787.265 ;
        RECT 99.840 11.735 174.240 787.265 ;
        RECT 176.640 11.735 251.040 787.265 ;
        RECT 253.440 11.735 287.665 787.265 ;
  END
END interconnect_inner
END LIBRARY

