magic
tech gf180mcuD
magscale 1 10
timestamp 1700096716
<< metal1 >>
rect 252242 305454 252254 305506
rect 252306 305503 252318 305506
rect 253026 305503 253038 305506
rect 252306 305457 253038 305503
rect 252306 305454 252318 305457
rect 253026 305454 253038 305457
rect 253090 305454 253102 305506
rect 185826 12910 185838 12962
rect 185890 12959 185902 12962
rect 186498 12959 186510 12962
rect 185890 12913 186510 12959
rect 185890 12910 185902 12913
rect 186498 12910 186510 12913
rect 186562 12910 186574 12962
<< via1 >>
rect 252254 305454 252306 305506
rect 253038 305454 253090 305506
rect 185838 12910 185890 12962
rect 186510 12910 186562 12962
<< metal2 >>
rect 11032 595672 11256 597000
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11004 595560 11256 595672
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 99260 595560 99512 595672
rect 121324 595560 121576 595672
rect 143388 595560 143640 595672
rect 165452 595560 165704 595672
rect 187516 595560 187768 595672
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 364056 595560 364308 595672
rect 4844 416724 4900 416734
rect 4844 394436 4900 416668
rect 4844 394370 4900 394380
rect 4956 403284 5012 403294
rect 4956 377188 5012 403228
rect 11004 378868 11060 595560
rect 19180 590996 19236 591006
rect 19180 380548 19236 590940
rect 33068 590996 33124 595560
rect 33068 590930 33124 590940
rect 55132 590884 55188 595560
rect 55132 590818 55188 590828
rect 77308 590772 77364 595560
rect 77308 590706 77364 590716
rect 99260 590660 99316 595560
rect 99260 590594 99316 590604
rect 121324 577332 121380 595560
rect 143388 590548 143444 595560
rect 143388 590482 143444 590492
rect 121324 577266 121380 577276
rect 162092 590212 162148 590222
rect 29260 577220 29316 577230
rect 28476 577108 28532 577118
rect 28476 574532 28532 577052
rect 29260 575092 29316 577164
rect 162092 576100 162148 590156
rect 165452 590212 165508 595560
rect 165452 590146 165508 590156
rect 162092 576034 162148 576044
rect 169708 577332 169764 577342
rect 169708 575988 169764 577276
rect 187516 577332 187572 595560
rect 193228 583828 193284 583838
rect 187516 577266 187572 577276
rect 188076 579348 188132 579358
rect 169708 575922 169764 575932
rect 188076 575876 188132 579292
rect 193228 579348 193284 583772
rect 209580 583828 209636 595560
rect 209580 583762 209636 583772
rect 225932 590212 225988 590222
rect 193228 579282 193284 579292
rect 225932 576324 225988 590156
rect 231644 590212 231700 595560
rect 231644 590146 231700 590156
rect 242732 590548 242788 590558
rect 225932 576258 225988 576268
rect 188076 575810 188132 575820
rect 242732 575652 242788 590492
rect 253708 590548 253764 595560
rect 253708 590482 253764 590492
rect 242732 575586 242788 575596
rect 268716 583044 268772 583054
rect 268716 575540 268772 582988
rect 275772 583044 275828 595560
rect 275772 582978 275828 582988
rect 295596 587972 295652 587982
rect 268716 575474 268772 575484
rect 292236 581364 292292 581374
rect 292236 575428 292292 581308
rect 295596 581364 295652 587916
rect 297836 587972 297892 595560
rect 317548 590212 317604 590222
rect 297836 587906 297892 587916
rect 314188 587972 314244 587982
rect 314188 584724 314244 587916
rect 317548 587972 317604 590156
rect 319900 590212 319956 595560
rect 319900 590146 319956 590156
rect 336812 590548 336868 590558
rect 317548 587906 317604 587916
rect 295596 581298 295652 581308
rect 314076 584668 314244 584724
rect 310828 579572 310884 579582
rect 310828 577220 310884 579516
rect 314076 579572 314132 584668
rect 314076 579506 314132 579516
rect 310828 577154 310884 577164
rect 336812 577108 336868 590492
rect 341964 590548 342020 595560
rect 341964 590482 342020 590492
rect 364252 590548 364308 595560
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 430248 595560 430500 595672
rect 452312 595560 452564 595672
rect 474376 595560 474628 595672
rect 496440 595560 496692 595672
rect 518504 595560 518756 595672
rect 540568 595560 540820 595672
rect 364252 590482 364308 590492
rect 380492 590548 380548 590558
rect 380492 577892 380548 590492
rect 386092 581364 386148 595560
rect 386092 581298 386148 581308
rect 394828 581364 394884 581374
rect 380492 577826 380548 577836
rect 383068 577892 383124 577902
rect 336812 577042 336868 577052
rect 292236 575362 292292 575372
rect 383068 575428 383124 577836
rect 394828 575540 394884 581308
rect 408268 575652 408324 595560
rect 430444 590548 430500 595560
rect 452508 590660 452564 595560
rect 474572 590772 474628 595560
rect 496636 590884 496692 595560
rect 518700 590996 518756 595560
rect 540764 591108 540820 595560
rect 540764 591042 540820 591052
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 518700 590930 518756 590940
rect 496636 590818 496692 590828
rect 474572 590706 474628 590716
rect 452508 590594 452564 590604
rect 430444 590482 430500 590492
rect 408268 575586 408324 575596
rect 394828 575474 394884 575484
rect 383068 575362 383124 575372
rect 29260 575026 29316 575036
rect 28476 574466 28532 574476
rect 19180 380482 19236 380492
rect 27692 389732 27748 389742
rect 11004 378802 11060 378812
rect 27692 377972 27748 389676
rect 27916 378980 27972 395080
rect 30268 394548 30324 394558
rect 30156 393204 30212 393214
rect 28476 393092 28532 393102
rect 28476 389844 28532 393036
rect 30156 391412 30212 393148
rect 30268 392532 30324 394492
rect 30268 392466 30324 392476
rect 31948 392308 32004 395080
rect 35980 392420 36036 395080
rect 35980 392354 36036 392364
rect 37772 392532 37828 392542
rect 31948 392242 32004 392252
rect 30156 391356 30324 391412
rect 28476 389778 28532 389788
rect 28588 389732 28644 389742
rect 28588 384804 28644 389676
rect 30268 389396 30324 391356
rect 30268 389330 30324 389340
rect 31052 389732 31108 389742
rect 28588 384738 28644 384748
rect 31052 384132 31108 389676
rect 35084 389732 35140 389742
rect 34412 389396 34468 389406
rect 31052 384066 31108 384076
rect 33404 384692 33460 384702
rect 33404 381892 33460 384636
rect 33404 381826 33460 381836
rect 33516 383012 33572 383022
rect 33516 379764 33572 382956
rect 34412 381444 34468 389340
rect 35084 387940 35140 389676
rect 37772 389732 37828 392476
rect 37772 389666 37828 389676
rect 35084 387874 35140 387884
rect 35196 389508 35252 389518
rect 35196 386372 35252 389452
rect 40012 387268 40068 395080
rect 40236 389732 40292 389742
rect 40236 388052 40292 389676
rect 40236 387996 40404 388052
rect 40012 387202 40068 387212
rect 35196 386306 35252 386316
rect 39004 386372 39060 386382
rect 34412 381378 34468 381388
rect 36764 384132 36820 384142
rect 33516 379698 33572 379708
rect 27916 378914 27972 378924
rect 27692 377906 27748 377916
rect 28700 377972 28756 377982
rect 36764 377972 36820 384076
rect 37772 381892 37828 381902
rect 36876 381444 36932 381454
rect 36876 379540 36932 381388
rect 36876 379474 36932 379484
rect 36764 377916 37044 377972
rect 4956 377122 5012 377132
rect 28700 375732 28756 377916
rect 36876 377412 36932 377422
rect 36876 375956 36932 377356
rect 36876 375890 36932 375900
rect 28700 375666 28756 375676
rect 36988 374276 37044 377916
rect 37772 375844 37828 381836
rect 39004 381444 39060 386316
rect 40348 385588 40404 387996
rect 40348 385522 40404 385532
rect 41132 387940 41188 387950
rect 41132 382228 41188 387884
rect 44044 387380 44100 395080
rect 44044 387314 44100 387324
rect 41132 382162 41188 382172
rect 47852 385588 47908 385598
rect 39004 381378 39060 381388
rect 42812 381444 42868 381454
rect 42028 379540 42084 379550
rect 42028 377412 42084 379484
rect 42028 377346 42084 377356
rect 37772 375778 37828 375788
rect 36988 374210 37044 374220
rect 42812 372484 42868 381388
rect 46956 379316 47012 379326
rect 46956 376292 47012 379260
rect 46956 376226 47012 376236
rect 47852 376180 47908 385532
rect 48076 384132 48132 395080
rect 52108 392644 52164 395080
rect 52108 392578 52164 392588
rect 56140 392532 56196 395080
rect 56140 392466 56196 392476
rect 57036 392420 57092 392430
rect 57036 390852 57092 392364
rect 60172 392420 60228 395080
rect 60172 392354 60228 392364
rect 63868 392644 63924 392654
rect 57036 390786 57092 390796
rect 60396 392308 60452 392318
rect 60396 388948 60452 392252
rect 63868 390964 63924 392588
rect 64204 391524 64260 395080
rect 64204 391458 64260 391468
rect 65660 391524 65716 391534
rect 63868 390898 63924 390908
rect 60396 388882 60452 388892
rect 65660 385588 65716 391468
rect 68236 385700 68292 395080
rect 70476 392532 70532 392542
rect 70476 387492 70532 392476
rect 72268 392308 72324 395080
rect 72268 392242 72324 392252
rect 70476 387426 70532 387436
rect 76300 385812 76356 395080
rect 80332 389060 80388 395080
rect 80332 388994 80388 389004
rect 84364 387604 84420 395080
rect 88396 387716 88452 395080
rect 88396 387650 88452 387660
rect 84364 387538 84420 387548
rect 76300 385746 76356 385756
rect 68236 385634 68292 385644
rect 65660 385522 65716 385532
rect 92428 384244 92484 395080
rect 96460 393092 96516 395080
rect 96460 393026 96516 393036
rect 100492 392532 100548 395080
rect 100492 392466 100548 392476
rect 104524 385924 104580 395080
rect 108556 386036 108612 395080
rect 112588 391076 112644 395080
rect 112588 391010 112644 391020
rect 116620 389172 116676 395080
rect 120652 389284 120708 395080
rect 120652 389218 120708 389228
rect 116620 389106 116676 389116
rect 108556 385970 108612 385980
rect 104524 385858 104580 385868
rect 124684 384356 124740 395080
rect 128716 392980 128772 395080
rect 128716 392914 128772 392924
rect 132748 391524 132804 395080
rect 136780 392756 136836 395080
rect 136780 392690 136836 392700
rect 140812 392644 140868 395080
rect 140812 392578 140868 392588
rect 132748 391458 132804 391468
rect 136108 391524 136164 391534
rect 136108 386148 136164 391468
rect 144844 391188 144900 395080
rect 144844 391122 144900 391132
rect 148876 387828 148932 395080
rect 148876 387762 148932 387772
rect 152236 394436 152292 394446
rect 136108 386082 136164 386092
rect 124684 384290 124740 384300
rect 92428 384178 92484 384188
rect 48076 384066 48132 384076
rect 48636 382228 48692 382238
rect 48636 381332 48692 382172
rect 48636 381266 48692 381276
rect 50428 381332 50484 381342
rect 50428 378084 50484 381276
rect 50428 378018 50484 378028
rect 57036 377972 57092 377982
rect 47852 376114 47908 376124
rect 48636 377412 48692 377422
rect 48636 374388 48692 377356
rect 48636 374322 48692 374332
rect 50428 376292 50484 376302
rect 50428 373044 50484 376236
rect 57036 376068 57092 377916
rect 57036 376002 57092 376012
rect 62188 376180 62244 376190
rect 62188 374500 62244 376124
rect 62188 374434 62244 374444
rect 151004 375956 151060 375966
rect 149324 374388 149380 374398
rect 149324 374164 149380 374332
rect 151004 374388 151060 375900
rect 151004 374322 151060 374332
rect 151116 374500 151172 374510
rect 149324 374108 149604 374164
rect 50428 372978 50484 372988
rect 42812 372418 42868 372428
rect 149548 370692 149604 374108
rect 151116 372988 151172 374444
rect 151116 372932 151284 372988
rect 149548 370626 149604 370636
rect 151116 372596 151172 372606
rect 151116 366212 151172 372540
rect 151228 369684 151284 372932
rect 151228 369618 151284 369628
rect 151452 370692 151508 370702
rect 151452 368004 151508 370636
rect 151452 367938 151508 367948
rect 151116 366156 151284 366212
rect 151228 364532 151284 366156
rect 151228 364466 151284 364476
rect 152236 58884 152292 394380
rect 152908 391300 152964 395080
rect 156940 394324 156996 395080
rect 156940 394258 156996 394268
rect 160972 392868 161028 395080
rect 160972 392802 161028 392812
rect 152908 391234 152964 391244
rect 164556 392420 164612 392430
rect 164556 390740 164612 392364
rect 165004 391636 165060 395080
rect 165004 391570 165060 391580
rect 164556 390674 164612 390684
rect 169036 390628 169092 395080
rect 169036 390562 169092 390572
rect 173068 387940 173124 395080
rect 173068 387874 173124 387884
rect 176316 391636 176372 391646
rect 176316 386260 176372 391580
rect 177100 389396 177156 395080
rect 181160 395052 181412 395108
rect 181356 391524 181412 395052
rect 185164 392420 185220 395080
rect 185164 392354 185220 392364
rect 186396 392980 186452 392990
rect 181356 391468 181524 391524
rect 177100 389330 177156 389340
rect 180124 390852 180180 390862
rect 176316 386194 176372 386204
rect 180124 381864 180180 390796
rect 181468 387156 181524 391468
rect 186396 391412 186452 392924
rect 186396 391346 186452 391356
rect 188972 392308 189028 392318
rect 187292 390964 187348 390974
rect 183708 387380 183764 387390
rect 181468 387090 181524 387100
rect 181916 387268 181972 387278
rect 181916 381864 181972 387212
rect 183708 381864 183764 387324
rect 185500 384132 185556 384142
rect 185500 381864 185556 384076
rect 187292 381864 187348 390908
rect 188972 390404 189028 392252
rect 189196 392308 189252 395080
rect 189196 392242 189252 392252
rect 188972 390338 189028 390348
rect 192668 390740 192724 390750
rect 189084 388948 189140 388958
rect 189084 381864 189140 388892
rect 190876 387492 190932 387502
rect 190876 381864 190932 387436
rect 192668 381864 192724 390684
rect 193228 390740 193284 395080
rect 193228 390674 193284 390684
rect 194908 392532 194964 392542
rect 194908 386372 194964 392476
rect 197260 388948 197316 395080
rect 197260 388882 197316 388892
rect 198044 390404 198100 390414
rect 194908 386306 194964 386316
rect 196252 385700 196308 385710
rect 194460 385588 194516 385598
rect 194460 381864 194516 385532
rect 196252 381864 196308 385644
rect 198044 381864 198100 390348
rect 201292 387380 201348 395080
rect 201292 387314 201348 387324
rect 201628 389060 201684 389070
rect 199836 385812 199892 385822
rect 199836 381864 199892 385756
rect 201628 381864 201684 389004
rect 205212 387716 205268 387726
rect 203420 387604 203476 387614
rect 203420 381864 203476 387548
rect 205212 381864 205268 387660
rect 205324 385588 205380 395080
rect 209384 395052 209972 395108
rect 205324 385522 205380 385532
rect 208796 393204 208852 393214
rect 207004 384244 207060 384254
rect 207004 381864 207060 384188
rect 208796 381864 208852 393148
rect 209916 391524 209972 395052
rect 209916 391468 210084 391524
rect 210028 385700 210084 391468
rect 210028 385634 210084 385644
rect 210588 386372 210644 386382
rect 210588 381864 210644 386316
rect 212380 385924 212436 385934
rect 212380 381864 212436 385868
rect 213388 385812 213444 395080
rect 215964 391076 216020 391086
rect 213388 385746 213444 385756
rect 214172 386036 214228 386046
rect 214172 381864 214228 385980
rect 215964 381864 216020 391020
rect 217420 387492 217476 395080
rect 221452 390852 221508 395080
rect 223468 392756 223524 392766
rect 221452 390786 221508 390796
rect 223132 391412 223188 391422
rect 219548 389284 219604 389294
rect 217420 387426 217476 387436
rect 217756 389172 217812 389182
rect 217756 381864 217812 389116
rect 219548 381864 219604 389228
rect 221340 384356 221396 384366
rect 221340 381864 221396 384300
rect 223132 381864 223188 391356
rect 223468 386372 223524 392700
rect 225484 391524 225540 395080
rect 229516 392756 229572 395080
rect 229516 392690 229572 392700
rect 225484 391458 225540 391468
rect 228508 392644 228564 392654
rect 223468 386306 223524 386316
rect 226716 386372 226772 386382
rect 224924 386148 224980 386158
rect 224924 381864 224980 386092
rect 226716 381864 226772 386316
rect 228508 381864 228564 392588
rect 233548 392532 233604 395080
rect 233548 392466 233604 392476
rect 235676 394324 235732 394334
rect 233884 391300 233940 391310
rect 230300 391188 230356 391198
rect 230300 381864 230356 391132
rect 232092 387828 232148 387838
rect 232092 381864 232148 387772
rect 233884 381864 233940 391244
rect 235676 381864 235732 394268
rect 237468 392868 237524 392878
rect 237468 381864 237524 392812
rect 237580 392644 237636 395080
rect 237580 392578 237636 392588
rect 238588 392756 238644 392766
rect 238588 389060 238644 392700
rect 238588 388994 238644 389004
rect 241052 390628 241108 390638
rect 239260 386260 239316 386270
rect 239260 381864 239316 386204
rect 241052 381864 241108 390572
rect 241612 390628 241668 395080
rect 241612 390562 241668 390572
rect 241948 392420 242004 392430
rect 241948 385924 242004 392364
rect 245644 392420 245700 395080
rect 245644 392354 245700 392364
rect 246988 392308 247044 392318
rect 244636 389396 244692 389406
rect 241948 385858 242004 385868
rect 242844 387940 242900 387950
rect 242844 381864 242900 387884
rect 244636 381864 244692 389340
rect 246428 387268 246484 387278
rect 246428 381864 246484 387212
rect 246988 386372 247044 392252
rect 249676 392308 249732 395080
rect 249676 392242 249732 392252
rect 251804 390740 251860 390750
rect 246988 386306 247044 386316
rect 250012 386372 250068 386382
rect 248220 385924 248276 385934
rect 248220 381864 248276 385868
rect 250012 381864 250068 386316
rect 251804 381864 251860 390684
rect 253708 389172 253764 395080
rect 253708 389106 253764 389116
rect 253596 388948 253652 388958
rect 253596 381864 253652 388892
rect 257740 388948 257796 395080
rect 257740 388882 257796 388892
rect 260316 392644 260372 392654
rect 255388 387380 255444 387390
rect 255388 381864 255444 387324
rect 260316 385924 260372 392588
rect 261772 389284 261828 395080
rect 263788 392532 263844 392542
rect 263788 390740 263844 392476
rect 265468 392420 265524 392430
rect 263788 390674 263844 390684
rect 264348 390852 264404 390862
rect 261772 389218 261828 389228
rect 260316 385858 260372 385868
rect 262556 387492 262612 387502
rect 260764 385812 260820 385822
rect 258972 385700 259028 385710
rect 257180 385588 257236 385598
rect 257180 381864 257236 385532
rect 258972 381864 259028 385644
rect 260764 381864 260820 385756
rect 262556 381864 262612 387436
rect 264348 381864 264404 390796
rect 265468 387268 265524 392364
rect 265468 387202 265524 387212
rect 265804 385588 265860 395080
rect 265804 385522 265860 385532
rect 266140 390964 266196 390974
rect 266140 381864 266196 390908
rect 269724 390740 269780 390750
rect 267932 389060 267988 389070
rect 267932 381864 267988 389004
rect 269724 381864 269780 390684
rect 269836 385700 269892 395080
rect 270396 392308 270452 392318
rect 270396 388052 270452 392252
rect 273868 392308 273924 395080
rect 273868 392242 273924 392252
rect 270396 387986 270452 387996
rect 273308 390628 273364 390638
rect 269836 385634 269892 385644
rect 271516 385924 271572 385934
rect 271516 381864 271572 385868
rect 273308 381864 273364 390572
rect 276892 388052 276948 388062
rect 275100 387268 275156 387278
rect 275100 381864 275156 387212
rect 276892 381864 276948 387996
rect 277900 385812 277956 395080
rect 277900 385746 277956 385756
rect 278684 389172 278740 389182
rect 278684 381864 278740 389116
rect 280476 388948 280532 388958
rect 280476 381864 280532 388892
rect 281932 387268 281988 395080
rect 281932 387202 281988 387212
rect 282268 389284 282324 389294
rect 282268 381864 282324 389228
rect 285964 386484 286020 395080
rect 285964 386418 286020 386428
rect 287644 392308 287700 392318
rect 285852 385700 285908 385710
rect 284060 385588 284116 385598
rect 284060 381864 284116 385532
rect 285852 381864 285908 385644
rect 287644 381864 287700 392252
rect 289996 392308 290052 395080
rect 289996 392242 290052 392252
rect 291228 387268 291284 387278
rect 289436 385812 289492 385822
rect 289436 381864 289492 385756
rect 291228 381864 291284 387212
rect 293020 386484 293076 386494
rect 293020 381864 293076 386428
rect 294028 386372 294084 395080
rect 294028 386306 294084 386316
rect 294812 392308 294868 392318
rect 294812 381864 294868 392252
rect 296604 386372 296660 386382
rect 296604 381864 296660 386316
rect 298060 381892 298116 395080
rect 301980 390740 302036 390750
rect 300188 388052 300244 388062
rect 298060 381836 298424 381892
rect 300188 381864 300244 387996
rect 301980 381864 302036 390684
rect 302092 388052 302148 395080
rect 306124 390740 306180 395080
rect 306124 390674 306180 390684
rect 305564 390628 305620 390638
rect 302092 387986 302148 387996
rect 303772 389732 303828 389742
rect 303772 381864 303828 389676
rect 305564 381864 305620 390572
rect 310156 389732 310212 395080
rect 310156 389666 310212 389676
rect 310940 392756 310996 392766
rect 309148 385700 309204 385710
rect 307356 385588 307412 385598
rect 307356 381864 307412 385532
rect 309148 381864 309204 385644
rect 310940 381864 310996 392700
rect 312732 392420 312788 392430
rect 312732 381864 312788 392364
rect 314188 390628 314244 395080
rect 314188 390562 314244 390572
rect 314524 392532 314580 392542
rect 314524 381864 314580 392476
rect 318108 392308 318164 392318
rect 316316 387268 316372 387278
rect 316316 381864 316372 387212
rect 318108 381864 318164 392252
rect 318220 385588 318276 395080
rect 321692 390628 321748 390638
rect 318220 385522 318276 385532
rect 319900 385588 319956 385598
rect 319900 381864 319956 385532
rect 321692 381864 321748 390572
rect 322252 385700 322308 395080
rect 326284 392756 326340 395080
rect 326284 392690 326340 392700
rect 325276 392644 325332 392654
rect 322252 385634 322308 385644
rect 323484 387380 323540 387390
rect 323484 381864 323540 387324
rect 325276 381864 325332 392588
rect 330316 392420 330372 395080
rect 334348 392532 334404 395080
rect 334348 392466 334404 392476
rect 334460 392756 334516 392766
rect 330316 392354 330372 392364
rect 334236 392420 334292 392430
rect 332444 389060 332500 389070
rect 328860 387492 328916 387502
rect 327068 386372 327124 386382
rect 327068 381864 327124 386316
rect 328860 381864 328916 387436
rect 330652 385700 330708 385710
rect 330652 381864 330708 385644
rect 332444 381864 332500 389004
rect 334236 381864 334292 392364
rect 334460 387380 334516 392700
rect 334460 387314 334516 387324
rect 336028 390964 336084 390974
rect 336028 386372 336084 390908
rect 336028 386306 336084 386316
rect 337820 390852 337876 390862
rect 336028 385924 336084 385934
rect 336028 381864 336084 385868
rect 337820 381864 337876 390796
rect 338380 387268 338436 395080
rect 342412 392308 342468 395080
rect 342412 392242 342468 392252
rect 343532 392532 343588 392542
rect 338380 387202 338436 387212
rect 340956 388276 341012 388286
rect 339612 386036 339668 386046
rect 339612 381864 339668 385980
rect 340956 385588 341012 388220
rect 340956 385522 341012 385532
rect 341404 387268 341460 387278
rect 341404 381864 341460 387212
rect 343532 385924 343588 392476
rect 346444 388276 346500 395080
rect 346444 388210 346500 388220
rect 348572 391300 348628 391310
rect 344540 387380 344596 387390
rect 344540 386036 344596 387324
rect 344540 385970 344596 385980
rect 344988 386036 345044 386046
rect 343532 385858 343588 385868
rect 343196 385812 343252 385822
rect 343196 381864 343252 385756
rect 344988 381864 345044 385980
rect 346780 385588 346836 385598
rect 346780 381864 346836 385532
rect 348572 381864 348628 391244
rect 350476 390628 350532 395080
rect 354508 392756 354564 395080
rect 354508 392690 354564 392700
rect 358540 392644 358596 395080
rect 358540 392578 358596 392588
rect 359548 392644 359604 392654
rect 355292 392308 355348 392318
rect 350476 390562 350532 390572
rect 351820 390628 351876 390638
rect 351036 389172 351092 389182
rect 350364 386372 350420 386382
rect 350364 381864 350420 386316
rect 351036 385700 351092 389116
rect 351820 386372 351876 390572
rect 351820 386306 351876 386316
rect 352828 388948 352884 388958
rect 351036 385634 351092 385644
rect 352828 384748 352884 388892
rect 355292 386036 355348 392252
rect 359324 390740 359380 390750
rect 355292 385970 355348 385980
rect 355740 386372 355796 386382
rect 352156 384692 352884 384748
rect 353948 385924 354004 385934
rect 352156 381864 352212 384692
rect 353948 381864 354004 385868
rect 355740 381864 355796 386316
rect 357532 385700 357588 385710
rect 357532 381864 357588 385644
rect 359324 381864 359380 390684
rect 359548 386372 359604 392588
rect 362572 390964 362628 395080
rect 362572 390898 362628 390908
rect 362796 391076 362852 391086
rect 359548 386306 359604 386316
rect 361116 384804 361172 384814
rect 361116 381864 361172 384748
rect 362796 384804 362852 391020
rect 366156 387940 366212 387950
rect 362796 384738 362852 384748
rect 362908 386260 362964 386270
rect 362908 381864 362964 386204
rect 366156 385812 366212 387884
rect 366604 387492 366660 395080
rect 366604 387426 366660 387436
rect 367948 391188 368004 391198
rect 366156 385746 366212 385756
rect 366492 386372 366548 386382
rect 364700 384244 364756 384254
rect 364700 381864 364756 384188
rect 366492 381864 366548 386316
rect 367948 386260 368004 391132
rect 370076 389620 370132 389630
rect 367948 386194 368004 386204
rect 368284 386260 368340 386270
rect 368284 381864 368340 386204
rect 370076 381864 370132 389564
rect 370636 389172 370692 395080
rect 370636 389106 370692 389116
rect 371868 389508 371924 389518
rect 371868 381864 371924 389452
rect 374668 389060 374724 395080
rect 378700 392420 378756 395080
rect 378700 392354 378756 392364
rect 381388 393092 381444 393102
rect 374668 388994 374724 389004
rect 378700 392196 378756 392206
rect 374556 387716 374612 387726
rect 374556 385924 374612 387660
rect 374556 385858 374612 385868
rect 377244 386148 377300 386158
rect 373660 384132 373716 384142
rect 373660 381864 373716 384076
rect 375452 384020 375508 384030
rect 375452 381864 375508 383964
rect 377244 381864 377300 386092
rect 378700 386148 378756 392140
rect 380828 390964 380884 390974
rect 378700 386082 378756 386092
rect 379036 386148 379092 386158
rect 379036 381864 379092 386092
rect 380828 381864 380884 390908
rect 381388 386148 381444 393036
rect 382732 392532 382788 395080
rect 382732 392466 382788 392476
rect 386764 390852 386820 395080
rect 386764 390786 386820 390796
rect 387996 389284 388052 389294
rect 381388 386082 381444 386092
rect 384412 387604 384468 387614
rect 382620 386036 382676 386046
rect 382620 381864 382676 385980
rect 384412 381864 384468 387548
rect 386204 385924 386260 385934
rect 386204 381864 386260 385868
rect 387996 381864 388052 389228
rect 390572 387828 390628 387838
rect 389788 385812 389844 385822
rect 389788 381864 389844 385756
rect 390572 385700 390628 387772
rect 390796 387380 390852 395080
rect 393372 392532 393428 392542
rect 390796 387314 390852 387324
rect 391580 387492 391636 387502
rect 390572 385634 390628 385644
rect 391580 381864 391636 387436
rect 393372 381864 393428 392476
rect 394828 387268 394884 395080
rect 396956 392420 397012 392430
rect 394828 387202 394884 387212
rect 395164 387380 395220 387390
rect 395164 381864 395220 387324
rect 396956 381864 397012 392364
rect 398748 390852 398804 390862
rect 398748 381864 398804 390796
rect 398860 387940 398916 395080
rect 402892 392308 402948 395080
rect 402892 392242 402948 392252
rect 404124 392308 404180 392318
rect 398860 387874 398916 387884
rect 401436 391524 401492 391534
rect 400540 385700 400596 385710
rect 400540 381864 400596 385644
rect 401436 385588 401492 391468
rect 401436 385522 401492 385532
rect 402332 389172 402388 389182
rect 402332 381864 402388 389116
rect 404124 381864 404180 392252
rect 406924 391524 406980 395080
rect 406924 391458 406980 391468
rect 407708 391412 407764 391422
rect 405916 387268 405972 387278
rect 405916 381864 405972 387212
rect 407708 381864 407764 391356
rect 410956 391300 411012 395080
rect 410956 391234 411012 391244
rect 414988 390628 415044 395080
rect 414988 390562 415044 390572
rect 419020 388948 419076 395080
rect 419020 388882 419076 388892
rect 423052 387716 423108 395080
rect 423052 387650 423108 387660
rect 424172 393988 424228 393998
rect 163772 380548 163828 380558
rect 154588 376068 154644 376078
rect 152908 375844 152964 375854
rect 152908 373044 152964 375788
rect 152908 372978 152964 372988
rect 154252 375732 154308 375742
rect 152796 372484 152852 372494
rect 152796 369572 152852 372428
rect 154252 371364 154308 375676
rect 154588 374500 154644 376012
rect 154588 374434 154644 374444
rect 157948 374500 158004 374510
rect 154364 374388 154420 374398
rect 154364 371476 154420 374332
rect 156156 374276 156212 374286
rect 156156 372988 156212 374220
rect 156156 372932 156436 372988
rect 154364 371420 154756 371476
rect 154252 371308 154644 371364
rect 153020 369684 153076 369694
rect 152796 369516 152964 369572
rect 152908 364420 152964 369516
rect 152908 364354 152964 364364
rect 153020 363076 153076 369628
rect 154588 368004 154644 371308
rect 154700 369236 154756 371420
rect 156380 369684 156436 372932
rect 157948 371364 158004 374444
rect 157948 371298 158004 371308
rect 159516 372932 159572 372942
rect 159516 371252 159572 372876
rect 159516 371196 159684 371252
rect 156380 369618 156436 369628
rect 154812 369236 154868 369246
rect 154700 369180 154812 369236
rect 154812 369170 154868 369180
rect 159516 369236 159572 369246
rect 154700 368004 154756 368014
rect 154588 367948 154700 368004
rect 154700 367938 154756 367948
rect 157052 368004 157108 368014
rect 153020 363010 153076 363020
rect 154476 364532 154532 364542
rect 154476 361228 154532 364476
rect 154588 364420 154644 364430
rect 154588 362740 154644 364364
rect 154588 362674 154644 362684
rect 154476 361172 154756 361228
rect 154700 354564 154756 361172
rect 154700 354498 154756 354508
rect 157052 352772 157108 367948
rect 159516 367892 159572 369180
rect 159628 368900 159684 371196
rect 162876 371140 162932 371150
rect 159628 368834 159684 368844
rect 160524 369572 160580 369582
rect 160412 367892 160468 367902
rect 159516 367836 159684 367892
rect 159628 365428 159684 367836
rect 159628 365362 159684 365372
rect 158060 362740 158116 362750
rect 158060 358820 158116 362684
rect 158060 358754 158116 358764
rect 157052 352706 157108 352716
rect 158844 354452 158900 354462
rect 158844 347844 158900 354396
rect 158844 347778 158900 347788
rect 160412 230244 160468 367836
rect 160524 257124 160580 369516
rect 162876 364532 162932 371084
rect 162876 364466 162932 364476
rect 162092 363076 162148 363086
rect 160860 352772 160916 352782
rect 160860 348740 160916 352716
rect 160860 348674 160916 348684
rect 160524 257058 160580 257068
rect 160412 230178 160468 230188
rect 152236 58818 152292 58828
rect 153692 79044 153748 79054
rect 150332 40068 150388 40078
rect 4172 36932 4228 36942
rect 3500 23492 3556 23502
rect 3500 17668 3556 23436
rect 3500 17602 3556 17612
rect 4172 16772 4228 36876
rect 150332 17668 150388 40012
rect 153692 32004 153748 78988
rect 162092 66052 162148 363020
rect 162204 358820 162260 358830
rect 162204 69636 162260 358764
rect 162204 69570 162260 69580
rect 162316 347732 162372 347742
rect 162316 66948 162372 347676
rect 162428 257124 162484 257134
rect 162428 67844 162484 257068
rect 162652 230244 162708 230254
rect 162652 68740 162708 230188
rect 162652 68674 162708 68684
rect 162428 67778 162484 67788
rect 162316 66882 162372 66892
rect 162092 65986 162148 65996
rect 163772 60676 163828 380492
rect 172172 378980 172228 378990
rect 166348 378868 166404 378878
rect 166012 377188 166068 377198
rect 163996 375620 164052 375630
rect 163996 61572 164052 375564
rect 164556 374612 164612 374622
rect 164332 374052 164388 374062
rect 164108 373940 164164 373950
rect 164108 63364 164164 373884
rect 164220 372372 164276 372382
rect 164220 65156 164276 372316
rect 164220 65090 164276 65100
rect 164108 63298 164164 63308
rect 164332 62468 164388 373996
rect 164556 64260 164612 374556
rect 164556 64194 164612 64204
rect 164332 62402 164388 62412
rect 163996 61506 164052 61516
rect 163772 60610 163828 60620
rect 166012 57316 166068 377132
rect 166348 60340 166404 378812
rect 166796 368900 166852 368910
rect 166796 366212 166852 368844
rect 166796 366146 166852 366156
rect 167244 365428 167300 365438
rect 167244 359604 167300 365372
rect 167244 359538 167300 359548
rect 167580 364532 167636 364542
rect 167580 354452 167636 364476
rect 171388 359492 171444 359502
rect 167580 354386 167636 354396
rect 170492 354452 170548 354462
rect 167132 348740 167188 348750
rect 167132 346164 167188 348684
rect 167132 346098 167188 346108
rect 170492 324660 170548 354396
rect 171388 349524 171444 359436
rect 171388 349458 171444 349468
rect 170492 324594 170548 324604
rect 171612 300692 171668 300702
rect 170940 79044 170996 79054
rect 170940 75880 170996 78988
rect 171612 75880 171668 300636
rect 172172 79940 172228 378924
rect 172396 366212 172452 366222
rect 172172 79874 172228 79884
rect 172284 298788 172340 298798
rect 172284 75880 172340 298732
rect 172396 243684 172452 366156
rect 420924 362852 420980 362862
rect 172396 243618 172452 243628
rect 173852 349524 173908 349534
rect 173852 99092 173908 349468
rect 173964 345716 174020 345726
rect 173964 337708 174020 345660
rect 420924 337764 420980 362796
rect 173964 337652 174132 337708
rect 420924 337698 420980 337708
rect 173852 99026 173908 99036
rect 173964 324660 174020 324670
rect 173628 93380 173684 93390
rect 172956 79044 173012 79054
rect 172956 75880 173012 78988
rect 173628 75880 173684 93324
rect 173964 83748 174020 324604
rect 174076 105252 174132 337652
rect 419132 333508 419188 333518
rect 418348 314244 418404 314254
rect 378364 308308 378420 308318
rect 378364 308242 378420 308252
rect 351036 308084 351092 308094
rect 385084 308084 385140 308094
rect 189308 305732 189364 305742
rect 185724 305620 185780 305630
rect 183484 305396 183540 305406
rect 183036 305284 183092 305294
rect 182588 305172 182644 305182
rect 177212 305060 177268 305070
rect 176204 300692 176260 300702
rect 174300 299908 174356 299918
rect 174076 105186 174132 105196
rect 174188 243684 174244 243694
rect 174188 85204 174244 243628
rect 174188 85138 174244 85148
rect 173964 83682 174020 83692
rect 174300 75880 174356 299852
rect 176204 298900 176260 300636
rect 176204 298844 176792 298900
rect 177212 298872 177268 305004
rect 179004 304948 179060 304958
rect 178108 303604 178164 303614
rect 177660 301588 177716 301598
rect 177660 298872 177716 301532
rect 178108 298872 178164 303548
rect 178556 303492 178612 303502
rect 178556 298872 178612 303436
rect 179004 298872 179060 304892
rect 180348 303940 180404 303950
rect 179900 303268 179956 303278
rect 179452 301700 179508 301710
rect 179452 298872 179508 301644
rect 179900 298872 179956 303212
rect 180348 298872 180404 303884
rect 180796 303828 180852 303838
rect 180796 298872 180852 303772
rect 181244 303716 181300 303726
rect 181244 298872 181300 303660
rect 182140 302036 182196 302046
rect 181692 301924 181748 301934
rect 181692 298872 181748 301868
rect 182140 298872 182196 301980
rect 182588 298872 182644 305116
rect 183036 298872 183092 305228
rect 183484 298872 183540 305340
rect 184380 303380 184436 303390
rect 183932 301812 183988 301822
rect 183932 298872 183988 301756
rect 184380 298872 184436 303324
rect 185724 298872 185780 305564
rect 187964 305508 188020 305518
rect 186620 304052 186676 304062
rect 186172 302260 186228 302270
rect 186172 298872 186228 302204
rect 186620 298872 186676 303996
rect 187068 303156 187124 303166
rect 187068 298872 187124 303100
rect 187516 300020 187572 300030
rect 187516 298872 187572 299964
rect 187964 298872 188020 305452
rect 188860 302372 188916 302382
rect 188412 301476 188468 301486
rect 188412 298872 188468 301420
rect 188860 298872 188916 302316
rect 189308 298872 189364 305676
rect 191100 305060 191156 308056
rect 191100 304994 191156 305004
rect 189756 304836 189812 304846
rect 189756 298872 189812 304780
rect 190204 302148 190260 302158
rect 190204 298872 190260 302092
rect 191548 301588 191604 308056
rect 191996 303604 192052 308056
rect 191996 303538 192052 303548
rect 192444 303492 192500 308056
rect 192892 304948 192948 308056
rect 192892 304882 192948 304892
rect 192444 303426 192500 303436
rect 192892 304724 192948 304734
rect 192444 303156 192500 303166
rect 191996 303044 192052 303054
rect 191548 301522 191604 301532
rect 191772 302932 191828 302942
rect 191100 299124 191156 299134
rect 191100 298872 191156 299068
rect 191772 298900 191828 302876
rect 191576 298844 191828 298900
rect 191996 298872 192052 302988
rect 192444 298872 192500 303100
rect 192892 298872 192948 304668
rect 193340 301700 193396 308056
rect 193788 303940 193844 308056
rect 193788 303874 193844 303884
rect 194236 303828 194292 308056
rect 194236 303762 194292 303772
rect 194684 303716 194740 308056
rect 194684 303650 194740 303660
rect 193340 301634 193396 301644
rect 193564 303604 193620 303614
rect 193564 298900 193620 303548
rect 193368 298844 193620 298900
rect 193788 303492 193844 303502
rect 193788 298872 193844 303436
rect 195132 301924 195188 308056
rect 195580 302036 195636 308056
rect 196028 305172 196084 308056
rect 196476 305284 196532 308056
rect 196924 305396 196980 308056
rect 196924 305330 196980 305340
rect 197260 308028 197400 308084
rect 196476 305218 196532 305228
rect 196028 305106 196084 305116
rect 195580 301970 195636 301980
rect 196028 304612 196084 304622
rect 195132 301858 195188 301868
rect 195580 301700 195636 301710
rect 194684 301588 194740 301598
rect 194236 301252 194292 301262
rect 194236 298872 194292 301196
rect 194684 298872 194740 301532
rect 195132 301364 195188 301374
rect 195132 298872 195188 301308
rect 195580 298872 195636 301644
rect 196028 298872 196084 304556
rect 197260 301812 197316 308028
rect 197820 303268 197876 308056
rect 197820 303202 197876 303212
rect 197932 303716 197988 303726
rect 197260 301746 197316 301756
rect 197372 302036 197428 302046
rect 197372 298872 197428 301980
rect 197932 298900 197988 303660
rect 198268 303380 198324 308056
rect 198716 305620 198772 308056
rect 198716 305554 198772 305564
rect 199052 308028 199192 308084
rect 198268 303314 198324 303324
rect 198492 305396 198548 305406
rect 198492 298900 198548 305340
rect 197848 298844 197988 298900
rect 198296 298844 198548 298900
rect 198716 305172 198772 305182
rect 198716 298872 198772 305116
rect 199052 302260 199108 308028
rect 199612 304052 199668 308056
rect 199612 303986 199668 303996
rect 199724 305060 199780 305070
rect 199052 302194 199108 302204
rect 199164 303268 199220 303278
rect 199164 298872 199220 303212
rect 199724 298900 199780 305004
rect 200060 304500 200116 308056
rect 200060 304434 200116 304444
rect 199640 298844 199780 298900
rect 200060 303828 200116 303838
rect 200060 298872 200116 303772
rect 200508 300020 200564 308056
rect 200844 301812 200900 301822
rect 200508 299954 200564 299964
rect 200732 301756 200844 301812
rect 200732 298900 200788 301756
rect 200844 301746 200900 301756
rect 200956 301476 201012 308056
rect 201404 305508 201460 308056
rect 201404 305442 201460 305452
rect 201404 305284 201460 305294
rect 201292 301924 201348 301934
rect 200956 301410 201012 301420
rect 201180 301868 201292 301924
rect 201180 298900 201236 301868
rect 201292 301858 201348 301868
rect 200536 298844 200788 298900
rect 200984 298844 201236 298900
rect 201404 298872 201460 305228
rect 201852 302372 201908 308056
rect 202300 305732 202356 308056
rect 202300 305666 202356 305676
rect 202748 304836 202804 308056
rect 202748 304770 202804 304780
rect 203084 305508 203140 305518
rect 201852 302306 201908 302316
rect 202748 304052 202804 304062
rect 202300 301476 202356 301486
rect 201852 299236 201908 299246
rect 201852 298872 201908 299180
rect 202300 298872 202356 301420
rect 202748 298872 202804 303996
rect 203084 298900 203140 305452
rect 203196 302148 203252 308056
rect 203644 302932 203700 308056
rect 204092 303044 204148 308056
rect 204092 302978 204148 302988
rect 204316 303940 204372 303950
rect 203644 302866 203700 302876
rect 203196 302082 203252 302092
rect 203644 302708 203700 302718
rect 203084 298844 203224 298900
rect 203644 298872 203700 302652
rect 204316 298900 204372 303884
rect 204540 303156 204596 308056
rect 204540 303090 204596 303100
rect 204764 304948 204820 304958
rect 204120 298844 204372 298900
rect 204540 302932 204596 302942
rect 204540 298872 204596 302876
rect 204764 299012 204820 304892
rect 204988 304724 205044 308056
rect 204988 304658 205044 304668
rect 205436 303604 205492 308056
rect 205436 303538 205492 303548
rect 204764 298946 204820 298956
rect 204988 303380 205044 303390
rect 204988 298872 205044 303324
rect 205436 303156 205492 303166
rect 205436 298872 205492 303100
rect 205884 301252 205940 308056
rect 205884 301186 205940 301196
rect 206108 305620 206164 305630
rect 206108 298900 206164 305564
rect 206332 303492 206388 308056
rect 206668 308028 206808 308084
rect 206332 303426 206388 303436
rect 206556 305732 206612 305742
rect 206556 298900 206612 305676
rect 206668 301588 206724 308028
rect 206668 301522 206724 301532
rect 206780 302148 206836 302158
rect 205912 298844 206164 298900
rect 206360 298844 206612 298900
rect 206780 298872 206836 302092
rect 207228 301364 207284 308056
rect 207676 301700 207732 308056
rect 208124 304612 208180 308056
rect 208124 304546 208180 304556
rect 208572 302036 208628 308056
rect 209020 303716 209076 308056
rect 209468 305396 209524 308056
rect 209468 305330 209524 305340
rect 209804 305396 209860 305406
rect 209468 304836 209524 304846
rect 209020 303650 209076 303660
rect 209132 304724 209188 304734
rect 208572 301970 208628 301980
rect 207676 301634 207732 301644
rect 208124 301700 208180 301710
rect 207228 301298 207284 301308
rect 207228 299348 207284 299358
rect 207228 298872 207284 299292
rect 208124 298872 208180 301644
rect 208572 300804 208628 300814
rect 208572 298872 208628 300748
rect 209132 298900 209188 304668
rect 209048 298844 209188 298900
rect 209468 298872 209524 304780
rect 209804 298900 209860 305340
rect 209916 305172 209972 308056
rect 209916 305106 209972 305116
rect 210364 303268 210420 308056
rect 210812 303828 210868 308056
rect 211260 305060 211316 308056
rect 211260 304994 211316 305004
rect 210812 303762 210868 303772
rect 211260 304612 211316 304622
rect 210364 303202 210420 303212
rect 210476 303492 210532 303502
rect 210476 298900 210532 303436
rect 209804 298844 209944 298900
rect 210392 298844 210532 298900
rect 210812 303268 210868 303278
rect 210812 298872 210868 303212
rect 211260 298872 211316 304556
rect 211708 301812 211764 308056
rect 211708 301746 211764 301756
rect 211932 302596 211988 302606
rect 211932 298900 211988 302540
rect 212156 301924 212212 308056
rect 212604 305284 212660 308056
rect 212604 305218 212660 305228
rect 213052 304052 213108 308056
rect 213500 305508 213556 308056
rect 213500 305442 213556 305452
rect 213052 303986 213108 303996
rect 212156 301858 212212 301868
rect 212380 303604 212436 303614
rect 212380 298900 212436 303548
rect 213948 302708 214004 308056
rect 213948 302642 214004 302652
rect 214172 304164 214228 304174
rect 213500 302484 213556 302494
rect 211736 298844 211988 298900
rect 212184 298844 212436 298900
rect 212604 299572 212660 299582
rect 212604 298872 212660 299516
rect 213052 298900 213108 298910
rect 213500 298872 213556 302428
rect 214172 298900 214228 304108
rect 214396 303940 214452 308056
rect 214396 303874 214452 303884
rect 214620 304276 214676 304286
rect 214620 298900 214676 304220
rect 214844 302932 214900 308056
rect 215292 303156 215348 308056
rect 215292 303090 215348 303100
rect 215516 305508 215572 305518
rect 214844 302866 214900 302876
rect 213976 298844 214228 298900
rect 214424 298844 214676 298900
rect 214844 301924 214900 301934
rect 214844 298872 214900 301868
rect 215516 298900 215572 305452
rect 215740 303380 215796 308056
rect 216188 305620 216244 308056
rect 216636 305732 216692 308056
rect 216636 305666 216692 305676
rect 216188 305554 216244 305564
rect 215740 303314 215796 303324
rect 215964 305060 216020 305070
rect 215964 298900 216020 305004
rect 215320 298844 215572 298900
rect 215768 298844 216020 298900
rect 216188 303940 216244 303950
rect 216188 298872 216244 303884
rect 216636 303828 216692 303838
rect 216636 298872 216692 303772
rect 217084 302148 217140 308056
rect 217084 302082 217140 302092
rect 217084 301812 217140 301822
rect 217084 298872 217140 301756
rect 217532 301700 217588 308056
rect 217532 301634 217588 301644
rect 217756 303380 217812 303390
rect 217756 298900 217812 303324
rect 217980 300804 218036 308056
rect 218428 304724 218484 308056
rect 218876 304836 218932 308056
rect 219324 305396 219380 308056
rect 219324 305330 219380 305340
rect 218876 304770 218932 304780
rect 218428 304658 218484 304668
rect 219324 304052 219380 304062
rect 218876 302260 218932 302270
rect 217980 300738 218036 300748
rect 218428 300804 218484 300814
rect 217560 298844 217812 298900
rect 217980 299460 218036 299470
rect 217980 298872 218036 299404
rect 218428 298872 218484 300748
rect 218876 298872 218932 302204
rect 219324 298872 219380 303996
rect 219772 303268 219828 308056
rect 220220 303492 220276 308056
rect 220668 304612 220724 308056
rect 220668 304546 220724 304556
rect 220220 303426 220276 303436
rect 219772 303202 219828 303212
rect 221116 302596 221172 308056
rect 221564 303604 221620 308056
rect 221564 303538 221620 303548
rect 221788 308028 222040 308084
rect 221116 302530 221172 302540
rect 221564 303268 221620 303278
rect 220668 302148 220724 302158
rect 220220 302036 220276 302046
rect 219772 301700 219828 301710
rect 219772 298872 219828 301644
rect 220220 298872 220276 301980
rect 220668 298872 220724 302092
rect 221116 301028 221172 301038
rect 221116 298872 221172 300972
rect 221564 298872 221620 303212
rect 221788 302484 221844 308028
rect 221788 302418 221844 302428
rect 222012 305172 222068 305182
rect 222012 298872 222068 305116
rect 222460 304164 222516 308056
rect 222908 304276 222964 308056
rect 222908 304210 222964 304220
rect 222460 304098 222516 304108
rect 222460 303492 222516 303502
rect 222460 298872 222516 303436
rect 223356 301924 223412 308056
rect 223356 301858 223412 301868
rect 223692 305844 223748 305854
rect 222908 300916 222964 300926
rect 222908 298872 222964 300860
rect 223356 299572 223412 299582
rect 223356 298872 223412 299516
rect 223692 298900 223748 305788
rect 223804 305508 223860 308056
rect 223804 305442 223860 305452
rect 224252 303940 224308 308056
rect 224252 303874 224308 303884
rect 224476 305284 224532 305294
rect 224476 298900 224532 305228
rect 224700 305060 224756 308056
rect 224700 304994 224756 305004
rect 223692 298844 223832 298900
rect 224280 298844 224532 298900
rect 224700 303940 224756 303950
rect 224700 298872 224756 303884
rect 225148 303828 225204 308056
rect 225148 303762 225204 303772
rect 225372 304276 225428 304286
rect 225372 298900 225428 304220
rect 225596 301812 225652 308056
rect 225596 301746 225652 301756
rect 225820 304388 225876 304398
rect 225820 298900 225876 304332
rect 226044 303380 226100 308056
rect 226044 303314 226100 303324
rect 226268 304500 226324 304510
rect 226268 298900 226324 304444
rect 226492 302260 226548 308056
rect 226492 302194 226548 302204
rect 226716 304612 226772 304622
rect 226716 298900 226772 304556
rect 226940 304052 226996 308056
rect 226940 303986 226996 303996
rect 225176 298844 225428 298900
rect 225624 298844 225876 298900
rect 226072 298844 226324 298900
rect 226520 298844 226772 298900
rect 226940 302484 226996 302494
rect 226940 298872 226996 302428
rect 227388 301700 227444 308056
rect 227836 302036 227892 308056
rect 228284 302148 228340 308056
rect 228284 302082 228340 302092
rect 228396 305060 228452 305070
rect 227836 301970 227892 301980
rect 228284 301924 228340 301934
rect 227388 301634 227444 301644
rect 227836 301812 227892 301822
rect 227388 301364 227444 301374
rect 227388 298872 227444 301308
rect 227836 298872 227892 301756
rect 228284 298872 228340 301868
rect 228396 299908 228452 305004
rect 228732 303268 228788 308056
rect 228732 303202 228788 303212
rect 229180 301028 229236 308056
rect 229628 305172 229684 308056
rect 229628 305106 229684 305116
rect 229180 300962 229236 300972
rect 229628 303716 229684 303726
rect 228396 299842 228452 299852
rect 228732 300804 228788 300814
rect 228732 298872 228788 300748
rect 229180 300804 229236 300814
rect 229180 298872 229236 300748
rect 229628 298872 229684 303660
rect 229964 303604 230020 303614
rect 229964 298900 230020 303548
rect 230076 303492 230132 308056
rect 230076 303426 230132 303436
rect 230524 300916 230580 308056
rect 230972 305284 231028 308056
rect 230972 305218 231028 305228
rect 230524 300850 230580 300860
rect 230748 304836 230804 304846
rect 230748 298900 230804 304780
rect 231420 303940 231476 308056
rect 231420 303874 231476 303884
rect 231644 305396 231700 305406
rect 229964 298844 230104 298900
rect 230552 298844 230804 298900
rect 230972 302036 231028 302046
rect 230972 298872 231028 301980
rect 231644 298900 231700 305340
rect 231868 304276 231924 308056
rect 232316 304388 232372 308056
rect 232764 304500 232820 308056
rect 232764 304434 232820 304444
rect 232876 308028 233240 308084
rect 232316 304322 232372 304332
rect 231868 304210 231924 304220
rect 232316 303380 232372 303390
rect 231448 298844 231700 298900
rect 231868 300804 231924 300814
rect 231868 298872 231924 300748
rect 232316 298872 232372 303324
rect 232876 302484 232932 308028
rect 232876 302418 232932 302428
rect 232988 305620 233044 305630
rect 232988 298900 233044 305564
rect 233660 304612 233716 308056
rect 233660 304546 233716 304556
rect 232792 298844 233044 298900
rect 233212 304276 233268 304286
rect 233212 298872 233268 304220
rect 233660 304164 233716 304174
rect 233660 298872 233716 304108
rect 234108 301364 234164 308056
rect 234108 301298 234164 301308
rect 234332 305508 234388 305518
rect 234332 298900 234388 305452
rect 234556 301812 234612 308056
rect 234892 308028 235032 308084
rect 234556 301746 234612 301756
rect 234780 305172 234836 305182
rect 234780 298900 234836 305116
rect 234892 301924 234948 308028
rect 234892 301858 234948 301868
rect 235004 303828 235060 303838
rect 234136 298844 234388 298900
rect 234584 298844 234836 298900
rect 235004 298872 235060 303772
rect 235452 303716 235508 308056
rect 235452 303650 235508 303660
rect 235564 308028 235928 308084
rect 235564 303604 235620 308028
rect 236348 304836 236404 308056
rect 236348 304770 236404 304780
rect 236572 305284 236628 305294
rect 235564 303538 235620 303548
rect 235900 304052 235956 304062
rect 235452 303492 235508 303502
rect 235452 298872 235508 303436
rect 235900 298872 235956 303996
rect 236572 298900 236628 305228
rect 236376 298844 236628 298900
rect 236684 303940 236740 303950
rect 236684 298900 236740 303884
rect 236796 302036 236852 308056
rect 237244 305396 237300 308056
rect 237244 305330 237300 305340
rect 236796 301970 236852 301980
rect 237244 301252 237300 301262
rect 236684 298844 236824 298900
rect 237244 298872 237300 301196
rect 237692 300804 237748 308056
rect 238140 303380 238196 308056
rect 238588 305620 238644 308056
rect 238588 305554 238644 305564
rect 239036 305508 239092 308056
rect 239036 305442 239092 305452
rect 239484 305172 239540 308056
rect 239484 305106 239540 305116
rect 239932 303828 239988 308056
rect 239932 303762 239988 303772
rect 240156 304612 240212 304622
rect 238140 303314 238196 303324
rect 237692 300738 237748 300748
rect 238140 302820 238196 302830
rect 237692 299572 237748 299582
rect 237692 298872 237748 299516
rect 238140 298872 238196 302764
rect 238588 302372 238644 302382
rect 238588 298872 238644 302316
rect 239036 302260 239092 302270
rect 239036 298872 239092 302204
rect 239484 302148 239540 302158
rect 239484 298872 239540 302092
rect 240156 298900 240212 304556
rect 240380 303492 240436 308056
rect 240828 304052 240884 308056
rect 241276 305284 241332 308056
rect 241276 305218 241332 305228
rect 240828 303986 240884 303996
rect 241276 304724 241332 304734
rect 240380 303426 240436 303436
rect 239960 298844 240212 298900
rect 240380 302036 240436 302046
rect 240380 298872 240436 301980
rect 240828 301924 240884 301934
rect 240828 298872 240884 301868
rect 241276 298872 241332 304668
rect 241724 303940 241780 308056
rect 241724 303874 241780 303884
rect 241836 304836 241892 304846
rect 241836 298900 241892 304780
rect 242172 301252 242228 308056
rect 242620 302372 242676 308056
rect 242620 302306 242676 302316
rect 242732 308028 243096 308084
rect 243180 308028 243544 308084
rect 242732 302260 242788 308028
rect 243068 303156 243124 303166
rect 242956 302596 243012 302606
rect 242732 302194 242788 302204
rect 242844 302540 242956 302596
rect 242172 301186 242228 301196
rect 241752 298844 241892 298900
rect 242172 300804 242228 300814
rect 242172 298872 242228 300748
rect 242844 298900 242900 302540
rect 242956 302530 243012 302540
rect 242648 298844 242900 298900
rect 243068 298872 243124 303100
rect 243180 302148 243236 308028
rect 243964 304612 244020 308056
rect 243964 304546 244020 304556
rect 244076 308028 244440 308084
rect 244524 308028 244888 308084
rect 243964 304388 244020 304398
rect 243180 302082 243236 302092
rect 243516 303268 243572 303278
rect 243516 298872 243572 303212
rect 243964 298872 244020 304332
rect 244076 302036 244132 308028
rect 244076 301970 244132 301980
rect 244412 304500 244468 304510
rect 244412 298872 244468 304444
rect 244524 301924 244580 308028
rect 245308 304724 245364 308056
rect 245756 304836 245812 308056
rect 245756 304770 245812 304780
rect 245308 304658 245364 304668
rect 246204 303156 246260 308056
rect 246652 303268 246708 308056
rect 247100 304388 247156 308056
rect 247548 304500 247604 308056
rect 247548 304434 247604 304444
rect 247660 308028 248024 308084
rect 247100 304322 247156 304332
rect 246652 303202 246708 303212
rect 246204 303090 246260 303100
rect 247548 303156 247604 303166
rect 245308 303044 245364 303054
rect 244524 301858 244580 301868
rect 244860 302372 244916 302382
rect 244860 298872 244916 302316
rect 245308 298872 245364 302988
rect 245756 302260 245812 302270
rect 245756 298872 245812 302204
rect 246204 302148 246260 302158
rect 246204 298872 246260 302092
rect 247100 301252 247156 301262
rect 246876 299012 246932 299022
rect 246876 298900 246932 298956
rect 246680 298844 246932 298900
rect 247100 298872 247156 301196
rect 247548 298872 247604 303100
rect 247660 302372 247716 308028
rect 247660 302306 247716 302316
rect 247996 303268 248052 303278
rect 247996 298872 248052 303212
rect 248444 303044 248500 308056
rect 248444 302978 248500 302988
rect 248892 302260 248948 308056
rect 249228 303828 249284 303838
rect 248892 302194 248948 302204
rect 249116 303772 249228 303828
rect 248444 301028 248500 301038
rect 248444 298872 248500 300972
rect 249116 298900 249172 303772
rect 249228 303762 249284 303772
rect 249340 302148 249396 308056
rect 249676 304052 249732 304062
rect 249340 302082 249396 302092
rect 249564 303996 249676 304052
rect 249564 298900 249620 303996
rect 249676 303986 249732 303996
rect 249788 303156 249844 308056
rect 250236 303268 250292 308056
rect 250236 303202 250292 303212
rect 249788 303090 249844 303100
rect 250684 301028 250740 308056
rect 250684 300962 250740 300972
rect 250908 303940 250964 303950
rect 250236 300916 250292 300926
rect 248920 298844 249172 298900
rect 249368 298844 249620 298900
rect 249788 300804 249844 300814
rect 249788 298872 249844 300748
rect 250236 298872 250292 300860
rect 250908 298900 250964 303884
rect 251132 303828 251188 308056
rect 251580 304052 251636 308056
rect 251580 303986 251636 303996
rect 251132 303762 251188 303772
rect 250712 298844 250964 298900
rect 251132 301140 251188 301150
rect 251132 298872 251188 301084
rect 251580 301028 251636 301038
rect 251580 298872 251636 300972
rect 252028 300804 252084 308056
rect 252364 308028 252504 308084
rect 252588 308028 252952 308084
rect 253036 308028 253400 308084
rect 252252 305508 252308 305518
rect 252028 300738 252084 300748
rect 252140 305506 252308 305508
rect 252140 305454 252254 305506
rect 252306 305454 252308 305506
rect 252140 305452 252308 305454
rect 252140 298900 252196 305452
rect 252252 305442 252308 305452
rect 252364 300916 252420 308028
rect 252364 300850 252420 300860
rect 252476 304052 252532 304062
rect 252056 298844 252196 298900
rect 252476 298872 252532 303996
rect 252588 303940 252644 308028
rect 253036 305506 253092 308028
rect 253036 305454 253038 305506
rect 253090 305454 253092 305506
rect 253036 305442 253092 305454
rect 253820 304052 253876 308056
rect 253820 303986 253876 303996
rect 252588 303874 252644 303884
rect 252924 303940 252980 303950
rect 252588 301252 252644 301262
rect 252588 300916 252644 301196
rect 252588 300850 252644 300860
rect 252924 298872 252980 303884
rect 254268 303940 254324 308056
rect 254268 303874 254324 303884
rect 253372 303828 253428 303838
rect 253372 298872 253428 303772
rect 254716 303828 254772 308056
rect 254716 303762 254772 303772
rect 254828 308028 255192 308084
rect 254828 303604 254884 308028
rect 253932 303548 254884 303604
rect 253932 298900 253988 303548
rect 255164 302932 255220 302942
rect 254716 302820 254772 302830
rect 253848 298844 253988 298900
rect 254268 302708 254324 302718
rect 254268 298872 254324 302652
rect 254716 298872 254772 302764
rect 255164 298872 255220 302876
rect 255612 302708 255668 308056
rect 256060 302820 256116 308056
rect 256508 302932 256564 308056
rect 256508 302866 256564 302876
rect 256620 308028 256984 308084
rect 257068 308028 257432 308084
rect 257516 308028 257880 308084
rect 257964 308028 258328 308084
rect 256060 302754 256116 302764
rect 255612 302642 255668 302652
rect 256284 302708 256340 302718
rect 256284 298900 256340 302652
rect 256620 298900 256676 308028
rect 257068 302428 257124 308028
rect 256088 298844 256340 298900
rect 256536 298844 256676 298900
rect 256956 302372 257124 302428
rect 256956 298872 257012 302372
rect 257516 298900 257572 308028
rect 257964 298900 258020 308028
rect 258748 302428 258804 308056
rect 258524 302372 258804 302428
rect 258860 308028 259224 308084
rect 259308 308028 259672 308084
rect 259756 308028 260120 308084
rect 260568 308028 260820 308084
rect 261016 308028 261268 308084
rect 261464 308028 261716 308084
rect 261912 308028 262052 308084
rect 262360 308028 262612 308084
rect 262808 308028 263060 308084
rect 263256 308028 263508 308084
rect 258524 298900 258580 302372
rect 258860 298900 258916 308028
rect 259308 298900 259364 308028
rect 259756 298900 259812 308028
rect 257432 298844 257572 298900
rect 257880 298844 258020 298900
rect 258328 298844 258580 298900
rect 258776 298844 258916 298900
rect 259224 298844 259364 298900
rect 259672 298844 259812 298900
rect 260540 300804 260596 300814
rect 260540 298872 260596 300748
rect 260764 298900 260820 308028
rect 261212 298900 261268 308028
rect 261660 298900 261716 308028
rect 261996 305172 262052 308028
rect 261996 305116 262164 305172
rect 262108 298900 262164 305116
rect 262556 298900 262612 308028
rect 263004 298900 263060 308028
rect 263452 298900 263508 308028
rect 263676 305284 263732 308056
rect 264152 308028 264404 308084
rect 264600 308028 264852 308084
rect 265048 308028 265300 308084
rect 265496 308028 265748 308084
rect 265944 308028 266196 308084
rect 266392 308028 266644 308084
rect 266840 308028 267092 308084
rect 267288 308028 267540 308084
rect 267736 308028 267988 308084
rect 268184 308028 268436 308084
rect 268632 308028 268772 308084
rect 269080 308028 269332 308084
rect 269528 308028 269780 308084
rect 269976 308028 270228 308084
rect 263676 305228 263844 305284
rect 263788 298900 263844 305228
rect 264348 298900 264404 308028
rect 264796 298900 264852 308028
rect 265244 305284 265300 308028
rect 265244 305228 265524 305284
rect 260764 298844 261016 298900
rect 261212 298844 261464 298900
rect 261660 298844 261912 298900
rect 262108 298844 262360 298900
rect 262556 298844 262808 298900
rect 263004 298844 263256 298900
rect 263452 298844 263704 298900
rect 263788 298844 264152 298900
rect 264348 298844 264600 298900
rect 264796 298844 265048 298900
rect 265468 298872 265524 305228
rect 265692 298900 265748 308028
rect 266140 298900 266196 308028
rect 266588 298900 266644 308028
rect 267036 305788 267092 308028
rect 267036 305732 267204 305788
rect 267148 298900 267204 305732
rect 267484 298900 267540 308028
rect 267932 298900 267988 308028
rect 268380 298900 268436 308028
rect 268716 305172 268772 308028
rect 268716 305116 268884 305172
rect 268828 298900 268884 305116
rect 269276 298900 269332 308028
rect 269724 298900 269780 308028
rect 270172 298900 270228 308028
rect 270396 305396 270452 308056
rect 270872 308028 271124 308084
rect 270396 305340 270900 305396
rect 265692 298844 265944 298900
rect 266140 298844 266392 298900
rect 266588 298844 266840 298900
rect 267148 298844 267288 298900
rect 267484 298844 267736 298900
rect 267932 298844 268184 298900
rect 268380 298844 268632 298900
rect 268828 298844 269080 298900
rect 269276 298844 269528 298900
rect 269724 298844 269976 298900
rect 270172 298844 270424 298900
rect 270844 298872 270900 305340
rect 271068 298900 271124 308028
rect 271292 304948 271348 308056
rect 271740 305508 271796 308056
rect 272188 305732 272244 308056
rect 272188 305666 272244 305676
rect 271740 305442 271796 305452
rect 272636 305172 272692 308056
rect 272636 305106 272692 305116
rect 272972 305396 273028 305406
rect 271292 304882 271348 304892
rect 271068 298844 271320 298900
rect 213052 298834 213108 298844
rect 207676 298788 207732 298798
rect 207676 298722 207732 298732
rect 196924 298676 196980 298686
rect 196924 298610 196980 298620
rect 190652 298564 190708 298574
rect 190652 298498 190708 298508
rect 196476 298452 196532 298462
rect 196476 298386 196532 298396
rect 184828 298340 184884 298350
rect 184828 298274 184884 298284
rect 185276 298340 185332 298350
rect 185276 298274 185332 298284
rect 255612 298340 255668 298350
rect 255612 298274 255668 298284
rect 260092 298340 260148 298350
rect 260092 298274 260148 298284
rect 191100 102004 191156 102014
rect 183036 101892 183092 101902
rect 181020 101780 181076 101790
rect 178332 101668 178388 101678
rect 174972 100212 175028 100222
rect 174972 75880 175028 100156
rect 177772 99092 177828 99102
rect 177772 96740 177828 99036
rect 177772 96674 177828 96684
rect 177212 94948 177268 94958
rect 176988 83188 177044 83198
rect 175644 80612 175700 80622
rect 175644 75880 175700 80556
rect 176316 80276 176372 80286
rect 176316 75880 176372 80220
rect 176988 75880 177044 83132
rect 177212 80612 177268 94892
rect 177212 80546 177268 80556
rect 177660 80612 177716 80622
rect 177660 75880 177716 80556
rect 178332 75880 178388 101612
rect 179676 99540 179732 99550
rect 179676 96628 179732 99484
rect 179676 96562 179732 96572
rect 180572 98532 180628 98542
rect 179676 91588 179732 91598
rect 179004 79828 179060 79838
rect 179004 75880 179060 79772
rect 179676 75880 179732 91532
rect 180348 83300 180404 83310
rect 180348 75880 180404 83244
rect 180572 80612 180628 98476
rect 180572 80546 180628 80556
rect 181020 75880 181076 101724
rect 181692 93492 181748 93502
rect 181692 75880 181748 93436
rect 182364 91700 182420 91710
rect 182364 75880 182420 91644
rect 183036 75880 183092 101836
rect 188412 98644 188468 98654
rect 185724 98420 185780 98430
rect 183708 95172 183764 95182
rect 183708 75880 183764 95116
rect 184380 91812 184436 91822
rect 184380 75880 184436 91756
rect 185052 80612 185108 80622
rect 185052 75880 185108 80556
rect 185724 75880 185780 98364
rect 187292 91924 187348 91934
rect 186396 89908 186452 89918
rect 186396 75880 186452 89852
rect 187068 81508 187124 81518
rect 187068 75880 187124 81452
rect 187292 80612 187348 91868
rect 187292 80546 187348 80556
rect 187740 86548 187796 86558
rect 187740 75880 187796 86492
rect 188412 75880 188468 98588
rect 189084 96852 189140 96862
rect 189084 75880 189140 96796
rect 189532 80612 189588 80622
rect 189532 75908 189588 80556
rect 190428 80612 190484 80622
rect 189532 75852 189784 75908
rect 190428 75880 190484 80556
rect 191100 75880 191156 101948
rect 199836 101556 199892 101566
rect 192444 100324 192500 100334
rect 191772 86660 191828 86670
rect 191772 75880 191828 86604
rect 192444 75880 192500 100268
rect 195804 96964 195860 96974
rect 195692 92036 195748 92046
rect 192668 90020 192724 90030
rect 192668 80612 192724 89964
rect 195132 88228 195188 88238
rect 193788 86772 193844 86782
rect 192668 80546 192724 80556
rect 193116 80612 193172 80622
rect 193116 75880 193172 80556
rect 193788 75880 193844 86716
rect 194460 78260 194516 78270
rect 194460 75880 194516 78204
rect 195132 75880 195188 88172
rect 195692 80612 195748 91980
rect 195692 80546 195748 80556
rect 195804 75880 195860 96908
rect 198156 90244 198212 90254
rect 197820 81620 197876 81630
rect 197148 80052 197204 80062
rect 196476 79044 196532 79054
rect 196476 75880 196532 78988
rect 197148 75880 197204 79996
rect 197820 75880 197876 81564
rect 198156 79044 198212 90188
rect 198156 78978 198212 78988
rect 198492 90132 198548 90142
rect 198492 75880 198548 90076
rect 199164 80388 199220 80398
rect 199164 75880 199220 80332
rect 199836 75880 199892 101500
rect 218652 101444 218708 101454
rect 203868 100436 203924 100446
rect 200508 98756 200564 98766
rect 200508 75880 200564 98700
rect 201180 92148 201236 92158
rect 201180 75880 201236 92092
rect 203196 90356 203252 90366
rect 201852 83412 201908 83422
rect 201852 75880 201908 83356
rect 202524 80612 202580 80622
rect 202524 75880 202580 80556
rect 203196 75880 203252 90300
rect 203868 75880 203924 100380
rect 205884 98868 205940 98878
rect 205212 90468 205268 90478
rect 204876 80612 204932 80622
rect 204876 75908 204932 80556
rect 204568 75852 204932 75908
rect 205212 75880 205268 90412
rect 205884 75880 205940 98812
rect 209916 97076 209972 97086
rect 209244 93716 209300 93726
rect 207900 93604 207956 93614
rect 207228 90580 207284 90590
rect 206556 80612 206612 80622
rect 206556 75880 206612 80556
rect 207228 75880 207284 90524
rect 207900 75880 207956 93548
rect 208572 80500 208628 80510
rect 208572 75880 208628 80444
rect 209244 75880 209300 93660
rect 209916 75880 209972 97020
rect 211260 95284 211316 95294
rect 210588 88340 210644 88350
rect 210588 75880 210644 88284
rect 211260 75880 211316 95228
rect 216748 88452 216804 88462
rect 212604 86884 212660 86894
rect 211932 84868 211988 84878
rect 211932 75880 211988 84812
rect 212604 75880 212660 86828
rect 215964 85092 216020 85102
rect 215292 84980 215348 84990
rect 213276 81732 213332 81742
rect 213276 75880 213332 81676
rect 213948 80612 214004 80622
rect 213948 75880 214004 80556
rect 214844 80612 214900 80622
rect 214844 75908 214900 80556
rect 214648 75852 214900 75908
rect 215292 75880 215348 84924
rect 215964 75880 216020 85036
rect 216636 83636 216692 83646
rect 216636 75880 216692 83580
rect 216748 80500 216804 88396
rect 218428 83748 218484 83758
rect 216748 80434 216804 80444
rect 217980 83524 218036 83534
rect 217308 80164 217364 80174
rect 217308 75880 217364 80108
rect 217980 75880 218036 83468
rect 218428 79044 218484 83692
rect 218428 78978 218484 78988
rect 218652 75880 218708 101388
rect 266252 100884 266308 100894
rect 246204 100660 246260 100670
rect 234332 100548 234388 100558
rect 221340 96740 221396 96750
rect 219996 95060 220052 95070
rect 219324 79940 219380 79950
rect 219324 75880 219380 79884
rect 219996 75880 220052 95004
rect 220668 80724 220724 80734
rect 220668 75880 220724 80668
rect 221340 75880 221396 96684
rect 223356 96628 223412 96638
rect 222684 85204 222740 85214
rect 222012 79044 222068 79054
rect 222012 75880 222068 78988
rect 222684 75880 222740 85148
rect 223356 75880 223412 96572
rect 224700 87108 224756 87118
rect 224028 80164 224084 80174
rect 224028 75880 224084 80108
rect 224700 75880 224756 87052
rect 225148 85204 225204 85214
rect 225148 80276 225204 85148
rect 230188 83860 230244 83870
rect 228620 83748 228676 83758
rect 226604 80612 226660 80622
rect 226044 80500 226100 80510
rect 225148 80210 225204 80220
rect 225372 80276 225428 80286
rect 225372 75880 225428 80220
rect 226044 75880 226100 80444
rect 226604 78988 226660 80556
rect 228396 80612 228452 80622
rect 226492 78932 226660 78988
rect 227388 79044 227444 79054
rect 226492 75796 226548 78932
rect 227388 75880 227444 78988
rect 228396 75908 228452 80556
rect 228620 80276 228676 83692
rect 229964 80612 230020 80622
rect 228620 80210 228676 80220
rect 228732 80500 228788 80510
rect 228088 75852 228452 75908
rect 228732 75880 228788 80444
rect 229964 78988 230020 80556
rect 230188 80164 230244 83804
rect 230188 80098 230244 80108
rect 232092 80612 232148 80622
rect 229852 78932 230020 78988
rect 230076 79716 230132 79726
rect 229852 75908 229908 78932
rect 229432 75852 229908 75908
rect 230076 75880 230132 79660
rect 231420 79604 231476 79614
rect 230748 79380 230804 79390
rect 230748 75880 230804 79324
rect 231420 75880 231476 79548
rect 232092 75880 232148 80556
rect 233436 80612 233492 80622
rect 232764 79492 232820 79502
rect 232764 75880 232820 79436
rect 233436 75880 233492 80556
rect 234108 80612 234164 80622
rect 234108 75880 234164 80556
rect 234332 79828 234388 100492
rect 244860 99988 244916 99998
rect 235452 98308 235508 98318
rect 234332 79762 234388 79772
rect 234780 79828 234836 79838
rect 234780 75880 234836 79772
rect 235452 75880 235508 98252
rect 242844 96628 242900 96638
rect 238588 90692 238644 90702
rect 237692 86996 237748 87006
rect 236124 80612 236180 80622
rect 236124 75880 236180 80556
rect 237468 80276 237524 80286
rect 236796 80164 236852 80174
rect 236796 75880 236852 80108
rect 237468 75880 237524 80220
rect 237692 80052 237748 86940
rect 237692 79986 237748 79996
rect 238476 80612 238532 80622
rect 238476 75908 238532 80556
rect 238588 80388 238644 90636
rect 241836 80612 241892 80622
rect 238588 80322 238644 80332
rect 240828 80388 240884 80398
rect 239484 80052 239540 80062
rect 238168 75852 238532 75908
rect 238812 79828 238868 79838
rect 238812 75880 238868 79772
rect 239484 75880 239540 79996
rect 240156 79940 240212 79950
rect 240156 75880 240212 79884
rect 240828 75880 240884 80332
rect 241836 75908 241892 80556
rect 241528 75852 241892 75908
rect 242172 80612 242228 80622
rect 242172 75880 242228 80556
rect 242844 75880 242900 96572
rect 243516 93268 243572 93278
rect 243516 75880 243572 93212
rect 244188 80612 244244 80622
rect 244188 75880 244244 80556
rect 244860 75880 244916 99932
rect 245532 96740 245588 96750
rect 245532 75880 245588 96684
rect 246204 75880 246260 100604
rect 248892 97524 248948 97534
rect 248220 95844 248276 95854
rect 247548 94164 247604 94174
rect 246876 80612 246932 80622
rect 246876 75880 246932 80556
rect 247548 75880 247604 94108
rect 248220 75880 248276 95788
rect 248892 75880 248948 97468
rect 258300 95956 258356 95966
rect 256284 94612 256340 94622
rect 250236 92596 250292 92606
rect 249564 80612 249620 80622
rect 249564 75880 249620 80556
rect 250236 75880 250292 92540
rect 252252 92484 252308 92494
rect 251916 80612 251972 80622
rect 250908 77364 250964 77374
rect 250908 75880 250964 77308
rect 251916 75908 251972 80556
rect 251608 75852 251972 75908
rect 252252 75880 252308 92428
rect 255612 90804 255668 90814
rect 253484 80612 253540 80622
rect 252924 79716 252980 79726
rect 252924 75880 252980 79660
rect 253484 78988 253540 80556
rect 253372 78932 253540 78988
rect 254268 80612 254324 80622
rect 253372 75796 253428 78932
rect 254268 75880 254324 80556
rect 254492 80500 254548 80510
rect 254492 75908 254548 80444
rect 254492 75852 254968 75908
rect 255612 75880 255668 90748
rect 256284 75880 256340 94556
rect 257628 94276 257684 94286
rect 256956 79716 257012 79726
rect 256956 75880 257012 79660
rect 257628 75880 257684 94220
rect 258300 75880 258356 95900
rect 260988 94388 261044 94398
rect 260316 92708 260372 92718
rect 259644 80612 259700 80622
rect 258972 79156 259028 79166
rect 258972 75880 259028 79100
rect 259644 75880 259700 80556
rect 260316 75880 260372 92652
rect 260988 75880 261044 94332
rect 226492 75740 226744 75796
rect 253372 75740 253624 75796
rect 166348 60274 166404 60284
rect 166012 57250 166068 57260
rect 153692 31938 153748 31948
rect 163772 42756 163828 42766
rect 163772 20020 163828 42700
rect 163772 19954 163828 19964
rect 163996 40964 164052 40974
rect 163996 19684 164052 40908
rect 164556 39172 164612 39182
rect 164444 37380 164500 37390
rect 164220 35588 164276 35598
rect 164220 20132 164276 35532
rect 164220 20066 164276 20076
rect 163996 19618 164052 19628
rect 164444 18340 164500 37324
rect 164556 18564 164612 39116
rect 164556 18498 164612 18508
rect 265244 18564 265300 18574
rect 164444 18274 164500 18284
rect 150332 17602 150388 17612
rect 4172 16706 4228 16716
rect 216860 16772 216916 16782
rect 216860 16706 216916 16716
rect 217532 16772 217588 16782
rect 217532 16706 217588 16716
rect 219100 16772 219156 16782
rect 219100 16706 219156 16716
rect 221116 16772 221172 16782
rect 221116 16706 221172 16716
rect 222460 16772 222516 16782
rect 222460 16706 222516 16716
rect 222908 16772 222964 16782
rect 222908 16706 222964 16716
rect 225820 16772 225876 16782
rect 225820 16706 225876 16716
rect 226268 16772 226324 16782
rect 226268 16706 226324 16716
rect 230748 16772 230804 16782
rect 230748 16706 230804 16716
rect 231196 16772 231252 16782
rect 231196 16706 231252 16716
rect 236572 16772 236628 16782
rect 236572 16706 236628 16716
rect 239260 16772 239316 16782
rect 239260 16706 239316 16716
rect 239932 16772 239988 16782
rect 239932 16706 239988 16716
rect 240380 16772 240436 16782
rect 240380 16706 240436 16716
rect 240604 16772 240660 16782
rect 240604 16706 240660 16716
rect 243740 16772 243796 16782
rect 243740 16706 243796 16716
rect 245084 16772 245140 16782
rect 245084 16706 245140 16716
rect 223132 16660 223188 16670
rect 223132 16594 223188 16604
rect 238588 16660 238644 16670
rect 238588 16594 238644 16604
rect 245308 16324 245364 16334
rect 245308 16258 245364 16268
rect 249564 16324 249620 16334
rect 216636 16212 216692 16222
rect 216636 16146 216692 16156
rect 248556 16212 248612 16222
rect 114268 16100 114324 16110
rect 197820 16100 197876 16110
rect 106540 14644 106596 14654
rect 69692 14532 69748 14542
rect 42812 14308 42868 14318
rect 37772 12628 37828 12638
rect 32508 10948 32564 10958
rect 24892 9268 24948 9278
rect 21084 7588 21140 7598
rect 17276 4228 17332 4238
rect 11564 3444 11620 3454
rect 11564 480 11620 3388
rect 13356 3444 13412 3454
rect 13356 480 13412 3388
rect 15372 2548 15428 2558
rect 15372 480 15428 2492
rect 17276 480 17332 4172
rect 19180 4228 19236 4238
rect 19180 480 19236 4172
rect 21084 480 21140 7532
rect 22988 4340 23044 4350
rect 22988 480 23044 4284
rect 24892 480 24948 9212
rect 30604 5908 30660 5918
rect 28700 4340 28756 4350
rect 26796 3444 26852 3454
rect 26796 480 26852 3388
rect 28700 480 28756 4284
rect 30604 480 30660 5852
rect 32508 480 32564 10892
rect 34412 6244 34468 6254
rect 34412 480 34468 6188
rect 36316 4116 36372 4126
rect 36316 480 36372 4060
rect 37772 4116 37828 12572
rect 42028 4116 42084 4126
rect 37772 4050 37828 4060
rect 41916 4060 42028 4116
rect 40124 3780 40180 3790
rect 38220 480 38388 532
rect 40124 480 40180 3724
rect 41916 480 41972 4060
rect 42028 4050 42084 4060
rect 42812 4116 42868 14252
rect 53228 13524 53284 13534
rect 49644 11284 49700 11294
rect 47740 11060 47796 11070
rect 42812 4050 42868 4060
rect 43932 4452 43988 4462
rect 43932 480 43988 4396
rect 45836 480 46004 532
rect 47740 480 47796 11004
rect 49644 480 49700 11228
rect 51548 6804 51604 6814
rect 51548 480 51604 6748
rect 11368 392 11620 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18984 392 19236 480
rect 20888 392 21140 480
rect 22792 392 23044 480
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30408 392 30660 480
rect 32312 392 32564 480
rect 34216 392 34468 480
rect 36120 392 36372 480
rect 38024 476 38388 480
rect 38024 392 38276 476
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 392
rect 38024 -960 38248 392
rect 38332 84 38388 476
rect 38332 18 38388 28
rect 39928 392 40180 480
rect 39928 -960 40152 392
rect 41832 -960 42056 480
rect 43736 392 43988 480
rect 45640 476 46004 480
rect 45640 392 45892 476
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 45948 196 46004 476
rect 45948 130 46004 140
rect 47544 392 47796 480
rect 49448 392 49700 480
rect 51352 392 51604 480
rect 53228 480 53284 13468
rect 54572 12740 54628 12750
rect 54572 6804 54628 12684
rect 54572 6738 54628 6748
rect 61068 9380 61124 9390
rect 55356 3892 55412 3902
rect 55356 480 55412 3836
rect 57260 2660 57316 2670
rect 57260 480 57316 2604
rect 59164 480 59332 532
rect 61068 480 61124 9324
rect 62972 7700 63028 7710
rect 62972 480 63028 7644
rect 66780 6020 66836 6030
rect 64876 480 65044 532
rect 66780 480 66836 5964
rect 68684 4116 68740 4126
rect 68684 480 68740 4060
rect 69692 4116 69748 14476
rect 104636 13748 104692 13758
rect 87500 13636 87556 13646
rect 81452 12964 81508 12974
rect 74172 12852 74228 12862
rect 72492 7588 72548 7598
rect 69692 4050 69748 4060
rect 70476 6132 70532 6142
rect 70476 480 70532 6076
rect 72492 480 72548 7532
rect 53228 392 53480 480
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 392
rect 53256 -960 53480 392
rect 55160 392 55412 480
rect 57064 392 57316 480
rect 58968 476 59332 480
rect 58968 392 59220 476
rect 55160 -960 55384 392
rect 57064 -960 57288 392
rect 58968 -960 59192 392
rect 59276 308 59332 476
rect 59276 242 59332 252
rect 60872 392 61124 480
rect 62776 392 63028 480
rect 64680 476 65044 480
rect 64680 392 64932 476
rect 64988 420 65044 476
rect 65436 420 65492 430
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 64988 364 65436 420
rect 65436 354 65492 364
rect 66584 392 66836 480
rect 68488 392 68740 480
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 480
rect 72296 392 72548 480
rect 74172 480 74228 12796
rect 78204 11172 78260 11182
rect 76412 532 76468 542
rect 76300 480 76412 532
rect 74172 392 74424 480
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 476 76412 480
rect 78204 480 78260 11116
rect 81452 7700 81508 12908
rect 85820 8484 85876 8494
rect 83916 7812 83972 7822
rect 81452 7634 81508 7644
rect 82012 7700 82068 7710
rect 80108 4564 80164 4574
rect 80108 480 80164 4508
rect 82012 480 82068 7644
rect 83916 480 83972 7756
rect 85820 480 85876 8428
rect 76104 392 76356 476
rect 76412 466 76468 476
rect 78008 392 78260 480
rect 79912 392 80164 480
rect 81816 392 82068 480
rect 83720 392 83972 480
rect 85624 392 85876 480
rect 87500 480 87556 13580
rect 92316 13076 92372 13086
rect 89628 9492 89684 9502
rect 89628 480 89684 9436
rect 92316 8484 92372 13020
rect 92316 8418 92372 8428
rect 97244 9604 97300 9614
rect 91532 7924 91588 7934
rect 91532 480 91588 7868
rect 93436 4676 93492 4686
rect 93436 480 93492 4620
rect 95340 2772 95396 2782
rect 95340 480 95396 2716
rect 97244 480 97300 9548
rect 99036 2884 99092 2894
rect 99036 480 99092 2828
rect 102956 756 103012 766
rect 101052 644 101108 654
rect 101052 480 101108 588
rect 102956 480 103012 700
rect 87500 392 87752 480
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89432 392 89684 480
rect 91336 392 91588 480
rect 93240 392 93492 480
rect 95144 392 95396 480
rect 97048 392 97300 480
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100856 392 101108 480
rect 102760 392 103012 480
rect 104636 480 104692 13692
rect 106540 480 106596 14588
rect 112476 9716 112532 9726
rect 108668 8036 108724 8046
rect 108668 480 108724 7980
rect 110572 2996 110628 3006
rect 110572 480 110628 2940
rect 112476 480 112532 9660
rect 114268 480 114324 16044
rect 137004 15988 137060 15998
rect 117964 15204 118020 15214
rect 116732 13188 116788 13198
rect 116284 6356 116340 6366
rect 116284 480 116340 6300
rect 116732 6244 116788 13132
rect 116732 6178 116788 6188
rect 104636 392 104888 480
rect 106540 392 106792 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 392 108724 480
rect 110376 392 110628 480
rect 112280 392 112532 480
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 480
rect 116088 392 116340 480
rect 117964 480 118020 15148
rect 133196 14756 133252 14766
rect 129612 11396 129668 11406
rect 127596 6580 127652 6590
rect 121996 6468 122052 6478
rect 120092 6244 120148 6254
rect 120092 480 120148 6188
rect 121996 480 122052 6412
rect 123900 3108 123956 3118
rect 123900 480 123956 3052
rect 125804 868 125860 878
rect 125804 480 125860 812
rect 127596 480 127652 6524
rect 129612 480 129668 11340
rect 131516 8260 131572 8270
rect 131516 480 131572 8204
rect 117964 392 118216 480
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 392 120148 480
rect 121800 392 122052 480
rect 123704 392 123956 480
rect 125608 392 125860 480
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129416 392 129668 480
rect 131320 392 131572 480
rect 133196 480 133252 14700
rect 135324 11508 135380 11518
rect 135324 480 135380 11452
rect 133196 392 133448 480
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 392 135380 480
rect 137004 480 137060 15932
rect 148428 15876 148484 15886
rect 142828 15316 142884 15326
rect 141036 11284 141092 11294
rect 139132 3220 139188 3230
rect 139132 480 139188 3164
rect 141036 480 141092 11228
rect 142828 480 142884 15260
rect 144620 14868 144676 14878
rect 144620 480 144676 14812
rect 146748 8148 146804 8158
rect 146748 480 146804 8092
rect 137004 392 137256 480
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 392 139188 480
rect 140840 392 141092 480
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 144648 -960 144872 392
rect 146552 392 146804 480
rect 148428 480 148484 15820
rect 167468 14420 167524 14430
rect 154140 13300 154196 13310
rect 152460 9828 152516 9838
rect 150556 3332 150612 3342
rect 150556 480 150612 3276
rect 152460 480 152516 9772
rect 148428 392 148680 480
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 392 150612 480
rect 152264 392 152516 480
rect 154140 480 154196 13244
rect 165564 12068 165620 12078
rect 158172 11620 158228 11630
rect 156156 4788 156212 4798
rect 156156 480 156212 4732
rect 158172 480 158228 11564
rect 160076 9940 160132 9950
rect 160076 480 160132 9884
rect 163884 6692 163940 6702
rect 161980 2436 162036 2446
rect 161980 480 162036 2380
rect 163884 480 163940 6636
rect 154140 392 154392 480
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 480
rect 157976 392 158228 480
rect 159880 392 160132 480
rect 161784 392 162036 480
rect 163688 392 163940 480
rect 165564 480 165620 12012
rect 167468 480 167524 14364
rect 179116 12404 179172 12414
rect 175308 11732 175364 11742
rect 171500 10836 171556 10846
rect 169596 10052 169652 10062
rect 169596 480 169652 9996
rect 171500 480 171556 10780
rect 173404 8372 173460 8382
rect 173404 480 173460 8316
rect 175308 480 175364 11676
rect 177212 9156 177268 9166
rect 177212 480 177268 9100
rect 179116 8260 179172 12348
rect 179116 8194 179172 8204
rect 184716 8260 184772 8270
rect 179116 7476 179172 7486
rect 179116 480 179172 7420
rect 181020 5796 181076 5806
rect 181020 480 181076 5740
rect 182924 4900 182980 4910
rect 182924 480 182980 4844
rect 184716 480 184772 8204
rect 185724 2548 185780 16072
rect 185836 12964 185892 12974
rect 185836 12870 185892 12908
rect 185948 12292 186004 16072
rect 185948 12226 186004 12236
rect 186172 12292 186228 16072
rect 186396 12516 186452 16072
rect 186508 12964 186564 12974
rect 186508 12870 186564 12908
rect 186396 12450 186452 12460
rect 186172 12226 186228 12236
rect 186620 4228 186676 16072
rect 186844 13412 186900 16072
rect 186844 13346 186900 13356
rect 187068 13412 187124 16072
rect 187068 13346 187124 13356
rect 187292 9268 187348 16072
rect 187516 12292 187572 16072
rect 187516 12226 187572 12236
rect 187292 9202 187348 9212
rect 186620 4162 186676 4172
rect 186732 5012 186788 5022
rect 185724 2482 185780 2492
rect 186060 1092 186116 1102
rect 186060 756 186116 1036
rect 186060 690 186116 700
rect 186732 480 186788 4956
rect 187740 4340 187796 16072
rect 187964 5908 188020 16072
rect 188188 10948 188244 16072
rect 188412 13188 188468 16072
rect 188412 13122 188468 13132
rect 188636 12628 188692 16072
rect 188636 12562 188692 12572
rect 188188 10882 188244 10892
rect 187964 5842 188020 5852
rect 188636 9268 188692 9278
rect 187740 4274 187796 4284
rect 188636 480 188692 9212
rect 165564 392 165816 480
rect 167468 392 167720 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 392 169652 480
rect 171304 392 171556 480
rect 173208 392 173460 480
rect 175112 392 175364 480
rect 177016 392 177268 480
rect 178920 392 179172 480
rect 180824 392 181076 480
rect 182728 392 182980 480
rect 169400 -960 169624 392
rect 171304 -960 171528 392
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 480
rect 186536 392 186788 480
rect 188440 392 188692 480
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 188860 84 188916 16072
rect 189084 12292 189140 16072
rect 189308 14308 189364 16072
rect 189308 14242 189364 14252
rect 189084 12226 189140 12236
rect 189308 12180 189364 12190
rect 189308 2660 189364 12124
rect 189532 4452 189588 16072
rect 189756 8428 189812 16072
rect 189980 11060 190036 16072
rect 190204 13188 190260 16072
rect 190204 13122 190260 13132
rect 190428 12740 190484 16072
rect 190652 13412 190708 16072
rect 190652 13346 190708 13356
rect 190428 12674 190484 12684
rect 190652 12740 190708 12750
rect 189980 10994 190036 11004
rect 189532 4386 189588 4396
rect 189644 8372 189812 8428
rect 190540 10948 190596 10958
rect 189308 2594 189364 2604
rect 189644 196 189700 8372
rect 190540 480 190596 10892
rect 190652 10836 190708 12684
rect 190876 12292 190932 16072
rect 190876 12226 190932 12236
rect 191100 12180 191156 16072
rect 191100 12114 191156 12124
rect 190652 10770 190708 10780
rect 189644 130 189700 140
rect 190344 392 190596 480
rect 188860 18 188916 28
rect 190344 -960 190568 392
rect 191324 308 191380 16072
rect 191436 12292 191492 12302
rect 191436 6132 191492 12236
rect 191548 9380 191604 16072
rect 191772 12964 191828 16072
rect 191772 12898 191828 12908
rect 191548 9314 191604 9324
rect 191436 6066 191492 6076
rect 191996 532 192052 16072
rect 192220 6020 192276 16072
rect 192444 14532 192500 16072
rect 192444 14466 192500 14476
rect 192556 12628 192612 12638
rect 192332 12516 192388 12526
rect 192332 7812 192388 12460
rect 192332 7746 192388 7756
rect 192444 12180 192500 12190
rect 192220 5954 192276 5964
rect 192444 4564 192500 12124
rect 192444 4498 192500 4508
rect 192556 4228 192612 12572
rect 192668 12292 192724 16072
rect 192668 12226 192724 12236
rect 192892 7588 192948 16072
rect 193116 13188 193172 16072
rect 193116 13122 193172 13132
rect 192892 7522 192948 7532
rect 192444 4172 192612 4228
rect 192444 480 192500 4172
rect 193340 756 193396 16072
rect 193452 12292 193508 12302
rect 193452 2772 193508 12236
rect 193564 11172 193620 16072
rect 193788 12180 193844 16072
rect 193788 12114 193844 12124
rect 193564 11106 193620 11116
rect 194012 7700 194068 16072
rect 194012 7634 194068 7644
rect 194124 12852 194180 12862
rect 193452 2706 193508 2716
rect 193340 690 193396 700
rect 191996 466 192052 476
rect 191324 242 191380 252
rect 192248 392 192500 480
rect 194124 480 194180 12796
rect 194236 12516 194292 16072
rect 194460 13076 194516 16072
rect 194684 13412 194740 16072
rect 194684 13346 194740 13356
rect 194460 13010 194516 13020
rect 194236 12450 194292 12460
rect 194908 9492 194964 16072
rect 194908 9426 194964 9436
rect 195132 7924 195188 16072
rect 195132 7858 195188 7868
rect 195356 4676 195412 16072
rect 195580 12292 195636 16072
rect 195580 12226 195636 12236
rect 195804 9604 195860 16072
rect 195804 9538 195860 9548
rect 195356 4610 195412 4620
rect 196028 2884 196084 16072
rect 196140 11060 196196 11070
rect 196140 8428 196196 11004
rect 196252 9604 196308 16072
rect 196252 9548 196420 9604
rect 196140 8372 196308 8428
rect 196028 2818 196084 2828
rect 196252 480 196308 8372
rect 196364 1204 196420 9548
rect 196364 1138 196420 1148
rect 196476 1092 196532 16072
rect 196700 13748 196756 16072
rect 196924 14644 196980 16072
rect 196924 14578 196980 14588
rect 196700 13682 196756 13692
rect 197148 8036 197204 16072
rect 197148 7970 197204 7980
rect 197372 2996 197428 16072
rect 197372 2930 197428 2940
rect 197484 12292 197540 12302
rect 196476 1026 196532 1036
rect 197484 868 197540 12236
rect 197596 9716 197652 16072
rect 200508 16100 200564 16110
rect 197820 16034 197876 16044
rect 197596 9650 197652 9660
rect 198044 6356 198100 16072
rect 198156 15204 198212 15214
rect 198268 15204 198324 16072
rect 198212 15148 198324 15204
rect 198156 15138 198212 15148
rect 198044 6290 198100 6300
rect 198492 6244 198548 16072
rect 198716 6468 198772 16072
rect 198716 6402 198772 6412
rect 198492 6178 198548 6188
rect 197484 802 197540 812
rect 198156 4228 198212 4238
rect 198156 480 198212 4172
rect 198940 3108 198996 16072
rect 199164 12292 199220 16072
rect 199164 12226 199220 12236
rect 199388 6580 199444 16072
rect 199500 11956 199556 11966
rect 199500 9828 199556 11900
rect 199612 11396 199668 16072
rect 199836 12404 199892 16072
rect 200060 14756 200116 16072
rect 200060 14690 200116 14700
rect 199836 12338 199892 12348
rect 200284 11508 200340 16072
rect 217308 16100 217364 16110
rect 200508 16034 200564 16044
rect 200284 11442 200340 11452
rect 199612 11330 199668 11340
rect 200396 10052 200452 10062
rect 199500 9762 199556 9772
rect 200060 9940 200116 9950
rect 199388 6514 199444 6524
rect 198940 3042 198996 3052
rect 200060 480 200116 9884
rect 200396 9716 200452 9996
rect 200396 9650 200452 9660
rect 200732 3220 200788 16072
rect 200956 11284 201012 16072
rect 201180 15316 201236 16072
rect 201180 15250 201236 15260
rect 201404 14868 201460 16072
rect 201404 14802 201460 14812
rect 200956 11218 201012 11228
rect 201292 11732 201348 11742
rect 201292 4788 201348 11676
rect 201628 8148 201684 16072
rect 201852 15876 201908 16072
rect 201852 15810 201908 15820
rect 201628 8082 201684 8092
rect 201964 10052 202020 10062
rect 201292 4722 201348 4732
rect 200732 3154 200788 3164
rect 201964 480 202020 9996
rect 202076 3332 202132 16072
rect 202300 11956 202356 16072
rect 202524 13300 202580 16072
rect 202524 13234 202580 13244
rect 202300 11890 202356 11900
rect 202748 11732 202804 16072
rect 202748 11666 202804 11676
rect 202972 11396 203028 16072
rect 202972 11330 203028 11340
rect 203196 9828 203252 16072
rect 203196 9762 203252 9772
rect 202076 3266 202132 3276
rect 203420 2436 203476 16072
rect 203644 6692 203700 16072
rect 203868 12068 203924 16072
rect 204092 14420 204148 16072
rect 204092 14354 204148 14364
rect 203868 12002 203924 12012
rect 204092 12292 204148 12302
rect 203644 6626 203700 6636
rect 203868 8484 203924 8494
rect 203420 2370 203476 2380
rect 203868 480 203924 8428
rect 204092 7476 204148 12236
rect 204316 9828 204372 16072
rect 204540 12740 204596 16072
rect 204540 12674 204596 12684
rect 204316 9762 204372 9772
rect 204764 8372 204820 16072
rect 204988 11508 205044 16072
rect 204988 11442 205044 11452
rect 205212 9156 205268 16072
rect 205436 12292 205492 16072
rect 205436 12226 205492 12236
rect 205548 13300 205604 13310
rect 205212 9090 205268 9100
rect 204764 8306 204820 8316
rect 204092 7410 204148 7420
rect 194124 392 194376 480
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 392 196308 480
rect 197960 392 198212 480
rect 199864 392 200116 480
rect 201768 392 202020 480
rect 203672 392 203924 480
rect 205548 480 205604 13244
rect 205660 5796 205716 16072
rect 205660 5730 205716 5740
rect 205884 4900 205940 16072
rect 206108 8260 206164 16072
rect 206108 8194 206164 8204
rect 206332 5012 206388 16072
rect 206556 9268 206612 16072
rect 206780 10948 206836 16072
rect 207004 12628 207060 16072
rect 207228 12852 207284 16072
rect 207228 12786 207284 12796
rect 207004 12562 207060 12572
rect 207452 11060 207508 16072
rect 207452 10994 207508 11004
rect 207564 13412 207620 13422
rect 206780 10882 206836 10892
rect 206556 9202 206612 9212
rect 206332 4946 206388 4956
rect 205884 4834 205940 4844
rect 207564 480 207620 13356
rect 207676 4228 207732 16072
rect 207900 9940 207956 16072
rect 208124 10052 208180 16072
rect 208124 9986 208180 9996
rect 207900 9874 207956 9884
rect 208348 8484 208404 16072
rect 208572 13300 208628 16072
rect 208796 13412 208852 16072
rect 208796 13346 208852 13356
rect 208572 13234 208628 13244
rect 208348 8418 208404 8428
rect 209020 8428 209076 16072
rect 209020 8372 209188 8428
rect 209132 4228 209188 8372
rect 209244 4452 209300 16072
rect 209468 13412 209524 16072
rect 209468 13346 209524 13356
rect 209692 13412 209748 16072
rect 209692 13346 209748 13356
rect 209916 13412 209972 16072
rect 209916 13346 209972 13356
rect 210140 13412 210196 16072
rect 210140 13346 210196 13356
rect 209244 4386 209300 4396
rect 210364 4228 210420 16072
rect 210588 6804 210644 16072
rect 210588 6738 210644 6748
rect 210812 4340 210868 16072
rect 211036 11620 211092 16072
rect 211036 11554 211092 11564
rect 211260 9380 211316 16072
rect 211260 9314 211316 9324
rect 211484 6468 211540 16072
rect 211484 6402 211540 6412
rect 211708 6132 211764 16072
rect 211932 12852 211988 16072
rect 211932 12786 211988 12796
rect 212156 12740 212212 16072
rect 212156 12674 212212 12684
rect 212380 11508 212436 16072
rect 212380 11442 212436 11452
rect 212604 9268 212660 16072
rect 212604 9202 212660 9212
rect 211708 6066 211764 6076
rect 210812 4274 210868 4284
rect 211260 4452 211316 4462
rect 209132 4172 209412 4228
rect 207676 4162 207732 4172
rect 209356 480 209412 4172
rect 210364 4162 210420 4172
rect 211260 480 211316 4396
rect 212828 4452 212884 16072
rect 212828 4386 212884 4396
rect 213052 4116 213108 16072
rect 213276 8148 213332 16072
rect 213500 11732 213556 16072
rect 213500 11666 213556 11676
rect 213276 8082 213332 8092
rect 213724 7588 213780 16072
rect 213948 8260 214004 16072
rect 213948 8194 214004 8204
rect 214172 7812 214228 16072
rect 214172 7746 214228 7756
rect 213724 7522 213780 7532
rect 214396 6356 214452 16072
rect 214620 15540 214676 16072
rect 214620 15474 214676 15484
rect 214396 6290 214452 6300
rect 214844 5908 214900 16072
rect 215068 12068 215124 16072
rect 215292 15652 215348 16072
rect 215292 15586 215348 15596
rect 215068 12002 215124 12012
rect 215516 7700 215572 16072
rect 215740 14308 215796 16072
rect 215964 15876 216020 16072
rect 215964 15810 216020 15820
rect 215740 14242 215796 14252
rect 216188 9716 216244 16072
rect 216412 13412 216468 16072
rect 216412 13346 216468 13356
rect 217084 13300 217140 16072
rect 219772 16100 219828 16110
rect 217308 16034 217364 16044
rect 217084 13234 217140 13244
rect 216188 9650 216244 9660
rect 216748 11732 216804 11742
rect 215516 7634 215572 7644
rect 214844 5842 214900 5852
rect 215068 6804 215124 6814
rect 213052 4050 213108 4060
rect 213164 4228 213220 4238
rect 213164 480 213220 4172
rect 215068 480 215124 6748
rect 216748 4676 216804 11676
rect 217756 11396 217812 16072
rect 217756 11330 217812 11340
rect 217980 6244 218036 16072
rect 218204 10164 218260 16072
rect 218428 10836 218484 16072
rect 218652 13412 218708 16072
rect 218876 14532 218932 16072
rect 218876 14466 218932 14476
rect 218652 13346 218708 13356
rect 218428 10770 218484 10780
rect 218876 11620 218932 11630
rect 218204 10098 218260 10108
rect 217980 6178 218036 6188
rect 216748 4610 216804 4620
rect 216972 4340 217028 4350
rect 216972 480 217028 4284
rect 218876 480 218932 11564
rect 219324 2660 219380 16072
rect 219548 6020 219604 16072
rect 226044 16100 226100 16110
rect 219772 16034 219828 16044
rect 219996 14980 220052 16072
rect 219996 14914 220052 14924
rect 220220 10500 220276 16072
rect 220444 13188 220500 16072
rect 220444 13122 220500 13132
rect 220668 12628 220724 16072
rect 220668 12562 220724 12572
rect 220892 12516 220948 16072
rect 221340 14980 221396 16072
rect 221340 14914 221396 14924
rect 220892 12450 220948 12460
rect 221564 10948 221620 16072
rect 221564 10882 221620 10892
rect 220220 10434 220276 10444
rect 219548 5954 219604 5964
rect 220780 9380 220836 9390
rect 219324 2594 219380 2604
rect 220780 480 220836 9324
rect 221788 3332 221844 16072
rect 222012 12964 222068 16072
rect 222236 14980 222292 16072
rect 222236 14914 222292 14924
rect 222012 12898 222068 12908
rect 222684 8372 222740 16072
rect 223356 12292 223412 16072
rect 223356 12226 223412 12236
rect 222684 8306 222740 8316
rect 221788 3266 221844 3276
rect 222684 6468 222740 6478
rect 222684 480 222740 6412
rect 223580 2324 223636 16072
rect 223804 11172 223860 16072
rect 224028 12404 224084 16072
rect 224028 12338 224084 12348
rect 223804 11106 223860 11116
rect 224252 9604 224308 16072
rect 224476 13412 224532 16072
rect 224476 13346 224532 13356
rect 224700 12292 224756 16072
rect 224700 12226 224756 12236
rect 224252 9538 224308 9548
rect 224924 9492 224980 16072
rect 224924 9426 224980 9436
rect 223580 2258 223636 2268
rect 224588 6132 224644 6142
rect 224588 480 224644 6076
rect 225148 3220 225204 16072
rect 225372 12404 225428 16072
rect 225372 12338 225428 12348
rect 225596 9380 225652 16072
rect 226044 16034 226100 16044
rect 226492 15764 226548 16072
rect 226492 15698 226548 15708
rect 225596 9314 225652 9324
rect 226492 12852 226548 12862
rect 225148 3154 225204 3164
rect 226492 480 226548 12796
rect 226716 12292 226772 16072
rect 226828 15428 226884 15438
rect 226828 13188 226884 15372
rect 226828 13122 226884 13132
rect 226716 12226 226772 12236
rect 226940 8036 226996 16072
rect 227164 15204 227220 16072
rect 227164 15138 227220 15148
rect 227388 12852 227444 16072
rect 227388 12786 227444 12796
rect 226940 7970 226996 7980
rect 227612 6132 227668 16072
rect 227836 11060 227892 16072
rect 228060 12292 228116 16072
rect 228060 12226 228116 12236
rect 228284 12180 228340 16072
rect 228508 14420 228564 16072
rect 228508 14354 228564 14364
rect 228284 12114 228340 12124
rect 228508 12740 228564 12750
rect 227836 10994 227892 11004
rect 227612 6066 227668 6076
rect 226828 5908 226884 5918
rect 226828 4564 226884 5852
rect 226828 4498 226884 4508
rect 228508 480 228564 12684
rect 228620 7812 228676 7822
rect 228620 4004 228676 7756
rect 228732 6692 228788 16072
rect 228956 11284 229012 16072
rect 229180 11732 229236 16072
rect 229404 12292 229460 16072
rect 229404 12226 229460 12236
rect 229180 11666 229236 11676
rect 228956 11218 229012 11228
rect 229628 7924 229684 16072
rect 229628 7858 229684 7868
rect 228732 6626 228788 6636
rect 228620 3938 228676 3948
rect 229852 2436 229908 16072
rect 230076 10052 230132 16072
rect 230188 13636 230244 13646
rect 230188 13300 230244 13580
rect 230188 13234 230244 13244
rect 230076 9986 230132 9996
rect 230188 11508 230244 11518
rect 230188 8428 230244 11452
rect 230300 9604 230356 16072
rect 230412 15316 230468 15326
rect 230412 13412 230468 15260
rect 230412 13346 230468 13356
rect 230300 9548 230468 9604
rect 230188 8372 230356 8428
rect 230188 6356 230244 6366
rect 230188 4116 230244 6300
rect 230188 4050 230244 4060
rect 229852 2370 229908 2380
rect 230188 3332 230244 3342
rect 230188 1092 230244 3276
rect 230188 1026 230244 1036
rect 230300 480 230356 8372
rect 230412 7812 230468 9548
rect 230412 7746 230468 7756
rect 230524 1316 230580 16072
rect 230972 5908 231028 16072
rect 231420 12740 231476 16072
rect 231420 12674 231476 12684
rect 231644 12292 231700 16072
rect 231644 12226 231700 12236
rect 231868 8428 231924 16072
rect 232092 12740 232148 16072
rect 232092 12674 232148 12684
rect 232204 9268 232260 9278
rect 231868 8372 232148 8428
rect 230972 5842 231028 5852
rect 230524 1250 230580 1260
rect 232092 644 232148 8372
rect 232092 578 232148 588
rect 232204 480 232260 9212
rect 232316 3108 232372 16072
rect 232540 12404 232596 16072
rect 232540 12338 232596 12348
rect 232316 3042 232372 3052
rect 232764 1652 232820 16072
rect 232988 12292 233044 16072
rect 232988 12226 233044 12236
rect 233212 2100 233268 16072
rect 233436 14084 233492 16072
rect 233324 14028 233492 14084
rect 233324 11732 233380 14028
rect 233436 13860 233492 13870
rect 233436 12068 233492 13804
rect 233436 12002 233492 12012
rect 233324 11666 233380 11676
rect 233436 7700 233492 7710
rect 233436 4452 233492 7644
rect 233436 4386 233492 4396
rect 233212 2034 233268 2044
rect 232764 1586 232820 1596
rect 233660 1540 233716 16072
rect 233884 14644 233940 16072
rect 233884 14578 233940 14588
rect 234108 8428 234164 16072
rect 234108 8372 234276 8428
rect 233660 1474 233716 1484
rect 234108 4340 234164 4350
rect 234108 480 234164 4284
rect 234220 2884 234276 8372
rect 234332 7700 234388 16072
rect 234332 7634 234388 7644
rect 234220 2818 234276 2828
rect 234556 1428 234612 16072
rect 234780 13188 234836 16072
rect 234780 13122 234836 13132
rect 234892 12740 234948 12750
rect 234892 9268 234948 12684
rect 234892 9202 234948 9212
rect 235004 3332 235060 16072
rect 235228 13300 235284 16072
rect 235228 13234 235284 13244
rect 235116 12404 235172 12414
rect 235116 9156 235172 12348
rect 235116 9090 235172 9100
rect 235116 7588 235172 7598
rect 235116 4900 235172 7532
rect 235116 4834 235172 4844
rect 235004 3266 235060 3276
rect 234556 1362 234612 1372
rect 235452 1204 235508 16072
rect 235676 7588 235732 16072
rect 235676 7522 235732 7532
rect 235900 2772 235956 16072
rect 236124 13412 236180 16072
rect 236124 13346 236180 13356
rect 235900 2706 235956 2716
rect 236012 4228 236068 4238
rect 235452 1138 235508 1148
rect 236012 480 236068 4172
rect 236348 532 236404 16072
rect 236796 12964 236852 16072
rect 236796 12898 236852 12908
rect 237020 11620 237076 16072
rect 237244 11844 237300 16072
rect 237244 11778 237300 11788
rect 237020 11554 237076 11564
rect 236796 8260 236852 8270
rect 236796 4228 236852 8204
rect 237468 6468 237524 16072
rect 237468 6402 237524 6412
rect 236796 4162 236852 4172
rect 237692 644 237748 16072
rect 237916 12404 237972 16072
rect 237916 12338 237972 12348
rect 237804 12292 237860 12302
rect 237804 6580 237860 12236
rect 238140 12068 238196 16072
rect 238364 12292 238420 16072
rect 238364 12226 238420 12236
rect 238140 12002 238196 12012
rect 238812 11844 238868 16072
rect 239036 12740 239092 16072
rect 239036 12674 239092 12684
rect 238812 11778 238868 11788
rect 238476 9716 238532 9726
rect 237804 6514 237860 6524
rect 237916 8148 237972 8158
rect 237692 578 237748 588
rect 205548 392 205800 480
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 392
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 -960 205800 392
rect 207480 -960 207704 480
rect 209356 392 209608 480
rect 211260 392 211512 480
rect 213164 392 213416 480
rect 215068 392 215320 480
rect 216972 392 217224 480
rect 218876 392 219128 480
rect 220780 392 221032 480
rect 222684 392 222936 480
rect 224588 392 224840 480
rect 226492 392 226744 480
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 392
rect 215096 -960 215320 392
rect 217000 -960 217224 392
rect 218904 -960 219128 392
rect 220808 -960 221032 392
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230300 392 230552 480
rect 232204 392 232456 480
rect 234108 392 234360 480
rect 236012 392 236264 480
rect 236348 466 236404 476
rect 237916 480 237972 8092
rect 238476 4788 238532 9660
rect 239484 5012 239540 16072
rect 239708 9940 239764 16072
rect 240156 12292 240212 16072
rect 240268 13748 240324 13758
rect 240268 12516 240324 13692
rect 240268 12450 240324 12460
rect 240492 12964 240548 12974
rect 240492 12516 240548 12908
rect 240828 12964 240884 16072
rect 240828 12898 240884 12908
rect 240492 12450 240548 12460
rect 240156 12226 240212 12236
rect 239708 9874 239764 9884
rect 241052 8260 241108 16072
rect 241276 12292 241332 16072
rect 241500 13412 241556 16072
rect 241500 13346 241556 13356
rect 241276 12226 241332 12236
rect 241724 9716 241780 16072
rect 241724 9650 241780 9660
rect 241052 8194 241108 8204
rect 239484 4946 239540 4956
rect 238476 4722 238532 4732
rect 241724 4900 241780 4910
rect 239820 4676 239876 4686
rect 239820 480 239876 4620
rect 241724 480 241780 4844
rect 241948 4900 242004 16072
rect 242172 12404 242228 16072
rect 242396 12852 242452 16072
rect 242396 12786 242452 12796
rect 242172 12338 242228 12348
rect 242620 11844 242676 16072
rect 242620 11778 242676 11788
rect 241948 4834 242004 4844
rect 242844 4340 242900 16072
rect 243068 14980 243124 16072
rect 243068 14914 243124 14924
rect 243292 13412 243348 16072
rect 243292 13346 243348 13356
rect 243292 12180 243348 12190
rect 243516 12180 243572 16072
rect 243348 12124 243572 12180
rect 243292 12114 243348 12124
rect 243964 4788 244020 16072
rect 244188 12852 244244 16072
rect 244188 12786 244244 12796
rect 244412 12404 244468 16072
rect 244412 12338 244468 12348
rect 244524 14644 244580 14654
rect 244412 12180 244468 12190
rect 244412 11956 244468 12124
rect 244412 11890 244468 11900
rect 244524 6356 244580 14588
rect 244636 12180 244692 16072
rect 244860 14980 244916 16072
rect 244860 14914 244916 14924
rect 244636 12114 244692 12124
rect 245532 12180 245588 16072
rect 245532 12114 245588 12124
rect 245756 8148 245812 16072
rect 245980 13412 246036 16072
rect 245980 13346 246036 13356
rect 247772 15428 247828 15438
rect 245756 8082 245812 8092
rect 244524 6290 244580 6300
rect 243964 4722 244020 4732
rect 242844 4274 242900 4284
rect 243628 4228 243684 4238
rect 243628 480 243684 4172
rect 247436 4116 247492 4126
rect 245532 4004 245588 4014
rect 245532 480 245588 3948
rect 247436 480 247492 4060
rect 247772 980 247828 15372
rect 248556 11956 248612 16156
rect 248556 11890 248612 11900
rect 249228 15540 249284 15550
rect 249228 8428 249284 15484
rect 249452 13300 249508 13310
rect 249452 12516 249508 13244
rect 249452 12450 249508 12460
rect 249340 11508 249396 11518
rect 249340 8932 249396 11452
rect 249452 10164 249508 10174
rect 249452 9156 249508 10108
rect 249452 9090 249508 9100
rect 249340 8866 249396 8876
rect 249228 8372 249396 8428
rect 248556 3668 248612 3678
rect 248556 3220 248612 3612
rect 248556 3154 248612 3164
rect 247772 914 247828 924
rect 248668 1316 248724 1326
rect 237916 392 238168 480
rect 239820 392 240072 480
rect 241724 392 241976 480
rect 243628 392 243880 480
rect 245532 392 245784 480
rect 247436 392 247688 480
rect 230328 -960 230552 392
rect 232232 -960 232456 392
rect 234136 -960 234360 392
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 239848 -960 240072 392
rect 241752 -960 241976 392
rect 243656 -960 243880 392
rect 245560 -960 245784 392
rect 247464 -960 247688 392
rect 248668 420 248724 1260
rect 249340 480 249396 8372
rect 249564 1204 249620 16268
rect 260764 15876 260820 15886
rect 255052 15652 255108 15662
rect 253708 15428 253764 15438
rect 253708 15092 253764 15372
rect 253708 15026 253764 15036
rect 253148 13860 253204 13870
rect 251916 11396 251972 11406
rect 249564 1138 249620 1148
rect 251244 4564 251300 4574
rect 251244 480 251300 4508
rect 251916 4116 251972 11340
rect 251916 4050 251972 4060
rect 253148 480 253204 13804
rect 255052 480 255108 15596
rect 258860 14308 258916 14318
rect 257068 8932 257124 8942
rect 257068 4676 257124 8876
rect 257068 4610 257124 4620
rect 257068 4452 257124 4462
rect 257068 480 257124 4396
rect 258860 480 258916 14252
rect 260764 480 260820 15820
rect 264572 13524 264628 13534
rect 264460 10164 264516 10174
rect 262668 4340 262724 4350
rect 262668 480 262724 4284
rect 264460 2996 264516 10108
rect 264460 2930 264516 2940
rect 264572 480 264628 13468
rect 265244 3108 265300 18508
rect 265468 15316 265524 15326
rect 265468 13412 265524 15260
rect 265468 13346 265524 13356
rect 265692 15092 265748 15102
rect 265468 11172 265524 11182
rect 265468 8260 265524 11116
rect 265692 11172 265748 15036
rect 266252 13188 266308 100828
rect 268156 96516 268212 96526
rect 266252 13122 266308 13132
rect 266364 94500 266420 94510
rect 265692 11106 265748 11116
rect 266364 9940 266420 94444
rect 266700 90916 266756 90926
rect 266588 81060 266644 81070
rect 266364 9874 266420 9884
rect 266476 16100 266532 16110
rect 265468 8194 265524 8204
rect 265804 8036 265860 8046
rect 265468 5124 265524 5134
rect 265468 4788 265524 5068
rect 265468 4722 265524 4732
rect 265692 4676 265748 4686
rect 265244 3042 265300 3052
rect 265580 3444 265636 3454
rect 265468 2548 265524 2558
rect 265468 980 265524 2492
rect 265580 2436 265636 3388
rect 265580 2370 265636 2380
rect 265692 2212 265748 4620
rect 265804 3108 265860 7980
rect 265804 3042 265860 3052
rect 265692 2146 265748 2156
rect 265468 914 265524 924
rect 266476 480 266532 16044
rect 266588 2884 266644 81004
rect 266700 8372 266756 90860
rect 266924 85316 266980 85326
rect 266700 8306 266756 8316
rect 266812 76356 266868 76366
rect 266812 6468 266868 76300
rect 266924 14980 266980 85260
rect 268156 83860 268212 96460
rect 269612 96068 269668 96078
rect 268156 83794 268212 83804
rect 268828 85764 268884 85774
rect 267932 83300 267988 83310
rect 267932 83076 267988 83244
rect 267932 83010 267988 83020
rect 268268 80836 268324 80846
rect 268156 78932 268212 78942
rect 266924 14914 266980 14924
rect 267036 78372 267092 78382
rect 267036 11620 267092 78316
rect 267932 78148 267988 78158
rect 267036 11554 267092 11564
rect 267820 13412 267876 13422
rect 266812 6402 266868 6412
rect 267820 4564 267876 13356
rect 267820 4498 267876 4508
rect 266588 2818 266644 2828
rect 267932 1540 267988 78092
rect 268044 77252 268100 77262
rect 268044 4900 268100 77196
rect 268044 4834 268100 4844
rect 268156 2772 268212 78876
rect 268268 13300 268324 80780
rect 268604 78596 268660 78606
rect 268268 13234 268324 13244
rect 268380 17108 268436 17118
rect 268156 2706 268212 2716
rect 267932 1474 267988 1484
rect 268380 480 268436 17052
rect 268604 16884 268660 78540
rect 268828 18452 268884 85708
rect 268828 18386 268884 18396
rect 268940 82404 268996 82414
rect 268940 18340 268996 82348
rect 268940 18274 268996 18284
rect 269500 17332 269556 17342
rect 268604 16818 268660 16828
rect 269388 17220 269444 17230
rect 269276 15988 269332 15998
rect 269164 15428 269220 15438
rect 268716 14644 268772 14654
rect 268492 13412 268548 13422
rect 268492 1428 268548 13356
rect 268716 13300 268772 14588
rect 268716 13234 268772 13244
rect 268716 12964 268772 12974
rect 268716 11732 268772 12908
rect 268716 11666 268772 11676
rect 268940 10948 268996 10958
rect 268940 6580 268996 10892
rect 269164 9156 269220 15372
rect 269164 9090 269220 9100
rect 269276 8148 269332 15932
rect 269388 9940 269444 17164
rect 269388 9874 269444 9884
rect 269276 8082 269332 8092
rect 269500 8036 269556 17276
rect 269612 13412 269668 96012
rect 272972 93492 273028 305340
rect 273084 305060 273140 308056
rect 273084 304994 273140 305004
rect 273084 218484 273140 218494
rect 273084 96516 273140 218428
rect 273084 96450 273140 96460
rect 273532 94948 273588 308056
rect 273980 305284 274036 308056
rect 273980 305218 274036 305228
rect 273532 94882 273588 94892
rect 273868 305172 273924 305182
rect 272972 93426 273028 93436
rect 273756 93492 273812 93502
rect 271292 91140 271348 91150
rect 269724 86100 269780 86110
rect 269724 16212 269780 86044
rect 270620 84532 270676 84542
rect 269836 84308 269892 84318
rect 269836 18564 269892 84252
rect 270284 84196 270340 84206
rect 270284 23156 270340 84140
rect 270620 77140 270676 84476
rect 271180 83300 271236 83310
rect 271180 78596 271236 83244
rect 271292 78932 271348 91084
rect 273756 87108 273812 93436
rect 273868 93380 273924 305116
rect 273868 93314 273924 93324
rect 273756 87042 273812 87052
rect 274428 83188 274484 308056
rect 274652 231028 274708 231038
rect 274652 218484 274708 230972
rect 274652 218418 274708 218428
rect 274876 98532 274932 308056
rect 275324 101668 275380 308056
rect 275324 101602 275380 101612
rect 275772 100548 275828 308056
rect 275772 100482 275828 100492
rect 274876 98466 274932 98476
rect 276220 91588 276276 308056
rect 276220 91522 276276 91532
rect 276332 91028 276388 91038
rect 276332 85316 276388 90972
rect 276332 85250 276388 85260
rect 274428 83122 274484 83132
rect 274652 83860 274708 83870
rect 271292 78866 271348 78876
rect 271180 78530 271236 78540
rect 274652 78484 274708 83804
rect 276668 83188 276724 308056
rect 277116 101780 277172 308056
rect 277116 101714 277172 101724
rect 277228 305508 277284 305518
rect 277228 100212 277284 305452
rect 277564 305396 277620 308056
rect 277564 305330 277620 305340
rect 277228 100146 277284 100156
rect 278012 91700 278068 308056
rect 278348 304948 278404 304958
rect 278012 91634 278068 91644
rect 278124 304388 278180 304398
rect 276668 83122 276724 83132
rect 278124 81508 278180 304332
rect 278348 96852 278404 304892
rect 278460 101892 278516 308056
rect 278460 101826 278516 101836
rect 278348 96786 278404 96796
rect 278908 95172 278964 308056
rect 279020 245252 279076 245262
rect 279020 236852 279076 245196
rect 279020 236786 279076 236796
rect 278908 95106 278964 95116
rect 279356 91812 279412 308056
rect 279804 91924 279860 308056
rect 280252 98420 280308 308056
rect 280252 98354 280308 98364
rect 279804 91858 279860 91868
rect 279356 91746 279412 91756
rect 280700 89908 280756 308056
rect 281148 304388 281204 308056
rect 281148 304322 281204 304332
rect 281372 305172 281428 305182
rect 281372 102004 281428 305116
rect 281372 101938 281428 101948
rect 280700 89842 280756 89852
rect 281596 86548 281652 308056
rect 282044 98644 282100 308056
rect 282492 304948 282548 308056
rect 282604 308028 282968 308084
rect 282604 305284 282660 308028
rect 282604 305218 282660 305228
rect 283052 305396 283108 305406
rect 282492 304882 282548 304892
rect 282044 98578 282100 98588
rect 283052 96964 283108 305340
rect 283052 96898 283108 96908
rect 283388 90020 283444 308056
rect 283836 305172 283892 308056
rect 283836 305106 283892 305116
rect 283388 89954 283444 89964
rect 284284 86660 284340 308056
rect 284732 305508 284788 308056
rect 284732 305442 284788 305452
rect 284732 305284 284788 305294
rect 284732 86772 284788 305228
rect 284956 305172 285012 305182
rect 284956 88228 285012 305116
rect 285180 92036 285236 308056
rect 285628 305284 285684 308056
rect 286104 308028 286356 308084
rect 285628 305218 285684 305228
rect 285740 305508 285796 305518
rect 285292 304948 285348 304958
rect 285292 93716 285348 304892
rect 285628 251972 285684 251982
rect 285628 245252 285684 251916
rect 285628 245186 285684 245196
rect 285740 100324 285796 305452
rect 286300 305284 286356 308028
rect 286300 305218 286356 305228
rect 286524 305172 286580 308056
rect 286972 305396 287028 308056
rect 286972 305330 287028 305340
rect 286524 305106 286580 305116
rect 286412 250292 286468 250302
rect 286412 231028 286468 250236
rect 286412 230962 286468 230972
rect 285740 100258 285796 100268
rect 285292 93650 285348 93660
rect 286412 96068 286468 96078
rect 285180 91970 285236 91980
rect 286412 89908 286468 96012
rect 287420 90244 287476 308056
rect 287420 90178 287476 90188
rect 286412 89842 286468 89852
rect 284956 88162 285012 88172
rect 284732 86706 284788 86716
rect 287308 87444 287364 87454
rect 284284 86594 284340 86604
rect 281596 86482 281652 86492
rect 282156 84420 282212 84430
rect 282156 83300 282212 84364
rect 287308 83972 287364 87388
rect 287868 86996 287924 308056
rect 287868 86930 287924 86940
rect 287308 83906 287364 83916
rect 282156 83234 282212 83244
rect 278124 81442 278180 81452
rect 282156 82516 282212 82526
rect 282156 79604 282212 82460
rect 288316 81620 288372 308056
rect 288764 90132 288820 308056
rect 289212 90692 289268 308056
rect 289660 101556 289716 308056
rect 289660 101490 289716 101500
rect 290108 98756 290164 308056
rect 290108 98690 290164 98700
rect 290556 92148 290612 308056
rect 290556 92082 290612 92092
rect 289212 90626 289268 90636
rect 288764 90066 288820 90076
rect 291004 83412 291060 308056
rect 291452 305284 291508 308056
rect 291452 305218 291508 305228
rect 291452 268772 291508 268782
rect 291452 250292 291508 268716
rect 291676 268660 291732 268670
rect 291676 251972 291732 268604
rect 291676 251906 291732 251916
rect 291452 250226 291508 250236
rect 291900 90356 291956 308056
rect 292348 100436 292404 308056
rect 292796 305284 292852 308056
rect 292796 305218 292852 305228
rect 292348 100370 292404 100380
rect 293244 90468 293300 308056
rect 293692 98868 293748 308056
rect 294140 305284 294196 308056
rect 294140 305218 294196 305228
rect 293692 98802 293748 98812
rect 294588 90580 294644 308056
rect 295036 93604 295092 308056
rect 295036 93538 295092 93548
rect 294588 90514 294644 90524
rect 293244 90402 293300 90412
rect 291900 90290 291956 90300
rect 295484 88452 295540 308056
rect 295932 304948 295988 308056
rect 295932 304882 295988 304892
rect 296380 97076 296436 308056
rect 296380 97010 296436 97020
rect 295484 88386 295540 88396
rect 296828 88340 296884 308056
rect 297276 95284 297332 308056
rect 297388 273924 297444 273934
rect 297388 268660 297444 273868
rect 297388 268594 297444 268604
rect 297276 95218 297332 95228
rect 296828 88274 296884 88284
rect 295596 88116 295652 88126
rect 291004 83346 291060 83356
rect 292236 86212 292292 86222
rect 288316 81554 288372 81564
rect 282156 79538 282212 79548
rect 287196 81508 287252 81518
rect 274652 78418 274708 78428
rect 287196 78372 287252 81452
rect 292236 80500 292292 86156
rect 295596 81844 295652 88060
rect 297724 84868 297780 308056
rect 298172 86884 298228 308056
rect 298172 86818 298228 86828
rect 298284 305172 298340 305182
rect 297724 84802 297780 84812
rect 298284 83636 298340 305116
rect 298284 83570 298340 83580
rect 295596 81778 295652 81788
rect 298620 81732 298676 308056
rect 299068 305396 299124 308056
rect 299068 305330 299124 305340
rect 299516 305284 299572 308056
rect 299516 305218 299572 305228
rect 298956 91140 299012 91150
rect 298956 84868 299012 91084
rect 299068 87444 299124 87454
rect 299068 85316 299124 87388
rect 299068 85250 299124 85260
rect 299180 85764 299236 85774
rect 298956 84802 299012 84812
rect 299180 83188 299236 85708
rect 299964 84980 300020 308056
rect 300412 85092 300468 308056
rect 300860 305172 300916 308056
rect 300860 305106 300916 305116
rect 300748 271348 300804 271358
rect 300748 268772 300804 271292
rect 300748 268706 300804 268716
rect 301308 85204 301364 308056
rect 301532 291508 301588 291518
rect 301532 273924 301588 291452
rect 301532 273858 301588 273868
rect 301308 85138 301364 85148
rect 300412 85026 300468 85036
rect 299964 84914 300020 84924
rect 301756 83524 301812 308056
rect 302204 101444 302260 308056
rect 302652 304948 302708 308056
rect 302652 304882 302708 304892
rect 303100 301700 303156 308056
rect 303548 303492 303604 308056
rect 303996 304052 304052 308056
rect 303996 303986 304052 303996
rect 304444 303716 304500 308056
rect 304892 306740 304948 308056
rect 304892 306674 304948 306684
rect 305340 306628 305396 308056
rect 305340 306562 305396 306572
rect 304444 303650 304500 303660
rect 303548 303426 303604 303436
rect 305788 303268 305844 308056
rect 305788 303202 305844 303212
rect 303100 301634 303156 301644
rect 306236 301588 306292 308056
rect 306684 305284 306740 308056
rect 306684 305218 306740 305228
rect 307132 305172 307188 308056
rect 307580 305396 307636 308056
rect 308028 305508 308084 308056
rect 308476 305732 308532 308056
rect 308476 305666 308532 305676
rect 308028 305442 308084 305452
rect 307580 305330 307636 305340
rect 307132 305106 307188 305116
rect 308924 304724 308980 308056
rect 308924 304658 308980 304668
rect 306236 301522 306292 301532
rect 309372 301364 309428 308056
rect 309820 301924 309876 308056
rect 309820 301858 309876 301868
rect 309372 301298 309428 301308
rect 310268 299908 310324 308056
rect 310716 306964 310772 308056
rect 310716 306898 310772 306908
rect 311164 306852 311220 308056
rect 311164 306786 311220 306796
rect 311612 303828 311668 308056
rect 311612 303762 311668 303772
rect 311836 304276 311892 304286
rect 310268 299842 310324 299852
rect 311164 280644 311220 280654
rect 311164 271348 311220 280588
rect 311164 271282 311220 271292
rect 302204 101378 302260 101388
rect 309148 94948 309204 94958
rect 309148 93492 309204 94892
rect 309148 93426 309204 93436
rect 311836 90020 311892 304220
rect 312060 303604 312116 308056
rect 312508 303940 312564 308056
rect 312508 303874 312564 303884
rect 312060 303538 312116 303548
rect 312956 301812 313012 308056
rect 313404 305620 313460 308056
rect 313404 305554 313460 305564
rect 312956 301746 313012 301756
rect 313852 300468 313908 308056
rect 314300 304836 314356 308056
rect 314300 304770 314356 304780
rect 314748 302260 314804 308056
rect 315196 304612 315252 308056
rect 315196 304546 315252 304556
rect 315084 304164 315140 304174
rect 314748 302194 314804 302204
rect 314972 302708 315028 302718
rect 313852 300402 313908 300412
rect 312508 296660 312564 296670
rect 312508 291508 312564 296604
rect 312508 291442 312564 291452
rect 311836 89954 311892 89964
rect 314972 86548 315028 302652
rect 315084 91588 315140 304108
rect 315644 303380 315700 308056
rect 316092 307412 316148 308056
rect 316092 307346 316148 307356
rect 316540 306516 316596 308056
rect 316540 306450 316596 306460
rect 315644 303314 315700 303324
rect 315084 91522 315140 91532
rect 315196 301028 315252 301038
rect 315196 87108 315252 300972
rect 316988 300132 317044 308056
rect 316988 300066 317044 300076
rect 317436 298116 317492 308056
rect 317884 307188 317940 308056
rect 317884 307122 317940 307132
rect 318332 304052 318388 308056
rect 318332 303986 318388 303996
rect 318444 305844 318500 305854
rect 317436 298050 317492 298060
rect 318332 302596 318388 302606
rect 316652 296772 316708 296782
rect 316652 280644 316708 296716
rect 316652 280578 316708 280588
rect 315196 87042 315252 87052
rect 315644 88004 315700 88014
rect 314972 86482 315028 86492
rect 315644 84980 315700 87948
rect 318332 86772 318388 302540
rect 318444 91700 318500 305788
rect 318444 91634 318500 91644
rect 318556 302484 318612 302494
rect 318556 86996 318612 302428
rect 318780 300020 318836 308056
rect 319228 303380 319284 308056
rect 319676 305284 319732 308056
rect 319676 305218 319732 305228
rect 320124 305284 320180 308056
rect 320124 305218 320180 305228
rect 319228 303314 319284 303324
rect 320572 302036 320628 308056
rect 321020 302484 321076 308056
rect 321020 302418 321076 302428
rect 321468 302148 321524 308056
rect 321916 307076 321972 308056
rect 322364 307300 322420 308056
rect 322364 307234 322420 307244
rect 321916 307010 321972 307020
rect 321468 302082 321524 302092
rect 320572 301970 320628 301980
rect 318780 299954 318836 299964
rect 318892 300916 318948 300926
rect 318668 298004 318724 298014
rect 318668 90356 318724 297948
rect 318668 90290 318724 90300
rect 318556 86930 318612 86940
rect 318892 86884 318948 300860
rect 322812 300356 322868 308056
rect 322812 300290 322868 300300
rect 323148 304948 323204 304958
rect 323148 298872 323204 304892
rect 323260 303156 323316 308056
rect 323260 303090 323316 303100
rect 323484 305284 323540 305294
rect 323484 301476 323540 305228
rect 323708 304388 323764 308056
rect 324156 305732 324212 308056
rect 324156 305666 324212 305676
rect 324604 305732 324660 308056
rect 324604 305666 324660 305676
rect 325052 304948 325108 308056
rect 325052 304882 325108 304892
rect 325388 306740 325444 306750
rect 323708 304322 323764 304332
rect 324940 303716 324996 303726
rect 324044 303492 324100 303502
rect 323484 301410 323540 301420
rect 323596 301700 323652 301710
rect 323596 298872 323652 301644
rect 324044 298872 324100 303436
rect 324492 302820 324548 302830
rect 324492 298872 324548 302764
rect 324940 298872 324996 303660
rect 325388 298872 325444 306684
rect 325500 304724 325556 308056
rect 325500 304658 325556 304668
rect 325948 304276 326004 308056
rect 325948 304210 326004 304220
rect 326284 306628 326340 306638
rect 325836 301364 325892 301374
rect 325836 298872 325892 301308
rect 326284 298872 326340 306572
rect 326396 304612 326452 308056
rect 326396 304546 326452 304556
rect 326508 304500 326564 304510
rect 326508 300804 326564 304444
rect 326508 300738 326564 300748
rect 326732 303268 326788 303278
rect 326732 298872 326788 303212
rect 326844 301700 326900 308056
rect 327292 305732 327348 308056
rect 327740 306628 327796 308056
rect 327740 306562 327796 306572
rect 327292 305666 327348 305676
rect 327180 305508 327236 305518
rect 327180 303716 327236 305452
rect 327180 303650 327236 303660
rect 327740 304164 327796 304174
rect 327740 302428 327796 304108
rect 328188 303492 328244 308056
rect 328188 303426 328244 303436
rect 328524 303716 328580 303726
rect 326844 301634 326900 301644
rect 327628 302372 327796 302428
rect 328076 302596 328132 302606
rect 327180 301588 327236 301598
rect 327180 298872 327236 301532
rect 327628 298872 327684 302372
rect 328076 298872 328132 302540
rect 328524 298872 328580 303660
rect 328636 303268 328692 308056
rect 329084 305508 329140 308056
rect 329084 305442 329140 305452
rect 328636 303202 328692 303212
rect 328972 300804 329028 300814
rect 328972 298872 329028 300748
rect 329420 300804 329476 300814
rect 329420 298872 329476 300748
rect 329532 300244 329588 308056
rect 329980 306740 330036 308056
rect 329980 306674 330036 306684
rect 330428 305732 330484 308056
rect 330428 305666 330484 305676
rect 330876 304388 330932 308056
rect 330876 304322 330932 304332
rect 331212 306964 331268 306974
rect 330316 301924 330372 301934
rect 329532 300178 329588 300188
rect 329868 300804 329924 300814
rect 329868 298872 329924 300748
rect 330316 298872 330372 301868
rect 330764 299908 330820 299918
rect 330764 298872 330820 299852
rect 331212 298872 331268 306908
rect 331324 305172 331380 308056
rect 331324 305106 331380 305116
rect 331660 306852 331716 306862
rect 331660 298872 331716 306796
rect 331772 305620 331828 308056
rect 332248 308028 332388 308084
rect 331772 305554 331828 305564
rect 332108 303828 332164 303838
rect 332108 298872 332164 303772
rect 319116 298340 319172 298350
rect 319116 290668 319172 298284
rect 322028 298340 322084 298350
rect 332332 298340 332388 308028
rect 332668 306852 332724 308056
rect 332668 306786 332724 306796
rect 333004 303940 333060 303950
rect 332556 303604 332612 303614
rect 332556 298872 332612 303548
rect 333004 298872 333060 303884
rect 333116 299908 333172 308056
rect 333564 303604 333620 308056
rect 334012 303940 334068 308056
rect 334012 303874 334068 303884
rect 333564 303538 333620 303548
rect 334460 303044 334516 308056
rect 334908 306964 334964 308056
rect 334908 306898 334964 306908
rect 335356 305732 335412 308056
rect 335356 305666 335412 305676
rect 334460 302978 334516 302988
rect 334796 305060 334852 305070
rect 333116 299842 333172 299852
rect 333452 301812 333508 301822
rect 333452 298872 333508 301756
rect 334348 300804 334404 300814
rect 333900 300468 333956 300478
rect 333900 298872 333956 300412
rect 334348 298872 334404 300748
rect 334796 298872 334852 305004
rect 335020 305060 335076 305070
rect 335020 304276 335076 305004
rect 335020 304210 335076 304220
rect 335692 303716 335748 303726
rect 335244 302260 335300 302270
rect 335244 298872 335300 302204
rect 335692 298872 335748 303660
rect 335804 301588 335860 308056
rect 336252 305396 336308 308056
rect 336252 305330 336308 305340
rect 336588 307412 336644 307422
rect 335804 301522 335860 301532
rect 336140 300916 336196 300926
rect 336140 298872 336196 300860
rect 336588 298872 336644 307356
rect 336700 304836 336756 308056
rect 336700 304770 336756 304780
rect 337036 306516 337092 306526
rect 337036 298872 337092 306460
rect 337148 301924 337204 308056
rect 337148 301858 337204 301868
rect 337596 301812 337652 308056
rect 338044 307412 338100 308056
rect 338044 307346 338100 307356
rect 337596 301746 337652 301756
rect 338380 307188 338436 307198
rect 337484 300132 337540 300142
rect 337484 298872 337540 300076
rect 338380 298872 338436 307132
rect 338492 303716 338548 308056
rect 338492 303650 338548 303660
rect 338828 304052 338884 304062
rect 338828 298872 338884 303996
rect 338940 303828 338996 308056
rect 339388 307188 339444 308056
rect 339388 307122 339444 307132
rect 338940 303762 338996 303772
rect 339724 305284 339780 305294
rect 339276 300020 339332 300030
rect 339276 298872 339332 299964
rect 339724 298872 339780 305228
rect 339836 303940 339892 308056
rect 339836 303874 339892 303884
rect 340172 303380 340228 303390
rect 340172 298872 340228 303324
rect 340284 300020 340340 308056
rect 340760 308028 340900 308084
rect 340284 299954 340340 299964
rect 340620 301476 340676 301486
rect 340620 298872 340676 301420
rect 322084 298284 322728 298340
rect 322028 298274 322084 298284
rect 332332 298274 332388 298284
rect 337932 298340 337988 298350
rect 337932 298274 337988 298284
rect 340844 298340 340900 308028
rect 341180 305172 341236 308056
rect 341180 305106 341236 305116
rect 341628 304500 341684 308056
rect 342076 305172 342132 308056
rect 342076 305106 342132 305116
rect 342412 307076 342468 307086
rect 341628 304434 341684 304444
rect 341516 302372 341572 302382
rect 341068 302036 341124 302046
rect 341068 298872 341124 301980
rect 341516 298872 341572 302316
rect 341964 302148 342020 302158
rect 341964 298872 342020 302092
rect 342412 298872 342468 307020
rect 342524 305732 342580 308056
rect 342524 305666 342580 305676
rect 342860 307300 342916 307310
rect 342524 304724 342580 304734
rect 342524 300916 342580 304668
rect 342524 300850 342580 300860
rect 342860 298872 342916 307244
rect 342972 305732 343028 308056
rect 343420 307076 343476 308056
rect 343868 307300 343924 308056
rect 343868 307234 343924 307244
rect 343420 307010 343476 307020
rect 342972 305666 343028 305676
rect 343756 303156 343812 303166
rect 343308 300356 343364 300366
rect 343308 298872 343364 300300
rect 343756 298872 343812 303100
rect 344204 302932 344260 302942
rect 344204 298872 344260 302876
rect 344316 302036 344372 308056
rect 344316 301970 344372 301980
rect 344652 304164 344708 304174
rect 344652 298872 344708 304108
rect 344764 304052 344820 308056
rect 344764 303986 344820 303996
rect 345212 303380 345268 308056
rect 345660 306404 345716 308056
rect 345660 306338 345716 306348
rect 345212 303314 345268 303324
rect 345996 304948 346052 304958
rect 345548 300916 345604 300926
rect 345100 300804 345156 300814
rect 345100 298872 345156 300748
rect 345548 298872 345604 300860
rect 345996 298872 346052 304892
rect 346108 300132 346164 308056
rect 346108 300066 346164 300076
rect 346444 305284 346500 305294
rect 346444 298872 346500 305228
rect 346556 304948 346612 308056
rect 347004 305620 347060 308056
rect 347004 305554 347060 305564
rect 346556 304882 346612 304892
rect 347340 301700 347396 301710
rect 346892 301140 346948 301150
rect 346892 298872 346948 301084
rect 347340 298872 347396 301644
rect 347452 301476 347508 308056
rect 347900 305284 347956 308056
rect 347900 305218 347956 305228
rect 348236 306628 348292 306638
rect 347452 301410 347508 301420
rect 347788 305172 347844 305182
rect 347788 301252 347844 305116
rect 347788 301186 347844 301196
rect 347788 301028 347844 301038
rect 347788 298872 347844 300972
rect 348236 298872 348292 306572
rect 348348 301140 348404 308056
rect 348796 306628 348852 308056
rect 348796 306562 348852 306572
rect 348348 301074 348404 301084
rect 348684 303492 348740 303502
rect 348684 298872 348740 303436
rect 349132 303268 349188 303278
rect 349132 298872 349188 303212
rect 349244 300356 349300 308056
rect 349356 304388 349412 304398
rect 349356 301028 349412 304332
rect 349692 303268 349748 308056
rect 350140 306516 350196 308056
rect 350140 306450 350196 306460
rect 350476 306740 350532 306750
rect 349692 303202 349748 303212
rect 349356 300962 349412 300972
rect 349580 302596 349636 302606
rect 349244 300290 349300 300300
rect 349580 298872 349636 302540
rect 350028 300244 350084 300254
rect 350028 298872 350084 300188
rect 350476 298872 350532 306684
rect 350588 300244 350644 308056
rect 351036 308018 351092 308028
rect 351148 304612 351204 304622
rect 350588 300178 350644 300188
rect 350924 301028 350980 301038
rect 350924 298872 350980 300972
rect 351148 301028 351204 304556
rect 351484 304612 351540 308056
rect 351484 304546 351540 304556
rect 351932 304276 351988 308056
rect 352380 305732 352436 308056
rect 352380 305666 352436 305676
rect 351932 304210 351988 304220
rect 352828 301700 352884 308056
rect 352828 301634 352884 301644
rect 353164 306852 353220 306862
rect 351148 300962 351204 300972
rect 351820 301364 351876 301374
rect 351372 300804 351428 300814
rect 351372 298872 351428 300748
rect 351820 298872 351876 301308
rect 352268 300916 352324 300926
rect 352268 298872 352324 300860
rect 353164 298872 353220 306796
rect 353276 302036 353332 308056
rect 353724 305508 353780 308056
rect 354172 306852 354228 308056
rect 354172 306786 354228 306796
rect 354620 306740 354676 308056
rect 354620 306674 354676 306684
rect 353724 305442 353780 305452
rect 353276 301970 353332 301980
rect 354060 303604 354116 303614
rect 353612 299908 353668 299918
rect 353612 298872 353668 299852
rect 354060 298872 354116 303548
rect 355068 303492 355124 308056
rect 355068 303426 355124 303436
rect 355404 306964 355460 306974
rect 354956 303044 355012 303054
rect 354508 302932 354564 302942
rect 354508 298872 354564 302876
rect 354956 298872 355012 302988
rect 355404 298872 355460 306908
rect 355516 303268 355572 308056
rect 355964 305732 356020 308056
rect 355964 305666 356020 305676
rect 356188 304948 356244 304958
rect 355516 303202 355572 303212
rect 355852 304164 355908 304174
rect 355852 298872 355908 304108
rect 356188 304164 356244 304892
rect 356412 304948 356468 308056
rect 356412 304882 356468 304892
rect 356188 304098 356244 304108
rect 356300 304836 356356 304846
rect 356300 298872 356356 304780
rect 356860 304724 356916 308056
rect 356860 304658 356916 304668
rect 357308 302148 357364 308056
rect 357756 302260 357812 308056
rect 357756 302194 357812 302204
rect 357308 302082 357364 302092
rect 357644 301924 357700 301934
rect 356748 301588 356804 301598
rect 356748 298872 356804 301532
rect 357196 301028 357252 301038
rect 357196 298872 357252 300972
rect 357644 298872 357700 301868
rect 358092 301812 358148 301822
rect 358092 298872 358148 301756
rect 358204 301588 358260 308056
rect 358204 301522 358260 301532
rect 358540 307412 358596 307422
rect 358540 298872 358596 307356
rect 358652 306964 358708 308056
rect 358652 306898 358708 306908
rect 358988 303716 359044 303726
rect 358988 298872 359044 303660
rect 359100 303604 359156 308056
rect 359100 303538 359156 303548
rect 359436 303828 359492 303838
rect 359436 298872 359492 303772
rect 359548 303716 359604 308056
rect 359996 307412 360052 308056
rect 359996 307346 360052 307356
rect 359548 303650 359604 303660
rect 359884 307188 359940 307198
rect 359884 298872 359940 307132
rect 360332 303940 360388 303950
rect 360332 298872 360388 303884
rect 360444 300580 360500 308056
rect 360892 305732 360948 308056
rect 360892 305666 360948 305676
rect 361340 302932 361396 308056
rect 361340 302866 361396 302876
rect 361676 305060 361732 305070
rect 361676 302820 361732 305004
rect 361788 304500 361844 308056
rect 361788 304434 361844 304444
rect 361676 302764 361956 302820
rect 360444 300514 360500 300524
rect 361676 302596 361732 302606
rect 360780 300020 360836 300030
rect 360780 298872 360836 299964
rect 361676 298872 361732 302540
rect 361900 298900 361956 302764
rect 362236 301812 362292 308056
rect 362684 305620 362740 308056
rect 363132 307188 363188 308056
rect 363132 307122 363188 307132
rect 363580 306292 363636 308056
rect 363580 306226 363636 306236
rect 363916 307076 363972 307086
rect 362684 305554 362740 305564
rect 362236 301746 362292 301756
rect 363468 302484 363524 302494
rect 363020 301364 363076 301374
rect 362572 301252 362628 301262
rect 361900 298844 362152 298900
rect 362572 298872 362628 301196
rect 363020 298872 363076 301308
rect 363468 298872 363524 302428
rect 363916 298872 363972 307020
rect 364028 303828 364084 308056
rect 364028 303762 364084 303772
rect 364140 308028 364504 308084
rect 340844 298274 340900 298284
rect 352716 298340 352772 298350
rect 352716 298274 352772 298284
rect 361228 298340 361284 298350
rect 361228 298274 361284 298284
rect 364140 298340 364196 308028
rect 364364 307300 364420 307310
rect 364364 298872 364420 307244
rect 364924 302820 364980 308056
rect 364924 302754 364980 302764
rect 365260 304052 365316 304062
rect 364812 300804 364868 300814
rect 364812 298872 364868 300748
rect 365260 298872 365316 303996
rect 365372 300468 365428 308056
rect 365820 305284 365876 308056
rect 365820 305218 365876 305228
rect 366156 306404 366212 306414
rect 365372 300402 365428 300412
rect 365708 303380 365764 303390
rect 365708 298872 365764 303324
rect 366156 298872 366212 306348
rect 366268 305396 366324 308056
rect 366268 305330 366324 305340
rect 366716 305060 366772 308056
rect 366716 304994 366772 305004
rect 366828 305508 366884 305518
rect 366604 300132 366660 300142
rect 366604 298872 366660 300076
rect 366828 298900 366884 305452
rect 367164 305508 367220 308056
rect 367164 305442 367220 305452
rect 367500 304164 367556 304174
rect 366828 298844 367080 298900
rect 367500 298872 367556 304108
rect 367612 302372 367668 308056
rect 367612 302306 367668 302316
rect 367948 301476 368004 301486
rect 367948 298872 368004 301420
rect 368060 300132 368116 308056
rect 368060 300066 368116 300076
rect 368396 304388 368452 304398
rect 368396 298872 368452 304332
rect 368508 304164 368564 308056
rect 368508 304098 368564 304108
rect 368956 303940 369012 308056
rect 368956 303874 369012 303884
rect 369292 306628 369348 306638
rect 368844 301140 368900 301150
rect 368844 298872 368900 301084
rect 369292 298872 369348 306572
rect 369404 305732 369460 308056
rect 369404 305666 369460 305676
rect 369740 300356 369796 300366
rect 369740 298872 369796 300300
rect 369852 300020 369908 308056
rect 370300 305620 370356 308056
rect 370300 305554 370356 305564
rect 370636 306516 370692 306526
rect 369852 299954 369908 299964
rect 370188 302932 370244 302942
rect 370188 298872 370244 302876
rect 370636 298872 370692 306460
rect 370748 305060 370804 308056
rect 370748 304994 370804 305004
rect 370860 308028 371224 308084
rect 364140 298274 364196 298284
rect 370860 298340 370916 308028
rect 371420 307972 371476 307982
rect 371196 304276 371252 304286
rect 371196 300916 371252 304220
rect 371308 304164 371364 304174
rect 371308 302932 371364 304108
rect 371308 302866 371364 302876
rect 371420 302428 371476 307916
rect 371644 305284 371700 308056
rect 372092 306516 372148 308056
rect 372540 306628 372596 308056
rect 372540 306562 372596 306572
rect 372092 306450 372148 306460
rect 371644 305218 371700 305228
rect 372988 304948 373044 308056
rect 372988 304882 373044 304892
rect 371980 304052 372036 304062
rect 371420 302372 371588 302428
rect 371196 300850 371252 300860
rect 371084 300244 371140 300254
rect 371084 298872 371140 300188
rect 371532 298872 371588 302372
rect 371980 298872 372036 303996
rect 373436 303380 373492 308056
rect 373884 304612 373940 308056
rect 373884 304546 373940 304556
rect 374220 305172 374276 305182
rect 373436 303314 373492 303324
rect 373772 302036 373828 302046
rect 373324 301700 373380 301710
rect 372876 300916 372932 300926
rect 372428 300804 372484 300814
rect 372428 298872 372484 300748
rect 372876 298872 372932 300860
rect 373324 298872 373380 301644
rect 373772 298872 373828 301980
rect 374220 298872 374276 305116
rect 374332 302148 374388 308056
rect 374332 302082 374388 302092
rect 374668 306852 374724 306862
rect 374668 298872 374724 306796
rect 374780 306404 374836 308056
rect 374780 306338 374836 306348
rect 375116 306740 375172 306750
rect 375116 298872 375172 306684
rect 375228 304836 375284 308056
rect 375228 304770 375284 304780
rect 375676 304052 375732 308056
rect 375676 303986 375732 303996
rect 375340 303268 375396 303278
rect 375340 298900 375396 303212
rect 376012 303156 376068 303166
rect 375340 298844 375592 298900
rect 376012 298872 376068 303100
rect 376124 301700 376180 308056
rect 376572 307076 376628 308056
rect 376572 307010 376628 307020
rect 376236 304612 376292 304622
rect 376236 303492 376292 304556
rect 376236 303426 376292 303436
rect 376460 304164 376516 304174
rect 376124 301634 376180 301644
rect 376460 298872 376516 304108
rect 376908 300916 376964 300926
rect 376908 298872 376964 300860
rect 377020 299908 377076 308056
rect 377244 304500 377300 304510
rect 377244 300916 377300 304444
rect 377468 303268 377524 308056
rect 377916 305732 377972 308056
rect 378812 307300 378868 308056
rect 378812 307234 378868 307244
rect 377916 305666 377972 305676
rect 379148 306964 379204 306974
rect 377468 303202 377524 303212
rect 378252 302260 378308 302270
rect 377244 300850 377300 300860
rect 377804 302036 377860 302046
rect 377020 299842 377076 299852
rect 377356 300804 377412 300814
rect 377356 298872 377412 300748
rect 377804 298872 377860 301980
rect 378252 298872 378308 302204
rect 378700 301588 378756 301598
rect 378700 298872 378756 301532
rect 379148 298872 379204 306908
rect 379260 301588 379316 308056
rect 379260 301522 379316 301532
rect 379596 303604 379652 303614
rect 379596 298872 379652 303548
rect 379708 301924 379764 308056
rect 380156 304612 380212 308056
rect 380156 304546 380212 304556
rect 380492 307412 380548 307422
rect 379708 301858 379764 301868
rect 380044 303716 380100 303726
rect 380044 298872 380100 303660
rect 380492 298872 380548 307356
rect 380604 304052 380660 308056
rect 381052 305732 381108 308056
rect 381500 306740 381556 308056
rect 381500 306674 381556 306684
rect 381052 305666 381108 305676
rect 380604 303986 380660 303996
rect 381948 303604 382004 308056
rect 382396 306852 382452 308056
rect 382396 306786 382452 306796
rect 381948 303538 382004 303548
rect 381388 303156 381444 303166
rect 380940 300580 380996 300590
rect 380940 298872 380996 300524
rect 381388 298872 381444 303100
rect 382732 301812 382788 301822
rect 381836 301364 381892 301374
rect 381836 298872 381892 301308
rect 382284 300916 382340 300926
rect 382284 298872 382340 300860
rect 382732 298872 382788 301756
rect 382844 300244 382900 308056
rect 383292 307412 383348 308056
rect 383292 307346 383348 307356
rect 383628 307188 383684 307198
rect 382844 300178 382900 300188
rect 383180 300804 383236 300814
rect 383180 298872 383236 300748
rect 383628 298872 383684 307132
rect 383740 301812 383796 308056
rect 384076 306292 384132 306302
rect 383964 304052 384020 304062
rect 383964 302148 384020 303996
rect 383964 302082 384020 302092
rect 383740 301746 383796 301756
rect 384076 298872 384132 306236
rect 384188 304500 384244 308056
rect 384188 304434 384244 304444
rect 384524 303828 384580 303838
rect 384524 298872 384580 303772
rect 384636 302036 384692 308056
rect 398860 308084 398916 308094
rect 385084 308018 385140 308028
rect 385532 306964 385588 308056
rect 385532 306898 385588 306908
rect 384636 301970 384692 301980
rect 385420 303044 385476 303054
rect 385420 298872 385476 302988
rect 385980 300580 386036 308056
rect 386428 303156 386484 308056
rect 386428 303090 386484 303100
rect 386764 305396 386820 305406
rect 385980 300514 386036 300524
rect 386316 301476 386372 301486
rect 385868 300468 385924 300478
rect 385868 298872 385924 300412
rect 386316 298872 386372 301420
rect 386764 298872 386820 305340
rect 386876 303828 386932 308056
rect 386876 303762 386932 303772
rect 387324 302820 387380 308056
rect 387324 302754 387380 302764
rect 387660 305172 387716 305182
rect 387212 302484 387268 302494
rect 387212 298872 387268 302428
rect 387660 298872 387716 305116
rect 387772 304836 387828 308056
rect 387772 304770 387828 304780
rect 388108 305620 388164 305630
rect 388108 304052 388164 305564
rect 388108 303986 388164 303996
rect 388108 300804 388164 300814
rect 388108 298872 388164 300748
rect 388220 300356 388276 308056
rect 388668 304724 388724 308056
rect 389116 305172 389172 308056
rect 389116 305106 389172 305116
rect 388668 304658 388724 304668
rect 389452 303940 389508 303950
rect 388220 300290 388276 300300
rect 389004 302932 389060 302942
rect 388556 300132 388612 300142
rect 388556 298872 388612 300076
rect 389004 298872 389060 302876
rect 389452 298872 389508 303884
rect 389564 302260 389620 308056
rect 390012 303828 390068 308056
rect 390012 303762 390068 303772
rect 389564 302194 389620 302204
rect 389900 303156 389956 303166
rect 389900 298872 389956 303100
rect 390460 300132 390516 308056
rect 390460 300066 390516 300076
rect 390796 304052 390852 304062
rect 390348 300020 390404 300030
rect 390348 298872 390404 299964
rect 390796 298872 390852 303996
rect 390908 303940 390964 308056
rect 390908 303874 390964 303884
rect 391244 305060 391300 305070
rect 391244 298872 391300 305004
rect 391356 304276 391412 308056
rect 391804 306292 391860 308056
rect 392252 307188 392308 308056
rect 392252 307122 392308 307132
rect 391804 306226 391860 306236
rect 392588 306516 392644 306526
rect 391356 304210 391412 304220
rect 392140 305284 392196 305294
rect 392140 298872 392196 305228
rect 392588 298872 392644 306460
rect 392700 305732 392756 308056
rect 392700 305666 392756 305676
rect 393036 306628 393092 306638
rect 393036 298872 393092 306572
rect 393148 305396 393204 308056
rect 393596 305508 393652 308056
rect 394044 305620 394100 308056
rect 394044 305554 394100 305564
rect 393596 305442 393652 305452
rect 393148 305330 393204 305340
rect 394492 305284 394548 308056
rect 394492 305218 394548 305228
rect 393484 304948 393540 304958
rect 393484 298872 393540 304892
rect 394828 304836 394884 304846
rect 393820 304612 393876 304622
rect 393708 303380 393764 303390
rect 393708 298900 393764 303324
rect 393820 301364 393876 304556
rect 393932 304500 393988 304510
rect 393932 301476 393988 304444
rect 393932 301410 393988 301420
rect 394380 303492 394436 303502
rect 393820 301298 393876 301308
rect 393708 298844 393960 298900
rect 394380 298872 394436 303436
rect 394828 302260 394884 304780
rect 394940 303492 394996 308056
rect 394940 303426 394996 303436
rect 395276 306404 395332 306414
rect 394828 302194 394884 302204
rect 394828 300804 394884 300814
rect 394828 298872 394884 300748
rect 395276 298872 395332 306348
rect 395388 305060 395444 308056
rect 395836 305284 395892 308056
rect 395836 305218 395892 305228
rect 395388 304994 395444 305004
rect 395724 304052 395780 304062
rect 395724 298872 395780 303996
rect 395948 304052 396004 304062
rect 395948 303716 396004 303996
rect 395948 303650 396004 303660
rect 396172 303716 396228 303726
rect 396172 303044 396228 303660
rect 396284 303380 396340 308056
rect 396732 304948 396788 308056
rect 396732 304882 396788 304892
rect 397068 307076 397124 307086
rect 396284 303314 396340 303324
rect 396172 302978 396228 302988
rect 396172 302372 396228 302382
rect 396172 298872 396228 302316
rect 396620 301700 396676 301710
rect 396620 298872 396676 301644
rect 397068 298872 397124 307020
rect 397964 303268 398020 303278
rect 397516 299908 397572 299918
rect 397516 298872 397572 299852
rect 397964 298872 398020 303212
rect 398412 303156 398468 303166
rect 398412 298872 398468 303100
rect 398860 298872 398916 308028
rect 405580 307972 405636 307982
rect 403788 307412 403844 307422
rect 399308 307300 399364 307310
rect 399308 298872 399364 307244
rect 402892 306852 402948 306862
rect 401996 306740 402052 306750
rect 401548 304164 401604 304174
rect 401100 302148 401156 302158
rect 400204 301924 400260 301934
rect 399756 301588 399812 301598
rect 399756 298872 399812 301532
rect 400204 298872 400260 301868
rect 400652 301364 400708 301374
rect 400652 298872 400708 301308
rect 401100 298872 401156 302092
rect 401548 298872 401604 304108
rect 401996 298872 402052 306684
rect 402332 304724 402388 304734
rect 402332 302484 402388 304668
rect 402332 302418 402388 302428
rect 402444 303604 402500 303614
rect 402444 298872 402500 303548
rect 402892 298872 402948 306796
rect 403340 300244 403396 300254
rect 403340 298872 403396 300188
rect 403788 298872 403844 307356
rect 405132 302036 405188 302046
rect 404236 301812 404292 301822
rect 404236 298872 404292 301756
rect 404684 301476 404740 301486
rect 404684 298872 404740 301420
rect 405132 298872 405188 301980
rect 405580 298872 405636 307916
rect 411516 307524 411572 307534
rect 406028 306964 406084 306974
rect 406028 298872 406084 306908
rect 409612 305172 409668 305182
rect 407372 304052 407428 304062
rect 406924 303716 406980 303726
rect 406476 300580 406532 300590
rect 406476 298872 406532 300524
rect 406924 298872 406980 303660
rect 407372 298872 407428 303996
rect 407820 303044 407876 303054
rect 407820 298872 407876 302988
rect 409164 302484 409220 302494
rect 408268 302260 408324 302270
rect 408268 298872 408324 302204
rect 408716 300356 408772 300366
rect 408716 298872 408772 300300
rect 409164 298872 409220 302428
rect 409612 298872 409668 305116
rect 411516 304164 411572 307468
rect 418348 307524 418404 314188
rect 418348 307458 418404 307468
rect 412748 307188 412804 307198
rect 411516 304098 411572 304108
rect 412300 306292 412356 306302
rect 411404 303940 411460 303950
rect 410508 303828 410564 303838
rect 410060 300804 410116 300814
rect 410060 298872 410116 300748
rect 410508 298872 410564 303772
rect 410956 300132 411012 300142
rect 410956 298872 411012 300076
rect 411404 298872 411460 303884
rect 411852 302932 411908 302942
rect 411852 298872 411908 302876
rect 412300 298872 412356 306236
rect 412748 298872 412804 307132
rect 413196 305732 413252 305742
rect 413196 298872 413252 305676
rect 414540 305620 414596 305630
rect 414092 305508 414148 305518
rect 413644 305396 413700 305406
rect 413644 298872 413700 305340
rect 414092 298872 414148 305452
rect 414540 298872 414596 305564
rect 416332 305284 416388 305294
rect 415884 305060 415940 305070
rect 415436 303492 415492 303502
rect 414988 300804 415044 300814
rect 414988 298872 415044 300748
rect 415436 298872 415492 303436
rect 415884 298872 415940 305004
rect 416332 298872 416388 305228
rect 417228 304948 417284 304958
rect 416780 303380 416836 303390
rect 416780 298872 416836 303324
rect 417228 298872 417284 304892
rect 370860 298274 370916 298284
rect 384972 298340 385028 298350
rect 384972 298274 385028 298284
rect 391692 298340 391748 298350
rect 391692 298274 391748 298284
rect 319004 290612 319172 290668
rect 319004 95060 319060 290612
rect 319004 94994 319060 95004
rect 419132 94948 419188 333452
rect 423276 320964 423332 320974
rect 423276 314244 423332 320908
rect 423276 314178 423332 314188
rect 420140 299124 420196 299134
rect 420028 298116 420084 298126
rect 420028 258692 420084 298060
rect 420140 285684 420196 299068
rect 420140 285618 420196 285628
rect 420028 258626 420084 258636
rect 419132 94882 419188 94892
rect 421596 89908 421652 89918
rect 318892 86818 318948 86828
rect 351036 88116 351092 88126
rect 318332 86706 318388 86716
rect 319116 86212 319172 86222
rect 315644 84914 315700 84924
rect 315756 85316 315812 85326
rect 301756 83458 301812 83468
rect 314972 84532 315028 84542
rect 299180 83122 299236 83132
rect 298620 81666 298676 81676
rect 292236 80434 292292 80444
rect 295596 81284 295652 81294
rect 287196 78306 287252 78316
rect 295596 78260 295652 81228
rect 295596 78194 295652 78204
rect 314972 78260 315028 84476
rect 315756 83300 315812 85260
rect 317324 84644 317380 84654
rect 317324 83860 317380 84588
rect 317324 83794 317380 83804
rect 317436 84532 317492 84542
rect 317436 83748 317492 84476
rect 319116 83972 319172 86156
rect 319116 83906 319172 83916
rect 340956 86100 341012 86110
rect 317436 83682 317492 83692
rect 340956 83524 341012 86044
rect 351036 83636 351092 88060
rect 421596 87332 421652 89852
rect 421596 87266 421652 87276
rect 414988 86100 415044 86110
rect 414988 83972 415044 86044
rect 414988 83906 415044 83916
rect 422828 84308 422884 84318
rect 351036 83570 351092 83580
rect 340956 83458 341012 83468
rect 315756 83234 315812 83244
rect 419132 83300 419188 83310
rect 416668 82628 416724 82638
rect 416668 81508 416724 82572
rect 416668 81442 416724 81452
rect 419132 78484 419188 83244
rect 422828 82292 422884 84252
rect 422828 82226 422884 82236
rect 424172 80164 424228 393932
rect 427084 392644 427140 395080
rect 427084 392578 427140 392588
rect 428428 392644 428484 392654
rect 428428 391412 428484 392588
rect 428428 391346 428484 391356
rect 431116 387828 431172 395080
rect 435148 390740 435204 395080
rect 439180 391076 439236 395080
rect 443212 391188 443268 395080
rect 443212 391122 443268 391132
rect 439180 391010 439236 391020
rect 435148 390674 435204 390684
rect 446796 390516 446852 390526
rect 431116 387762 431172 387772
rect 442652 389396 442708 389406
rect 430892 383908 430948 383918
rect 429212 380548 429268 380558
rect 425852 373828 425908 373838
rect 424396 372148 424452 372158
rect 424396 80276 424452 372092
rect 424956 341012 425012 341022
rect 424956 333508 425012 340956
rect 424956 333442 425012 333452
rect 425068 324324 425124 324334
rect 425068 320964 425124 324268
rect 425068 320898 425124 320908
rect 425180 84868 425236 84878
rect 425068 83188 425124 83198
rect 425068 80612 425124 83132
rect 425068 80546 425124 80556
rect 425180 80500 425236 84812
rect 425180 80434 425236 80444
rect 425852 80388 425908 373772
rect 426748 368900 426804 368910
rect 426748 362852 426804 368844
rect 426748 362786 426804 362796
rect 427532 368788 427588 368798
rect 427532 341012 427588 368732
rect 427532 340946 427588 340956
rect 428764 92820 428820 92830
rect 425852 80322 425908 80332
rect 428204 82740 428260 82750
rect 424396 80210 424452 80220
rect 424172 80098 424228 80108
rect 419132 78418 419188 78428
rect 314972 78194 315028 78204
rect 270620 77074 270676 77084
rect 270284 23090 270340 23100
rect 269836 18498 269892 18508
rect 269724 16146 269780 16156
rect 270396 16772 270452 16782
rect 269948 15764 270004 15774
rect 269612 13346 269668 13356
rect 269724 13748 269780 13758
rect 269500 7970 269556 7980
rect 268940 6514 268996 6524
rect 269724 6468 269780 13692
rect 269836 12628 269892 12638
rect 269836 10164 269892 12572
rect 269948 10388 270004 15708
rect 269948 10322 270004 10332
rect 270284 13636 270340 13646
rect 269836 10108 270004 10164
rect 269724 6402 269780 6412
rect 269836 9940 269892 9950
rect 269836 1652 269892 9884
rect 269948 5796 270004 10108
rect 269948 5730 270004 5740
rect 270172 8260 270228 8270
rect 270172 4452 270228 8204
rect 270172 4386 270228 4396
rect 269836 1586 269892 1596
rect 268492 1362 268548 1372
rect 270284 480 270340 13580
rect 270396 4340 270452 16716
rect 270620 14532 270676 14542
rect 270396 4274 270452 4284
rect 270508 11172 270564 11182
rect 270508 3220 270564 11116
rect 270508 3154 270564 3164
rect 270620 532 270676 14476
rect 275324 10500 275380 10510
rect 275212 10052 275268 10062
rect 275212 5348 275268 9996
rect 275212 5282 275268 5292
rect 275324 4452 275380 10444
rect 312396 10500 312452 10510
rect 287084 10388 287140 10398
rect 277228 9828 277284 9838
rect 275436 7028 275492 7038
rect 275436 5236 275492 6972
rect 275436 5170 275492 5180
rect 275660 5348 275716 5358
rect 275324 4386 275380 4396
rect 275548 5124 275604 5134
rect 274092 4340 274148 4350
rect 249340 392 249592 480
rect 251244 392 251496 480
rect 253148 392 253400 480
rect 255052 392 255304 480
rect 248668 354 248724 364
rect 249368 -960 249592 392
rect 251272 -960 251496 392
rect 253176 -960 253400 392
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 260764 392 261016 480
rect 262668 392 262920 480
rect 264572 392 264824 480
rect 266476 392 266728 480
rect 268380 392 268632 480
rect 270284 392 270536 480
rect 270620 466 270676 476
rect 272188 4228 272244 4238
rect 272188 480 272244 4172
rect 274092 480 274148 4284
rect 275548 2548 275604 5068
rect 275548 2482 275604 2492
rect 275660 2100 275716 5292
rect 277228 4900 277284 9772
rect 277564 9156 277620 9166
rect 277452 8820 277508 8830
rect 277340 8708 277396 8718
rect 277340 8372 277396 8652
rect 277340 8306 277396 8316
rect 277228 4834 277284 4844
rect 275996 4004 276052 4014
rect 275772 3556 275828 3566
rect 275772 3220 275828 3500
rect 275772 3154 275828 3164
rect 275660 2034 275716 2044
rect 275996 480 276052 3948
rect 277452 3108 277508 8764
rect 277452 3042 277508 3052
rect 277564 2436 277620 9100
rect 279132 8596 279188 8606
rect 278908 8484 278964 8494
rect 277564 2370 277620 2380
rect 277900 6244 277956 6254
rect 277900 480 277956 6188
rect 278908 3332 278964 8428
rect 278908 3266 278964 3276
rect 279132 1428 279188 8540
rect 283612 8260 283668 8270
rect 280812 7028 280868 7038
rect 280812 6356 280868 6972
rect 280812 6290 280868 6300
rect 281708 6916 281764 6926
rect 279132 1362 279188 1372
rect 279804 4900 279860 4910
rect 279804 480 279860 4844
rect 280476 3668 280532 3678
rect 280364 2772 280420 2782
rect 280364 1092 280420 2716
rect 280476 1652 280532 3612
rect 280476 1586 280532 1596
rect 280364 1026 280420 1036
rect 281708 480 281764 6860
rect 282156 3780 282212 3790
rect 282156 1652 282212 3724
rect 282156 1586 282212 1596
rect 283612 480 283668 8204
rect 285852 7028 285908 7038
rect 285628 6916 285684 6926
rect 285628 6468 285684 6860
rect 285628 6402 285684 6412
rect 285740 5236 285796 5246
rect 285628 3780 285684 3790
rect 285628 2324 285684 3724
rect 285740 3108 285796 5180
rect 285852 3388 285908 6972
rect 287084 6356 287140 10332
rect 310716 10164 310772 10174
rect 290668 8820 290724 8830
rect 288988 8708 289044 8718
rect 288988 8372 289044 8652
rect 288988 8306 289044 8316
rect 289100 8596 289156 8606
rect 289100 6692 289156 8540
rect 289100 6626 289156 6636
rect 290668 6692 290724 8764
rect 297164 8820 297220 8830
rect 290668 6626 290724 6636
rect 293132 8148 293188 8158
rect 287084 6290 287140 6300
rect 291228 6020 291284 6030
rect 287308 4900 287364 4910
rect 285852 3332 286132 3388
rect 285740 3042 285796 3052
rect 286076 2660 286132 3332
rect 286076 2594 286132 2604
rect 285628 2258 285684 2268
rect 287308 2212 287364 4844
rect 287308 2146 287364 2156
rect 287420 3668 287476 3678
rect 285404 532 285460 542
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 275996 392 276248 480
rect 277900 392 278152 480
rect 279804 392 280056 480
rect 281708 392 281960 480
rect 283612 392 283864 480
rect 285460 480 285572 532
rect 287420 480 287476 3612
rect 289324 2772 289380 2782
rect 289324 480 289380 2716
rect 291228 480 291284 5964
rect 293132 480 293188 8092
rect 295820 7028 295876 7038
rect 295820 6692 295876 6972
rect 295820 6626 295876 6636
rect 297164 6468 297220 8764
rect 304108 8708 304164 8718
rect 297164 6402 297220 6412
rect 302652 7140 302708 7150
rect 295372 6244 295428 6254
rect 294028 3220 294084 3230
rect 294028 1428 294084 3164
rect 294028 1362 294084 1372
rect 295036 2436 295092 2446
rect 295036 480 295092 2380
rect 295372 2436 295428 6188
rect 300748 5796 300804 5806
rect 295372 2370 295428 2380
rect 295484 5236 295540 5246
rect 295484 2100 295540 5180
rect 296492 5124 296548 5134
rect 296492 4900 296548 5068
rect 296492 4834 296548 4844
rect 298844 4900 298900 4910
rect 295484 2034 295540 2044
rect 296940 4452 296996 4462
rect 296940 480 296996 4396
rect 297388 3780 297444 3790
rect 297388 2884 297444 3724
rect 297388 2818 297444 2828
rect 297612 3556 297668 3566
rect 297612 2772 297668 3500
rect 297612 2706 297668 2716
rect 298844 480 298900 4844
rect 300748 480 300804 5740
rect 302652 480 302708 7084
rect 303996 6916 304052 6926
rect 303996 5124 304052 6860
rect 303996 5058 304052 5068
rect 304108 3332 304164 8652
rect 308364 6580 308420 6590
rect 304108 3266 304164 3276
rect 307356 5124 307412 5134
rect 307356 3220 307412 5068
rect 307356 3154 307412 3164
rect 304556 2660 304612 2670
rect 304556 480 304612 2604
rect 308252 2660 308308 2670
rect 308252 2436 308308 2604
rect 308252 2370 308308 2380
rect 305676 1988 305732 1998
rect 305676 1540 305732 1932
rect 305676 1474 305732 1484
rect 306796 532 306852 542
rect 306684 480 306796 532
rect 285460 476 285768 480
rect 285404 466 285460 476
rect 285516 392 285768 476
rect 287420 392 287672 480
rect 289324 392 289576 480
rect 291228 392 291480 480
rect 293132 392 293384 480
rect 295036 392 295288 480
rect 296940 392 297192 480
rect 298844 392 299096 480
rect 300748 392 301000 480
rect 302652 392 302904 480
rect 304556 392 304808 480
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262696 -960 262920 392
rect 264600 -960 264824 392
rect 266504 -960 266728 392
rect 268408 -960 268632 392
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277928 -960 278152 392
rect 279832 -960 280056 392
rect 281736 -960 281960 392
rect 283640 -960 283864 392
rect 285544 -960 285768 392
rect 287448 -960 287672 392
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 293160 -960 293384 392
rect 295064 -960 295288 392
rect 296968 -960 297192 392
rect 298872 -960 299096 392
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304584 -960 304808 392
rect 306488 476 306796 480
rect 306488 392 306740 476
rect 306796 466 306852 476
rect 308364 480 308420 6524
rect 310716 6020 310772 10108
rect 310716 5954 310772 5964
rect 310268 3780 310324 3790
rect 309148 3556 309204 3566
rect 309148 1988 309204 3500
rect 309148 1922 309204 1932
rect 310268 480 310324 3724
rect 312396 480 312452 10444
rect 420700 10500 420756 10510
rect 413084 10388 413140 10398
rect 314188 9940 314244 9950
rect 314188 480 314244 9884
rect 365484 9716 365540 9726
rect 331212 9604 331268 9614
rect 319788 8036 319844 8046
rect 318108 4452 318164 4462
rect 315980 3444 316036 3454
rect 315980 480 316036 3388
rect 318108 480 318164 4396
rect 308364 392 308616 480
rect 310268 392 310520 480
rect 306488 -960 306712 392
rect 308392 -960 308616 392
rect 310296 -960 310520 392
rect 312200 392 312452 480
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 316008 -960 316232 392
rect 317912 392 318164 480
rect 319788 480 319844 7980
rect 324268 5236 324324 5246
rect 320908 4788 320964 4798
rect 320908 2884 320964 4732
rect 323820 3780 323876 3790
rect 320908 2818 320964 2828
rect 321692 3556 321748 3566
rect 321692 480 321748 3500
rect 323820 480 323876 3724
rect 324268 3220 324324 5180
rect 324268 3154 324324 3164
rect 327404 4340 327460 4350
rect 319788 392 320040 480
rect 321692 392 321944 480
rect 317912 -960 318136 392
rect 319816 -960 320040 392
rect 321720 -960 321944 392
rect 323624 392 323876 480
rect 325500 2772 325556 2782
rect 325500 480 325556 2716
rect 327404 480 327460 4284
rect 329532 4340 329588 4350
rect 329532 480 329588 4284
rect 325500 392 325752 480
rect 327404 392 327656 480
rect 323624 -960 323848 392
rect 325528 -960 325752 392
rect 327432 -960 327656 392
rect 329336 392 329588 480
rect 331212 480 331268 9548
rect 336924 9492 336980 9502
rect 333116 4564 333172 4574
rect 333116 480 333172 4508
rect 335244 4564 335300 4574
rect 335244 480 335300 4508
rect 331212 392 331464 480
rect 333116 392 333368 480
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 335048 392 335300 480
rect 336924 480 336980 9436
rect 358092 9492 358148 9502
rect 342748 9380 342804 9390
rect 340956 6244 341012 6254
rect 338828 1764 338884 1774
rect 338828 480 338884 1708
rect 340956 480 341012 6188
rect 342748 480 342804 9324
rect 346668 9380 346724 9390
rect 344540 4676 344596 4686
rect 344540 480 344596 4620
rect 346668 480 346724 9324
rect 357196 8596 357252 8606
rect 357196 8260 357252 8540
rect 357196 8194 357252 8204
rect 354060 7028 354116 7038
rect 336924 392 337176 480
rect 338828 392 339080 480
rect 335048 -960 335272 392
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 340760 392 341012 480
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344540 392 344792 480
rect 344568 -960 344792 392
rect 346472 392 346724 480
rect 348348 6468 348404 6478
rect 348348 480 348404 6412
rect 350252 6356 350308 6366
rect 350252 480 350308 6300
rect 352716 4228 352772 4238
rect 352380 4116 352436 4126
rect 352380 480 352436 4060
rect 352716 2772 352772 4172
rect 352716 2706 352772 2716
rect 348348 392 348600 480
rect 350252 392 350504 480
rect 346472 -960 346696 392
rect 348376 -960 348600 392
rect 350280 -960 350504 392
rect 352184 392 352436 480
rect 354060 480 354116 6972
rect 355964 3108 356020 3118
rect 355964 480 356020 3052
rect 358092 480 358148 9436
rect 361676 8260 361732 8270
rect 354060 392 354312 480
rect 355964 392 356216 480
rect 352184 -960 352408 392
rect 354088 -960 354312 392
rect 355992 -960 356216 392
rect 357896 392 358148 480
rect 359772 6132 359828 6142
rect 359772 480 359828 6076
rect 361676 480 361732 8204
rect 363804 7028 363860 7038
rect 362796 6132 362852 6142
rect 362796 4116 362852 6076
rect 362796 4050 362852 4060
rect 363804 480 363860 6972
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 392 363860 480
rect 365484 480 365540 9660
rect 398188 9716 398244 9726
rect 370412 9604 370468 9614
rect 370412 7028 370468 9548
rect 398076 8036 398132 8046
rect 397964 7980 398076 8036
rect 370412 6962 370468 6972
rect 376908 7924 376964 7934
rect 373100 6916 373156 6926
rect 367388 4788 367444 4798
rect 367388 480 367444 4732
rect 369516 3444 369572 3454
rect 369516 480 369572 3388
rect 371308 3220 371364 3230
rect 371308 480 371364 3164
rect 373100 480 373156 6860
rect 375228 3668 375284 3678
rect 375228 480 375284 3612
rect 365484 392 365736 480
rect 367388 392 367640 480
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 369320 392 369572 480
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373100 392 373352 480
rect 373128 -960 373352 392
rect 375032 392 375284 480
rect 376908 480 376964 7868
rect 380940 7924 380996 7934
rect 378812 3556 378868 3566
rect 378812 480 378868 3500
rect 380940 480 380996 7868
rect 376908 392 377160 480
rect 378812 392 379064 480
rect 375032 -960 375256 392
rect 376936 -960 377160 392
rect 378840 -960 379064 392
rect 380744 392 380996 480
rect 382620 7812 382676 7822
rect 382620 480 382676 7756
rect 386652 7812 386708 7822
rect 384412 480 384580 532
rect 386652 480 386708 7756
rect 390460 6916 390516 6926
rect 382620 392 382872 480
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 384412 476 384776 480
rect 384412 420 384468 476
rect 384524 392 384776 476
rect 384412 354 384468 364
rect 384552 -960 384776 392
rect 386456 392 386708 480
rect 388332 5908 388388 5918
rect 388332 480 388388 5852
rect 390460 480 390516 6860
rect 394828 6468 394884 6478
rect 392364 5908 392420 5918
rect 392364 480 392420 5852
rect 394828 4452 394884 6412
rect 394828 4386 394884 4396
rect 388332 392 388584 480
rect 386456 -960 386680 392
rect 388360 -960 388584 392
rect 390264 392 390516 480
rect 392168 392 392420 480
rect 394044 3444 394100 3454
rect 394044 480 394100 3388
rect 397740 3444 397796 3454
rect 397740 532 397796 3388
rect 395836 480 396004 532
rect 394044 392 394296 480
rect 390264 -960 390488 392
rect 392168 -960 392392 392
rect 394072 -960 394296 392
rect 395836 476 396200 480
rect 395836 308 395892 476
rect 395948 392 396200 476
rect 397964 480 398020 7980
rect 398076 7970 398132 7980
rect 398188 6916 398244 9660
rect 398188 6850 398244 6860
rect 399868 9268 399924 9278
rect 398076 3668 398132 3678
rect 398076 1652 398132 3612
rect 398076 1586 398132 1596
rect 399868 480 399924 9212
rect 408268 9268 408324 9278
rect 403788 8148 403844 8158
rect 401884 6356 401940 6366
rect 401884 480 401940 6300
rect 403788 480 403844 8092
rect 408268 6468 408324 9212
rect 408268 6402 408324 6412
rect 411180 6804 411236 6814
rect 407596 4452 407652 4462
rect 406588 3444 406644 3454
rect 397740 466 397796 476
rect 395836 242 395892 252
rect 395976 -960 396200 392
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 392 401940 480
rect 403592 392 403844 480
rect 405468 2996 405524 3006
rect 405468 480 405524 2940
rect 406588 1540 406644 3388
rect 406588 1474 406644 1484
rect 407596 480 407652 4396
rect 409500 4228 409556 4238
rect 409500 480 409556 4172
rect 405468 392 405720 480
rect 401688 -960 401912 392
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 407400 392 407652 480
rect 409304 392 409556 480
rect 411180 480 411236 6748
rect 413084 480 413140 10332
rect 413196 8260 413252 8270
rect 413196 4564 413252 8204
rect 419020 4900 419076 4910
rect 417116 4788 417172 4798
rect 413196 4498 413252 4508
rect 415212 4564 415268 4574
rect 415212 480 415268 4508
rect 416668 3780 416724 3790
rect 416668 3108 416724 3724
rect 416668 3042 416724 3052
rect 417116 480 417172 4732
rect 419020 480 419076 4844
rect 420700 4452 420756 10444
rect 428204 9716 428260 82684
rect 428204 9650 428260 9660
rect 428428 7700 428484 7710
rect 425068 6804 425124 6814
rect 425068 4788 425124 6748
rect 425068 4722 425124 4732
rect 420700 4386 420756 4396
rect 422604 4228 422660 4238
rect 420924 4116 420980 4126
rect 420924 480 420980 4060
rect 411180 392 411432 480
rect 413084 392 413336 480
rect 407400 -960 407624 392
rect 409304 -960 409528 392
rect 411208 -960 411432 392
rect 413112 -960 413336 392
rect 415016 392 415268 480
rect 416920 392 417172 480
rect 418824 392 419076 480
rect 420728 392 420980 480
rect 422604 480 422660 4172
rect 424508 4228 424564 4238
rect 424508 480 424564 4172
rect 426636 4228 426692 4238
rect 426636 480 426692 4172
rect 428428 480 428484 7644
rect 428764 6804 428820 92764
rect 428988 84420 429044 84430
rect 428988 34468 429044 84364
rect 428988 34402 429044 34412
rect 429100 82516 429156 82526
rect 429100 14644 429156 82460
rect 429212 80052 429268 380492
rect 429324 338660 429380 338670
rect 429324 324324 429380 338604
rect 429324 324258 429380 324268
rect 430108 299348 430164 299358
rect 429660 89124 429716 89134
rect 429436 87892 429492 87902
rect 429212 79986 429268 79996
rect 429324 84644 429380 84654
rect 429100 14578 429156 14588
rect 428764 6738 428820 6748
rect 429324 4340 429380 84588
rect 429436 8036 429492 87836
rect 429436 7970 429492 7980
rect 429548 82628 429604 82638
rect 429548 5908 429604 82572
rect 429660 22708 429716 89068
rect 429660 22642 429716 22652
rect 429884 84980 429940 84990
rect 429884 14756 429940 84924
rect 429996 80500 430052 80510
rect 429996 22820 430052 80444
rect 429996 22754 430052 22764
rect 429884 14690 429940 14700
rect 429548 5842 429604 5852
rect 429324 4274 429380 4284
rect 430108 4116 430164 299292
rect 430220 298452 430276 298462
rect 430220 4228 430276 298396
rect 430220 4162 430276 4172
rect 430332 87332 430388 87342
rect 430108 4050 430164 4060
rect 430332 480 430388 87276
rect 430892 79940 430948 383852
rect 434252 375508 434308 375518
rect 430892 79874 430948 79884
rect 431004 95956 431060 95966
rect 430892 78484 430948 78494
rect 430892 11284 430948 78428
rect 431004 20132 431060 95900
rect 432796 94612 432852 94622
rect 432572 94164 432628 94174
rect 431004 20066 431060 20076
rect 431116 92708 431172 92718
rect 431116 18452 431172 92652
rect 431116 18386 431172 18396
rect 431228 86100 431284 86110
rect 430892 11218 430948 11228
rect 431228 10948 431284 86044
rect 431452 83524 431508 83534
rect 431452 11172 431508 83468
rect 432572 18228 432628 94108
rect 432572 18162 432628 18172
rect 432684 87668 432740 87678
rect 432684 14868 432740 87612
rect 432796 19572 432852 94556
rect 432796 19506 432852 19516
rect 432908 92596 432964 92606
rect 432908 18004 432964 92540
rect 434028 83636 434084 83646
rect 433020 80724 433076 80734
rect 433020 32004 433076 80668
rect 433020 31938 433076 31948
rect 432908 17938 432964 17948
rect 432684 14802 432740 14812
rect 431452 11106 431508 11116
rect 431228 10882 431284 10892
rect 432124 4228 432180 4238
rect 432124 480 432180 4172
rect 434028 480 434084 83580
rect 434252 79828 434308 375452
rect 435932 373044 435988 373054
rect 435932 93268 435988 372988
rect 440188 372484 440244 372494
rect 436044 372372 436100 372382
rect 436044 338660 436100 372316
rect 437612 372260 437668 372270
rect 437612 368900 437668 372204
rect 437612 368834 437668 368844
rect 440188 368788 440244 372428
rect 440188 368722 440244 368732
rect 436044 338594 436100 338604
rect 435932 93202 435988 93212
rect 437612 296996 437668 297006
rect 434252 79762 434308 79772
rect 435932 90804 435988 90814
rect 434476 79268 434532 79278
rect 434476 19684 434532 79212
rect 434476 19618 434532 19628
rect 435932 17892 435988 90748
rect 435932 17826 435988 17836
rect 436044 87556 436100 87566
rect 436044 16436 436100 87500
rect 436716 85988 436772 85998
rect 436268 85876 436324 85886
rect 436044 16370 436100 16380
rect 436156 84532 436212 84542
rect 436156 13188 436212 84476
rect 436268 16324 436324 85820
rect 436716 16548 436772 85932
rect 436716 16482 436772 16492
rect 436268 16258 436324 16268
rect 436156 13122 436212 13132
rect 435932 12628 435988 12638
rect 435932 480 435988 12572
rect 437612 4564 437668 296940
rect 439740 100884 439796 100894
rect 439404 94276 439460 94286
rect 437724 92484 437780 92494
rect 437724 19460 437780 92428
rect 439292 90916 439348 90926
rect 437724 19394 437780 19404
rect 437836 29428 437892 29438
rect 437836 14532 437892 29372
rect 438508 17668 438564 17678
rect 438508 15092 438564 17612
rect 438508 15026 438564 15036
rect 437836 14466 437892 14476
rect 439292 7924 439348 90860
rect 439404 17780 439460 94220
rect 439404 17714 439460 17724
rect 439516 80948 439572 80958
rect 439516 16660 439572 80892
rect 439516 16594 439572 16604
rect 439292 7858 439348 7868
rect 437612 4498 437668 4508
rect 437836 4228 437892 4238
rect 437836 480 437892 4172
rect 439740 480 439796 100828
rect 442652 94052 442708 389340
rect 446796 386372 446852 390460
rect 446796 386306 446852 386316
rect 443212 386148 443268 386158
rect 442764 373268 442820 373278
rect 442764 96628 442820 373212
rect 442876 371476 442932 371486
rect 442876 100660 442932 371420
rect 443100 371364 443156 371374
rect 442876 100594 442932 100604
rect 442988 370692 443044 370702
rect 442764 96562 442820 96572
rect 442876 97524 442932 97534
rect 442652 93986 442708 93996
rect 442764 94388 442820 94398
rect 442652 88564 442708 88574
rect 442428 80836 442484 80846
rect 441644 34468 441700 34478
rect 439964 22820 440020 22830
rect 439964 15876 440020 22764
rect 440076 22708 440132 22718
rect 440076 19236 440132 22652
rect 440076 19170 440132 19180
rect 439964 15810 440020 15820
rect 441644 480 441700 34412
rect 441868 15092 441924 15102
rect 441868 11060 441924 15036
rect 442428 13412 442484 80780
rect 442428 13346 442484 13356
rect 442652 13076 442708 88508
rect 442652 13010 442708 13020
rect 441868 10994 441924 11004
rect 442764 7140 442820 94332
rect 442876 19348 442932 97468
rect 442988 96740 443044 370636
rect 443100 99988 443156 371308
rect 443212 296548 443268 386092
rect 447244 384244 447300 395080
rect 451276 390516 451332 395080
rect 451276 390450 451332 390460
rect 455308 386260 455364 395080
rect 459340 389620 459396 395080
rect 459340 389554 459396 389564
rect 463372 389508 463428 395080
rect 463372 389442 463428 389452
rect 455308 386194 455364 386204
rect 447244 384178 447300 384188
rect 467404 384132 467460 395080
rect 467404 384066 467460 384076
rect 471436 384020 471492 395080
rect 475468 392196 475524 395080
rect 479500 393092 479556 395080
rect 479500 393026 479556 393036
rect 475468 392130 475524 392140
rect 483532 390964 483588 395080
rect 483532 390898 483588 390908
rect 487564 386036 487620 395080
rect 491596 387604 491652 395080
rect 491596 387538 491652 387548
rect 487564 385970 487620 385980
rect 495628 385924 495684 395080
rect 499660 389284 499716 395080
rect 499660 389218 499716 389228
rect 495628 385858 495684 385868
rect 503692 385812 503748 395080
rect 507724 387492 507780 395080
rect 511756 392532 511812 395080
rect 511756 392466 511812 392476
rect 507724 387426 507780 387436
rect 515788 387380 515844 395080
rect 519820 392420 519876 395080
rect 519820 392354 519876 392364
rect 523852 390852 523908 395080
rect 523852 390786 523908 390796
rect 515788 387314 515844 387324
rect 503692 385746 503748 385756
rect 527884 385700 527940 395080
rect 531916 389172 531972 395080
rect 535948 392308 536004 395080
rect 535948 392242 536004 392252
rect 531916 389106 531972 389116
rect 539980 387268 540036 395080
rect 544012 392644 544068 395080
rect 544012 392578 544068 392588
rect 539980 387202 540036 387212
rect 527884 385634 527940 385644
rect 471436 383954 471492 383964
rect 562604 380660 562660 595560
rect 562604 380594 562660 380604
rect 584668 378868 584724 595560
rect 587132 575428 587188 575438
rect 587132 385588 587188 575372
rect 587244 535780 587300 535790
rect 587244 388948 587300 535724
rect 590828 522564 590884 522574
rect 590492 469700 590548 469710
rect 587244 388882 587300 388892
rect 590380 403620 590436 403630
rect 587132 385522 587188 385532
rect 584668 378802 584724 378812
rect 544236 374612 544292 374622
rect 535052 373940 535108 373950
rect 535052 372484 535108 373884
rect 535052 372418 535108 372428
rect 544236 372372 544292 374556
rect 590380 373828 590436 403564
rect 590380 373762 590436 373772
rect 544236 372306 544292 372316
rect 590492 372148 590548 469644
rect 590716 456484 590772 456494
rect 590604 443268 590660 443278
rect 590604 375508 590660 443212
rect 590716 390740 590772 456428
rect 590828 394324 590884 522508
rect 591052 496132 591108 496142
rect 590828 394258 590884 394268
rect 590940 430164 590996 430174
rect 590716 390674 590772 390684
rect 590940 380548 590996 430108
rect 591052 394212 591108 496076
rect 591276 482916 591332 482926
rect 591052 394146 591108 394156
rect 591164 416836 591220 416846
rect 591164 383908 591220 416780
rect 591276 393988 591332 482860
rect 591276 393922 591332 393932
rect 591164 383842 591220 383852
rect 590940 380482 590996 380492
rect 590604 375442 590660 375452
rect 591052 373268 591108 373278
rect 590492 372082 590548 372092
rect 590604 373156 590660 373166
rect 590492 370692 590548 370702
rect 590492 311332 590548 370636
rect 590604 337652 590660 373100
rect 590828 373044 590884 373054
rect 590604 337586 590660 337596
rect 590716 371476 590772 371486
rect 590492 311266 590548 311276
rect 590716 298116 590772 371420
rect 590828 350980 590884 372988
rect 590828 350914 590884 350924
rect 590940 371364 590996 371374
rect 590940 324548 590996 371308
rect 591052 364196 591108 373212
rect 591052 364130 591108 364140
rect 590940 324482 590996 324492
rect 590716 298050 590772 298060
rect 443212 296482 443268 296492
rect 443996 296884 444052 296894
rect 443996 290668 444052 296828
rect 443996 290612 444276 290668
rect 443100 99922 443156 99932
rect 442988 96674 443044 96684
rect 443212 97748 443268 97758
rect 442876 19282 442932 19292
rect 442988 90020 443044 90030
rect 442988 8148 443044 89964
rect 443100 86324 443156 86334
rect 443100 12964 443156 86268
rect 443100 12898 443156 12908
rect 442988 8082 443044 8092
rect 442764 7074 442820 7084
rect 443212 4228 443268 97692
rect 444108 97636 444164 97646
rect 443436 94500 443492 94510
rect 443324 84084 443380 84094
rect 443324 12852 443380 84028
rect 443324 12786 443380 12796
rect 443436 4452 443492 94444
rect 443436 4386 443492 4396
rect 443548 90132 443604 90142
rect 443212 4162 443268 4172
rect 443548 480 443604 90076
rect 444108 7812 444164 97580
rect 444108 7746 444164 7756
rect 444220 4676 444276 290612
rect 587132 284676 587188 284686
rect 464492 19236 464548 19246
rect 460684 17556 460740 17566
rect 447356 15876 447412 15886
rect 444220 4610 444276 4620
rect 445452 7588 445508 7598
rect 445452 480 445508 7532
rect 447356 480 447412 15820
rect 458780 13412 458836 13422
rect 449260 8148 449316 8158
rect 449260 480 449316 8092
rect 456988 8036 457044 8046
rect 451164 6020 451220 6030
rect 451164 480 451220 5964
rect 454972 4900 455028 4910
rect 452956 480 453124 532
rect 454972 480 455028 4844
rect 456988 480 457044 7980
rect 458780 480 458836 13356
rect 460684 480 460740 17500
rect 462588 5908 462644 5918
rect 462588 480 462644 5852
rect 464492 480 464548 19180
rect 587132 17668 587188 284620
rect 587356 271460 587412 271470
rect 587244 178948 587300 178958
rect 587244 19460 587300 178892
rect 587244 19394 587300 19404
rect 587356 18228 587412 271404
rect 587580 218596 587636 218606
rect 587468 99652 587524 99662
rect 587468 19572 587524 99596
rect 587468 19506 587524 19516
rect 587356 18162 587412 18172
rect 587580 18004 587636 218540
rect 590828 165732 590884 165742
rect 587804 139300 587860 139310
rect 587804 18116 587860 139244
rect 590492 112868 590548 112878
rect 590268 60004 590324 60014
rect 590044 46788 590100 46798
rect 589820 33684 589876 33694
rect 589820 20020 589876 33628
rect 589820 19954 589876 19964
rect 590044 19684 590100 46732
rect 590268 20132 590324 59948
rect 590268 20066 590324 20076
rect 590044 19618 590100 19628
rect 587804 18050 587860 18060
rect 587580 17938 587636 17948
rect 590492 17892 590548 112812
rect 590828 20916 590884 165676
rect 590828 20850 590884 20860
rect 590940 152516 590996 152526
rect 590940 19908 590996 152460
rect 591052 126084 591108 126094
rect 591052 21028 591108 126028
rect 591276 86436 591332 86446
rect 591052 20962 591108 20972
rect 591164 73220 591220 73230
rect 590940 19842 590996 19852
rect 590492 17826 590548 17836
rect 591164 17780 591220 73164
rect 591276 20692 591332 86380
rect 591276 20626 591332 20636
rect 591276 20356 591332 20366
rect 591276 18452 591332 20300
rect 591276 18386 591332 18396
rect 591164 17714 591220 17724
rect 587132 17602 587188 17612
rect 487340 16772 487396 16782
rect 472108 13300 472164 13310
rect 468300 11284 468356 11294
rect 466396 4788 466452 4798
rect 466396 480 466452 4732
rect 468300 480 468356 11228
rect 470204 644 470260 654
rect 470204 480 470260 588
rect 472108 480 472164 13244
rect 481628 13188 481684 13198
rect 477820 4564 477876 4574
rect 475916 1764 475972 1774
rect 474012 644 474068 654
rect 474012 480 474068 588
rect 475916 480 475972 1708
rect 477820 480 477876 4508
rect 479724 4116 479780 4126
rect 479724 480 479780 4060
rect 481628 480 481684 13132
rect 483532 4676 483588 4686
rect 483532 480 483588 4620
rect 485548 644 485604 654
rect 485548 480 485604 588
rect 487340 480 487396 16716
rect 491148 16660 491204 16670
rect 489244 2884 489300 2894
rect 489244 480 489300 2828
rect 491148 480 491204 16604
rect 514108 16548 514164 16558
rect 508284 14868 508340 14878
rect 493052 13076 493108 13086
rect 493052 480 493108 13020
rect 498764 12964 498820 12974
rect 496860 4452 496916 4462
rect 494956 2660 495012 2670
rect 494956 480 495012 2604
rect 496860 480 496916 4396
rect 498764 480 498820 12908
rect 504476 12852 504532 12862
rect 500668 7924 500724 7934
rect 500668 480 500724 7868
rect 502572 2548 502628 2558
rect 502572 480 502628 2492
rect 504476 480 504532 12796
rect 506380 3444 506436 3454
rect 506380 480 506436 3388
rect 508284 480 508340 14812
rect 510188 12740 510244 12750
rect 510188 480 510244 12684
rect 512092 3444 512148 3454
rect 512092 480 512148 3388
rect 514108 480 514164 16492
rect 525420 16436 525476 16446
rect 519708 14756 519764 14766
rect 514220 8484 514276 8494
rect 514220 6804 514276 8428
rect 514220 6738 514276 6748
rect 517804 3444 517860 3454
rect 515900 1764 515956 1774
rect 515900 480 515956 1708
rect 517804 480 517860 3388
rect 519708 480 519764 14700
rect 521612 6804 521668 6814
rect 521612 480 521668 6748
rect 523516 4340 523572 4350
rect 523516 480 523572 4284
rect 525420 480 525476 16380
rect 538748 16324 538804 16334
rect 529228 14644 529284 14654
rect 527324 644 527380 654
rect 527324 480 527380 588
rect 529228 480 529284 14588
rect 531132 4340 531188 4350
rect 531132 480 531188 4284
rect 534940 3444 534996 3454
rect 533036 644 533092 654
rect 533036 480 533092 588
rect 534940 480 534996 3388
rect 536844 2772 536900 2782
rect 536844 480 536900 2716
rect 538748 480 538804 16268
rect 565404 16212 565460 16222
rect 546812 14532 546868 14542
rect 544460 11172 544516 11182
rect 540652 4004 540708 4014
rect 540652 480 540708 3948
rect 542668 1764 542724 1774
rect 542668 480 542724 1708
rect 544460 480 544516 11116
rect 546812 5012 546868 14476
rect 561596 11060 561652 11070
rect 552076 7812 552132 7822
rect 546812 4946 546868 4956
rect 550172 5012 550228 5022
rect 548268 4340 548324 4350
rect 546364 3892 546420 3902
rect 546364 480 546420 3836
rect 548268 480 548324 4284
rect 550172 480 550228 4956
rect 552076 480 552132 7756
rect 557788 3780 557844 3790
rect 555884 3444 555940 3454
rect 553980 644 554036 654
rect 553980 480 554036 588
rect 555884 480 555940 3388
rect 557788 480 557844 3724
rect 559692 3444 559748 3454
rect 559692 480 559748 3388
rect 561596 480 561652 11004
rect 563500 10948 563556 10958
rect 563500 480 563556 10892
rect 565404 480 565460 16156
rect 567308 16100 567364 16110
rect 567308 480 567364 16044
rect 578732 15988 578788 15998
rect 569212 14420 569268 14430
rect 569212 480 569268 14364
rect 576828 14308 576884 14318
rect 574924 6804 574980 6814
rect 573020 4228 573076 4238
rect 571228 3444 571284 3454
rect 571228 480 571284 3388
rect 573020 480 573076 4172
rect 574924 480 574980 6748
rect 576828 480 576884 14252
rect 578732 480 578788 15932
rect 584444 12628 584500 12638
rect 580636 7700 580692 7710
rect 580636 480 580692 7644
rect 582540 4228 582596 4238
rect 582540 480 582596 4172
rect 584444 480 584500 12572
rect 422604 392 422856 480
rect 424508 392 424760 480
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418824 -960 419048 392
rect 420728 -960 420952 392
rect 422632 -960 422856 392
rect 424536 -960 424760 392
rect 426440 392 426692 480
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432124 392 432376 480
rect 434028 392 434280 480
rect 435932 392 436184 480
rect 437836 392 438088 480
rect 439740 392 439992 480
rect 441644 392 441896 480
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 447356 392 447608 480
rect 449260 392 449512 480
rect 451164 392 451416 480
rect 432152 -960 432376 392
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 447384 -960 447608 392
rect 449288 -960 449512 392
rect 451192 -960 451416 392
rect 452956 476 453320 480
rect 452956 196 453012 476
rect 453068 392 453320 476
rect 454972 392 455224 480
rect 452956 130 453012 140
rect 453096 -960 453320 392
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 460684 392 460936 480
rect 462588 392 462840 480
rect 464492 392 464744 480
rect 466396 392 466648 480
rect 468300 392 468552 480
rect 470204 392 470456 480
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 475916 392 476168 480
rect 477820 392 478072 480
rect 479724 392 479976 480
rect 481628 392 481880 480
rect 483532 392 483784 480
rect 458808 -960 459032 392
rect 460712 -960 460936 392
rect 462616 -960 462840 392
rect 464520 -960 464744 392
rect 466424 -960 466648 392
rect 468328 -960 468552 392
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475944 -960 476168 392
rect 477848 -960 478072 392
rect 479752 -960 479976 392
rect 481656 -960 481880 392
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487340 392 487592 480
rect 489244 392 489496 480
rect 491148 392 491400 480
rect 493052 392 493304 480
rect 494956 392 495208 480
rect 496860 392 497112 480
rect 498764 392 499016 480
rect 500668 392 500920 480
rect 502572 392 502824 480
rect 504476 392 504728 480
rect 506380 392 506632 480
rect 508284 392 508536 480
rect 510188 392 510440 480
rect 512092 392 512344 480
rect 487368 -960 487592 392
rect 489272 -960 489496 392
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 494984 -960 495208 392
rect 496888 -960 497112 392
rect 498792 -960 499016 392
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504504 -960 504728 392
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 510216 -960 510440 392
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 517804 392 518056 480
rect 519708 392 519960 480
rect 521612 392 521864 480
rect 523516 392 523768 480
rect 525420 392 525672 480
rect 527324 392 527576 480
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 533036 392 533288 480
rect 534940 392 535192 480
rect 536844 392 537096 480
rect 538748 392 539000 480
rect 540652 392 540904 480
rect 515928 -960 516152 392
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 521640 -960 521864 392
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 533064 -960 533288 392
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 538776 -960 539000 392
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 550172 392 550424 480
rect 552076 392 552328 480
rect 553980 392 554232 480
rect 555884 392 556136 480
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 563500 392 563752 480
rect 565404 392 565656 480
rect 567308 392 567560 480
rect 569212 392 569464 480
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 550200 -960 550424 392
rect 552104 -960 552328 392
rect 554008 -960 554232 392
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 567336 -960 567560 392
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 574924 392 575176 480
rect 576828 392 577080 480
rect 578732 392 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 573048 -960 573272 392
rect 574952 -960 575176 392
rect 576856 -960 577080 392
rect 578760 -960 578984 392
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 4844 416668 4900 416724
rect 4844 394380 4900 394436
rect 4956 403228 5012 403284
rect 19180 590940 19236 590996
rect 33068 590940 33124 590996
rect 55132 590828 55188 590884
rect 77308 590716 77364 590772
rect 99260 590604 99316 590660
rect 143388 590492 143444 590548
rect 121324 577276 121380 577332
rect 162092 590156 162148 590212
rect 29260 577164 29316 577220
rect 28476 577052 28532 577108
rect 165452 590156 165508 590212
rect 162092 576044 162148 576100
rect 169708 577276 169764 577332
rect 193228 583772 193284 583828
rect 187516 577276 187572 577332
rect 188076 579292 188132 579348
rect 169708 575932 169764 575988
rect 209580 583772 209636 583828
rect 225932 590156 225988 590212
rect 193228 579292 193284 579348
rect 231644 590156 231700 590212
rect 242732 590492 242788 590548
rect 225932 576268 225988 576324
rect 188076 575820 188132 575876
rect 253708 590492 253764 590548
rect 242732 575596 242788 575652
rect 268716 582988 268772 583044
rect 275772 582988 275828 583044
rect 295596 587916 295652 587972
rect 268716 575484 268772 575540
rect 292236 581308 292292 581364
rect 317548 590156 317604 590212
rect 297836 587916 297892 587972
rect 314188 587916 314244 587972
rect 319900 590156 319956 590212
rect 336812 590492 336868 590548
rect 317548 587916 317604 587972
rect 295596 581308 295652 581364
rect 310828 579516 310884 579572
rect 314076 579516 314132 579572
rect 310828 577164 310884 577220
rect 341964 590492 342020 590548
rect 364252 590492 364308 590548
rect 380492 590492 380548 590548
rect 386092 581308 386148 581364
rect 394828 581308 394884 581364
rect 380492 577836 380548 577892
rect 383068 577836 383124 577892
rect 336812 577052 336868 577108
rect 292236 575372 292292 575428
rect 540764 591052 540820 591108
rect 518700 590940 518756 590996
rect 496636 590828 496692 590884
rect 474572 590716 474628 590772
rect 452508 590604 452564 590660
rect 430444 590492 430500 590548
rect 408268 575596 408324 575652
rect 394828 575484 394884 575540
rect 383068 575372 383124 575428
rect 29260 575036 29316 575092
rect 28476 574476 28532 574532
rect 19180 380492 19236 380548
rect 27692 389676 27748 389732
rect 11004 378812 11060 378868
rect 30268 394492 30324 394548
rect 30156 393148 30212 393204
rect 28476 393036 28532 393092
rect 30268 392476 30324 392532
rect 35980 392364 36036 392420
rect 37772 392476 37828 392532
rect 31948 392252 32004 392308
rect 28476 389788 28532 389844
rect 28588 389676 28644 389732
rect 30268 389340 30324 389396
rect 31052 389676 31108 389732
rect 28588 384748 28644 384804
rect 35084 389676 35140 389732
rect 34412 389340 34468 389396
rect 31052 384076 31108 384132
rect 33404 384636 33460 384692
rect 33404 381836 33460 381892
rect 33516 382956 33572 383012
rect 37772 389676 37828 389732
rect 35084 387884 35140 387940
rect 35196 389452 35252 389508
rect 40236 389676 40292 389732
rect 40012 387212 40068 387268
rect 35196 386316 35252 386372
rect 39004 386316 39060 386372
rect 34412 381388 34468 381444
rect 36764 384076 36820 384132
rect 33516 379708 33572 379764
rect 27916 378924 27972 378980
rect 27692 377916 27748 377972
rect 28700 377916 28756 377972
rect 37772 381836 37828 381892
rect 36876 381388 36932 381444
rect 36876 379484 36932 379540
rect 4956 377132 5012 377188
rect 36876 377356 36932 377412
rect 36876 375900 36932 375956
rect 28700 375676 28756 375732
rect 40348 385532 40404 385588
rect 41132 387884 41188 387940
rect 44044 387324 44100 387380
rect 41132 382172 41188 382228
rect 47852 385532 47908 385588
rect 39004 381388 39060 381444
rect 42812 381388 42868 381444
rect 42028 379484 42084 379540
rect 42028 377356 42084 377412
rect 37772 375788 37828 375844
rect 36988 374220 37044 374276
rect 46956 379260 47012 379316
rect 46956 376236 47012 376292
rect 52108 392588 52164 392644
rect 56140 392476 56196 392532
rect 57036 392364 57092 392420
rect 60172 392364 60228 392420
rect 63868 392588 63924 392644
rect 57036 390796 57092 390852
rect 60396 392252 60452 392308
rect 64204 391468 64260 391524
rect 65660 391468 65716 391524
rect 63868 390908 63924 390964
rect 60396 388892 60452 388948
rect 70476 392476 70532 392532
rect 72268 392252 72324 392308
rect 70476 387436 70532 387492
rect 80332 389004 80388 389060
rect 88396 387660 88452 387716
rect 84364 387548 84420 387604
rect 76300 385756 76356 385812
rect 68236 385644 68292 385700
rect 65660 385532 65716 385588
rect 96460 393036 96516 393092
rect 100492 392476 100548 392532
rect 112588 391020 112644 391076
rect 120652 389228 120708 389284
rect 116620 389116 116676 389172
rect 108556 385980 108612 386036
rect 104524 385868 104580 385924
rect 128716 392924 128772 392980
rect 136780 392700 136836 392756
rect 140812 392588 140868 392644
rect 132748 391468 132804 391524
rect 136108 391468 136164 391524
rect 144844 391132 144900 391188
rect 148876 387772 148932 387828
rect 152236 394380 152292 394436
rect 136108 386092 136164 386148
rect 124684 384300 124740 384356
rect 92428 384188 92484 384244
rect 48076 384076 48132 384132
rect 48636 382172 48692 382228
rect 48636 381276 48692 381332
rect 50428 381276 50484 381332
rect 50428 378028 50484 378084
rect 57036 377916 57092 377972
rect 47852 376124 47908 376180
rect 48636 377356 48692 377412
rect 48636 374332 48692 374388
rect 50428 376236 50484 376292
rect 57036 376012 57092 376068
rect 62188 376124 62244 376180
rect 62188 374444 62244 374500
rect 151004 375900 151060 375956
rect 149324 374332 149380 374388
rect 151004 374332 151060 374388
rect 151116 374444 151172 374500
rect 50428 372988 50484 373044
rect 42812 372428 42868 372484
rect 149548 370636 149604 370692
rect 151116 372540 151172 372596
rect 151228 369628 151284 369684
rect 151452 370636 151508 370692
rect 151452 367948 151508 368004
rect 151228 364476 151284 364532
rect 156940 394268 156996 394324
rect 160972 392812 161028 392868
rect 152908 391244 152964 391300
rect 164556 392364 164612 392420
rect 165004 391580 165060 391636
rect 164556 390684 164612 390740
rect 169036 390572 169092 390628
rect 173068 387884 173124 387940
rect 176316 391580 176372 391636
rect 185164 392364 185220 392420
rect 186396 392924 186452 392980
rect 177100 389340 177156 389396
rect 180124 390796 180180 390852
rect 176316 386204 176372 386260
rect 186396 391356 186452 391412
rect 188972 392252 189028 392308
rect 187292 390908 187348 390964
rect 183708 387324 183764 387380
rect 181468 387100 181524 387156
rect 181916 387212 181972 387268
rect 185500 384076 185556 384132
rect 189196 392252 189252 392308
rect 188972 390348 189028 390404
rect 192668 390684 192724 390740
rect 189084 388892 189140 388948
rect 190876 387436 190932 387492
rect 193228 390684 193284 390740
rect 194908 392476 194964 392532
rect 197260 388892 197316 388948
rect 198044 390348 198100 390404
rect 194908 386316 194964 386372
rect 196252 385644 196308 385700
rect 194460 385532 194516 385588
rect 201292 387324 201348 387380
rect 201628 389004 201684 389060
rect 199836 385756 199892 385812
rect 205212 387660 205268 387716
rect 203420 387548 203476 387604
rect 205324 385532 205380 385588
rect 208796 393148 208852 393204
rect 207004 384188 207060 384244
rect 210028 385644 210084 385700
rect 210588 386316 210644 386372
rect 212380 385868 212436 385924
rect 215964 391020 216020 391076
rect 213388 385756 213444 385812
rect 214172 385980 214228 386036
rect 223468 392700 223524 392756
rect 221452 390796 221508 390852
rect 223132 391356 223188 391412
rect 219548 389228 219604 389284
rect 217420 387436 217476 387492
rect 217756 389116 217812 389172
rect 221340 384300 221396 384356
rect 229516 392700 229572 392756
rect 225484 391468 225540 391524
rect 228508 392588 228564 392644
rect 223468 386316 223524 386372
rect 226716 386316 226772 386372
rect 224924 386092 224980 386148
rect 233548 392476 233604 392532
rect 235676 394268 235732 394324
rect 233884 391244 233940 391300
rect 230300 391132 230356 391188
rect 232092 387772 232148 387828
rect 237468 392812 237524 392868
rect 237580 392588 237636 392644
rect 238588 392700 238644 392756
rect 238588 389004 238644 389060
rect 241052 390572 241108 390628
rect 239260 386204 239316 386260
rect 241612 390572 241668 390628
rect 241948 392364 242004 392420
rect 245644 392364 245700 392420
rect 246988 392252 247044 392308
rect 244636 389340 244692 389396
rect 241948 385868 242004 385924
rect 242844 387884 242900 387940
rect 246428 387212 246484 387268
rect 249676 392252 249732 392308
rect 251804 390684 251860 390740
rect 246988 386316 247044 386372
rect 250012 386316 250068 386372
rect 248220 385868 248276 385924
rect 253708 389116 253764 389172
rect 253596 388892 253652 388948
rect 257740 388892 257796 388948
rect 260316 392588 260372 392644
rect 255388 387324 255444 387380
rect 263788 392476 263844 392532
rect 265468 392364 265524 392420
rect 263788 390684 263844 390740
rect 264348 390796 264404 390852
rect 261772 389228 261828 389284
rect 260316 385868 260372 385924
rect 262556 387436 262612 387492
rect 260764 385756 260820 385812
rect 258972 385644 259028 385700
rect 257180 385532 257236 385588
rect 265468 387212 265524 387268
rect 265804 385532 265860 385588
rect 266140 390908 266196 390964
rect 269724 390684 269780 390740
rect 267932 389004 267988 389060
rect 270396 392252 270452 392308
rect 273868 392252 273924 392308
rect 270396 387996 270452 388052
rect 273308 390572 273364 390628
rect 269836 385644 269892 385700
rect 271516 385868 271572 385924
rect 276892 387996 276948 388052
rect 275100 387212 275156 387268
rect 277900 385756 277956 385812
rect 278684 389116 278740 389172
rect 280476 388892 280532 388948
rect 281932 387212 281988 387268
rect 282268 389228 282324 389284
rect 285964 386428 286020 386484
rect 287644 392252 287700 392308
rect 285852 385644 285908 385700
rect 284060 385532 284116 385588
rect 289996 392252 290052 392308
rect 291228 387212 291284 387268
rect 289436 385756 289492 385812
rect 293020 386428 293076 386484
rect 294028 386316 294084 386372
rect 294812 392252 294868 392308
rect 296604 386316 296660 386372
rect 301980 390684 302036 390740
rect 300188 387996 300244 388052
rect 306124 390684 306180 390740
rect 305564 390572 305620 390628
rect 302092 387996 302148 388052
rect 303772 389676 303828 389732
rect 310156 389676 310212 389732
rect 310940 392700 310996 392756
rect 309148 385644 309204 385700
rect 307356 385532 307412 385588
rect 312732 392364 312788 392420
rect 314188 390572 314244 390628
rect 314524 392476 314580 392532
rect 318108 392252 318164 392308
rect 316316 387212 316372 387268
rect 321692 390572 321748 390628
rect 318220 385532 318276 385588
rect 319900 385532 319956 385588
rect 326284 392700 326340 392756
rect 325276 392588 325332 392644
rect 322252 385644 322308 385700
rect 323484 387324 323540 387380
rect 334348 392476 334404 392532
rect 334460 392700 334516 392756
rect 330316 392364 330372 392420
rect 334236 392364 334292 392420
rect 332444 389004 332500 389060
rect 328860 387436 328916 387492
rect 327068 386316 327124 386372
rect 330652 385644 330708 385700
rect 334460 387324 334516 387380
rect 336028 390908 336084 390964
rect 336028 386316 336084 386372
rect 337820 390796 337876 390852
rect 336028 385868 336084 385924
rect 342412 392252 342468 392308
rect 343532 392476 343588 392532
rect 338380 387212 338436 387268
rect 340956 388220 341012 388276
rect 339612 385980 339668 386036
rect 340956 385532 341012 385588
rect 341404 387212 341460 387268
rect 346444 388220 346500 388276
rect 348572 391244 348628 391300
rect 344540 387324 344596 387380
rect 344540 385980 344596 386036
rect 344988 385980 345044 386036
rect 343532 385868 343588 385924
rect 343196 385756 343252 385812
rect 346780 385532 346836 385588
rect 354508 392700 354564 392756
rect 358540 392588 358596 392644
rect 359548 392588 359604 392644
rect 355292 392252 355348 392308
rect 350476 390572 350532 390628
rect 351820 390572 351876 390628
rect 351036 389116 351092 389172
rect 350364 386316 350420 386372
rect 351820 386316 351876 386372
rect 352828 388892 352884 388948
rect 351036 385644 351092 385700
rect 359324 390684 359380 390740
rect 355292 385980 355348 386036
rect 355740 386316 355796 386372
rect 353948 385868 354004 385924
rect 357532 385644 357588 385700
rect 362572 390908 362628 390964
rect 362796 391020 362852 391076
rect 359548 386316 359604 386372
rect 361116 384748 361172 384804
rect 366156 387884 366212 387940
rect 362796 384748 362852 384804
rect 362908 386204 362964 386260
rect 366604 387436 366660 387492
rect 367948 391132 368004 391188
rect 366156 385756 366212 385812
rect 366492 386316 366548 386372
rect 364700 384188 364756 384244
rect 370076 389564 370132 389620
rect 367948 386204 368004 386260
rect 368284 386204 368340 386260
rect 370636 389116 370692 389172
rect 371868 389452 371924 389508
rect 378700 392364 378756 392420
rect 381388 393036 381444 393092
rect 374668 389004 374724 389060
rect 378700 392140 378756 392196
rect 374556 387660 374612 387716
rect 374556 385868 374612 385924
rect 377244 386092 377300 386148
rect 373660 384076 373716 384132
rect 375452 383964 375508 384020
rect 380828 390908 380884 390964
rect 378700 386092 378756 386148
rect 379036 386092 379092 386148
rect 382732 392476 382788 392532
rect 386764 390796 386820 390852
rect 387996 389228 388052 389284
rect 381388 386092 381444 386148
rect 384412 387548 384468 387604
rect 382620 385980 382676 386036
rect 386204 385868 386260 385924
rect 390572 387772 390628 387828
rect 389788 385756 389844 385812
rect 393372 392476 393428 392532
rect 390796 387324 390852 387380
rect 391580 387436 391636 387492
rect 390572 385644 390628 385700
rect 396956 392364 397012 392420
rect 394828 387212 394884 387268
rect 395164 387324 395220 387380
rect 398748 390796 398804 390852
rect 402892 392252 402948 392308
rect 404124 392252 404180 392308
rect 398860 387884 398916 387940
rect 401436 391468 401492 391524
rect 400540 385644 400596 385700
rect 401436 385532 401492 385588
rect 402332 389116 402388 389172
rect 406924 391468 406980 391524
rect 407708 391356 407764 391412
rect 405916 387212 405972 387268
rect 410956 391244 411012 391300
rect 414988 390572 415044 390628
rect 419020 388892 419076 388948
rect 423052 387660 423108 387716
rect 424172 393932 424228 393988
rect 163772 380492 163828 380548
rect 154588 376012 154644 376068
rect 152908 375788 152964 375844
rect 152908 372988 152964 373044
rect 154252 375676 154308 375732
rect 152796 372428 152852 372484
rect 154588 374444 154644 374500
rect 157948 374444 158004 374500
rect 154364 374332 154420 374388
rect 156156 374220 156212 374276
rect 153020 369628 153076 369684
rect 152908 364364 152964 364420
rect 157948 371308 158004 371364
rect 159516 372876 159572 372932
rect 156380 369628 156436 369684
rect 154812 369180 154868 369236
rect 159516 369180 159572 369236
rect 154700 367948 154756 368004
rect 157052 367948 157108 368004
rect 153020 363020 153076 363076
rect 154476 364476 154532 364532
rect 154588 364364 154644 364420
rect 154588 362684 154644 362740
rect 154700 354508 154756 354564
rect 162876 371084 162932 371140
rect 159628 368844 159684 368900
rect 160524 369516 160580 369572
rect 159628 365372 159684 365428
rect 160412 367836 160468 367892
rect 158060 362684 158116 362740
rect 158060 358764 158116 358820
rect 157052 352716 157108 352772
rect 158844 354396 158900 354452
rect 158844 347788 158900 347844
rect 162876 364476 162932 364532
rect 162092 363020 162148 363076
rect 160860 352716 160916 352772
rect 160860 348684 160916 348740
rect 160524 257068 160580 257124
rect 160412 230188 160468 230244
rect 152236 58828 152292 58884
rect 153692 78988 153748 79044
rect 150332 40012 150388 40068
rect 4172 36876 4228 36932
rect 3500 23436 3556 23492
rect 3500 17612 3556 17668
rect 162204 358764 162260 358820
rect 162204 69580 162260 69636
rect 162316 347676 162372 347732
rect 162428 257068 162484 257124
rect 162652 230188 162708 230244
rect 162652 68684 162708 68740
rect 162428 67788 162484 67844
rect 162316 66892 162372 66948
rect 162092 65996 162148 66052
rect 172172 378924 172228 378980
rect 166348 378812 166404 378868
rect 166012 377132 166068 377188
rect 163996 375564 164052 375620
rect 164556 374556 164612 374612
rect 164332 373996 164388 374052
rect 164108 373884 164164 373940
rect 164220 372316 164276 372372
rect 164220 65100 164276 65156
rect 164108 63308 164164 63364
rect 164556 64204 164612 64260
rect 164332 62412 164388 62468
rect 163996 61516 164052 61572
rect 163772 60620 163828 60676
rect 166796 368844 166852 368900
rect 166796 366156 166852 366212
rect 167244 365372 167300 365428
rect 167244 359548 167300 359604
rect 167580 364476 167636 364532
rect 171388 359436 171444 359492
rect 167580 354396 167636 354452
rect 170492 354396 170548 354452
rect 167132 348684 167188 348740
rect 167132 346108 167188 346164
rect 171388 349468 171444 349524
rect 170492 324604 170548 324660
rect 171612 300636 171668 300692
rect 170940 78988 170996 79044
rect 172396 366156 172452 366212
rect 172172 79884 172228 79940
rect 172284 298732 172340 298788
rect 420924 362796 420980 362852
rect 172396 243628 172452 243684
rect 173852 349468 173908 349524
rect 173964 345660 174020 345716
rect 420924 337708 420980 337764
rect 173852 99036 173908 99092
rect 173964 324604 174020 324660
rect 173628 93324 173684 93380
rect 172956 78988 173012 79044
rect 419132 333452 419188 333508
rect 418348 314188 418404 314244
rect 378364 308252 378420 308308
rect 189308 305676 189364 305732
rect 185724 305564 185780 305620
rect 183484 305340 183540 305396
rect 183036 305228 183092 305284
rect 182588 305116 182644 305172
rect 177212 305004 177268 305060
rect 176204 300636 176260 300692
rect 174300 299852 174356 299908
rect 174076 105196 174132 105252
rect 174188 243628 174244 243684
rect 174188 85148 174244 85204
rect 173964 83692 174020 83748
rect 179004 304892 179060 304948
rect 178108 303548 178164 303604
rect 177660 301532 177716 301588
rect 178556 303436 178612 303492
rect 180348 303884 180404 303940
rect 179900 303212 179956 303268
rect 179452 301644 179508 301700
rect 180796 303772 180852 303828
rect 181244 303660 181300 303716
rect 182140 301980 182196 302036
rect 181692 301868 181748 301924
rect 184380 303324 184436 303380
rect 183932 301756 183988 301812
rect 187964 305452 188020 305508
rect 186620 303996 186676 304052
rect 186172 302204 186228 302260
rect 187068 303100 187124 303156
rect 187516 299964 187572 300020
rect 188860 302316 188916 302372
rect 188412 301420 188468 301476
rect 191100 305004 191156 305060
rect 189756 304780 189812 304836
rect 190204 302092 190260 302148
rect 191996 303548 192052 303604
rect 192892 304892 192948 304948
rect 192444 303436 192500 303492
rect 192892 304668 192948 304724
rect 192444 303100 192500 303156
rect 191996 302988 192052 303044
rect 191548 301532 191604 301588
rect 191772 302876 191828 302932
rect 191100 299068 191156 299124
rect 193788 303884 193844 303940
rect 194236 303772 194292 303828
rect 194684 303660 194740 303716
rect 193340 301644 193396 301700
rect 193564 303548 193620 303604
rect 193788 303436 193844 303492
rect 196924 305340 196980 305396
rect 196476 305228 196532 305284
rect 196028 305116 196084 305172
rect 195580 301980 195636 302036
rect 196028 304556 196084 304612
rect 195132 301868 195188 301924
rect 195580 301644 195636 301700
rect 194684 301532 194740 301588
rect 194236 301196 194292 301252
rect 195132 301308 195188 301364
rect 197820 303212 197876 303268
rect 197932 303660 197988 303716
rect 197260 301756 197316 301812
rect 197372 301980 197428 302036
rect 198716 305564 198772 305620
rect 198268 303324 198324 303380
rect 198492 305340 198548 305396
rect 198716 305116 198772 305172
rect 199612 303996 199668 304052
rect 199724 305004 199780 305060
rect 199052 302204 199108 302260
rect 199164 303212 199220 303268
rect 200060 304444 200116 304500
rect 200060 303772 200116 303828
rect 200508 299964 200564 300020
rect 200844 301756 200900 301812
rect 201404 305452 201460 305508
rect 201404 305228 201460 305284
rect 200956 301420 201012 301476
rect 201292 301868 201348 301924
rect 202300 305676 202356 305732
rect 202748 304780 202804 304836
rect 203084 305452 203140 305508
rect 201852 302316 201908 302372
rect 202748 303996 202804 304052
rect 202300 301420 202356 301476
rect 201852 299180 201908 299236
rect 204092 302988 204148 303044
rect 204316 303884 204372 303940
rect 203644 302876 203700 302932
rect 203196 302092 203252 302148
rect 203644 302652 203700 302708
rect 204540 303100 204596 303156
rect 204764 304892 204820 304948
rect 204540 302876 204596 302932
rect 204988 304668 205044 304724
rect 205436 303548 205492 303604
rect 204764 298956 204820 299012
rect 204988 303324 205044 303380
rect 205436 303100 205492 303156
rect 205884 301196 205940 301252
rect 206108 305564 206164 305620
rect 206332 303436 206388 303492
rect 206556 305676 206612 305732
rect 206668 301532 206724 301588
rect 206780 302092 206836 302148
rect 208124 304556 208180 304612
rect 209468 305340 209524 305396
rect 209804 305340 209860 305396
rect 209468 304780 209524 304836
rect 209020 303660 209076 303716
rect 209132 304668 209188 304724
rect 208572 301980 208628 302036
rect 207676 301644 207732 301700
rect 208124 301644 208180 301700
rect 207228 301308 207284 301364
rect 207228 299292 207284 299348
rect 208572 300748 208628 300804
rect 209916 305116 209972 305172
rect 211260 305004 211316 305060
rect 210812 303772 210868 303828
rect 211260 304556 211316 304612
rect 210364 303212 210420 303268
rect 210476 303436 210532 303492
rect 210812 303212 210868 303268
rect 211708 301756 211764 301812
rect 211932 302540 211988 302596
rect 212604 305228 212660 305284
rect 213500 305452 213556 305508
rect 213052 303996 213108 304052
rect 212156 301868 212212 301924
rect 212380 303548 212436 303604
rect 213948 302652 214004 302708
rect 214172 304108 214228 304164
rect 213500 302428 213556 302484
rect 212604 299516 212660 299572
rect 213052 298844 213108 298900
rect 214396 303884 214452 303940
rect 214620 304220 214676 304276
rect 215292 303100 215348 303156
rect 215516 305452 215572 305508
rect 214844 302876 214900 302932
rect 214844 301868 214900 301924
rect 216636 305676 216692 305732
rect 216188 305564 216244 305620
rect 215740 303324 215796 303380
rect 215964 305004 216020 305060
rect 216188 303884 216244 303940
rect 216636 303772 216692 303828
rect 217084 302092 217140 302148
rect 217084 301756 217140 301812
rect 217532 301644 217588 301700
rect 217756 303324 217812 303380
rect 219324 305340 219380 305396
rect 218876 304780 218932 304836
rect 218428 304668 218484 304724
rect 219324 303996 219380 304052
rect 218876 302204 218932 302260
rect 217980 300748 218036 300804
rect 218428 300748 218484 300804
rect 217980 299404 218036 299460
rect 220668 304556 220724 304612
rect 220220 303436 220276 303492
rect 219772 303212 219828 303268
rect 221564 303548 221620 303604
rect 221116 302540 221172 302596
rect 221564 303212 221620 303268
rect 220668 302092 220724 302148
rect 220220 301980 220276 302036
rect 219772 301644 219828 301700
rect 221116 300972 221172 301028
rect 221788 302428 221844 302484
rect 222012 305116 222068 305172
rect 222908 304220 222964 304276
rect 222460 304108 222516 304164
rect 222460 303436 222516 303492
rect 223356 301868 223412 301924
rect 223692 305788 223748 305844
rect 222908 300860 222964 300916
rect 223356 299516 223412 299572
rect 223804 305452 223860 305508
rect 224252 303884 224308 303940
rect 224476 305228 224532 305284
rect 224700 305004 224756 305060
rect 224700 303884 224756 303940
rect 225148 303772 225204 303828
rect 225372 304220 225428 304276
rect 225596 301756 225652 301812
rect 225820 304332 225876 304388
rect 226044 303324 226100 303380
rect 226268 304444 226324 304500
rect 226492 302204 226548 302260
rect 226716 304556 226772 304612
rect 226940 303996 226996 304052
rect 226940 302428 226996 302484
rect 228284 302092 228340 302148
rect 228396 305004 228452 305060
rect 227836 301980 227892 302036
rect 228284 301868 228340 301924
rect 227388 301644 227444 301700
rect 227836 301756 227892 301812
rect 227388 301308 227444 301364
rect 228732 303212 228788 303268
rect 229628 305116 229684 305172
rect 229180 300972 229236 301028
rect 229628 303660 229684 303716
rect 228396 299852 228452 299908
rect 228732 300748 228788 300804
rect 229180 300748 229236 300804
rect 229964 303548 230020 303604
rect 230076 303436 230132 303492
rect 230972 305228 231028 305284
rect 230524 300860 230580 300916
rect 230748 304780 230804 304836
rect 231420 303884 231476 303940
rect 231644 305340 231700 305396
rect 230972 301980 231028 302036
rect 232764 304444 232820 304500
rect 232316 304332 232372 304388
rect 231868 304220 231924 304276
rect 232316 303324 232372 303380
rect 231868 300748 231924 300804
rect 232876 302428 232932 302484
rect 232988 305564 233044 305620
rect 233660 304556 233716 304612
rect 233212 304220 233268 304276
rect 233660 304108 233716 304164
rect 234108 301308 234164 301364
rect 234332 305452 234388 305508
rect 234556 301756 234612 301812
rect 234780 305116 234836 305172
rect 234892 301868 234948 301924
rect 235004 303772 235060 303828
rect 235452 303660 235508 303716
rect 236348 304780 236404 304836
rect 236572 305228 236628 305284
rect 235564 303548 235620 303604
rect 235900 303996 235956 304052
rect 235452 303436 235508 303492
rect 236684 303884 236740 303940
rect 237244 305340 237300 305396
rect 236796 301980 236852 302036
rect 237244 301196 237300 301252
rect 238588 305564 238644 305620
rect 239036 305452 239092 305508
rect 239484 305116 239540 305172
rect 239932 303772 239988 303828
rect 240156 304556 240212 304612
rect 238140 303324 238196 303380
rect 237692 300748 237748 300804
rect 238140 302764 238196 302820
rect 237692 299516 237748 299572
rect 238588 302316 238644 302372
rect 239036 302204 239092 302260
rect 239484 302092 239540 302148
rect 241276 305228 241332 305284
rect 240828 303996 240884 304052
rect 241276 304668 241332 304724
rect 240380 303436 240436 303492
rect 240380 301980 240436 302036
rect 240828 301868 240884 301924
rect 241724 303884 241780 303940
rect 241836 304780 241892 304836
rect 242620 302316 242676 302372
rect 243068 303100 243124 303156
rect 242732 302204 242788 302260
rect 242956 302540 243012 302596
rect 242172 301196 242228 301252
rect 242172 300748 242228 300804
rect 243964 304556 244020 304612
rect 243964 304332 244020 304388
rect 243180 302092 243236 302148
rect 243516 303212 243572 303268
rect 244076 301980 244132 302036
rect 244412 304444 244468 304500
rect 245756 304780 245812 304836
rect 245308 304668 245364 304724
rect 247548 304444 247604 304500
rect 247100 304332 247156 304388
rect 246652 303212 246708 303268
rect 246204 303100 246260 303156
rect 247548 303100 247604 303156
rect 245308 302988 245364 303044
rect 244524 301868 244580 301924
rect 244860 302316 244916 302372
rect 245756 302204 245812 302260
rect 246204 302092 246260 302148
rect 247100 301196 247156 301252
rect 246876 298956 246932 299012
rect 247660 302316 247716 302372
rect 247996 303212 248052 303268
rect 248444 302988 248500 303044
rect 248892 302204 248948 302260
rect 249228 303772 249284 303828
rect 248444 300972 248500 301028
rect 249340 302092 249396 302148
rect 249676 303996 249732 304052
rect 250236 303212 250292 303268
rect 249788 303100 249844 303156
rect 250684 300972 250740 301028
rect 250908 303884 250964 303940
rect 250236 300860 250292 300916
rect 249788 300748 249844 300804
rect 251580 303996 251636 304052
rect 251132 303772 251188 303828
rect 251132 301084 251188 301140
rect 251580 300972 251636 301028
rect 252028 300748 252084 300804
rect 252364 300860 252420 300916
rect 252476 303996 252532 304052
rect 253820 303996 253876 304052
rect 252588 303884 252644 303940
rect 252924 303884 252980 303940
rect 252588 301196 252644 301252
rect 252588 300860 252644 300916
rect 254268 303884 254324 303940
rect 253372 303772 253428 303828
rect 254716 303772 254772 303828
rect 255164 302876 255220 302932
rect 254716 302764 254772 302820
rect 254268 302652 254324 302708
rect 256508 302876 256564 302932
rect 256060 302764 256116 302820
rect 255612 302652 255668 302708
rect 256284 302652 256340 302708
rect 260540 300748 260596 300804
rect 272188 305676 272244 305732
rect 271740 305452 271796 305508
rect 272636 305116 272692 305172
rect 272972 305340 273028 305396
rect 271292 304892 271348 304948
rect 207676 298732 207732 298788
rect 196924 298620 196980 298676
rect 190652 298508 190708 298564
rect 196476 298396 196532 298452
rect 184828 298284 184884 298340
rect 185276 298284 185332 298340
rect 255612 298284 255668 298340
rect 260092 298284 260148 298340
rect 191100 101948 191156 102004
rect 183036 101836 183092 101892
rect 181020 101724 181076 101780
rect 178332 101612 178388 101668
rect 174972 100156 175028 100212
rect 177772 99036 177828 99092
rect 177772 96684 177828 96740
rect 177212 94892 177268 94948
rect 176988 83132 177044 83188
rect 175644 80556 175700 80612
rect 176316 80220 176372 80276
rect 177212 80556 177268 80612
rect 177660 80556 177716 80612
rect 179676 99484 179732 99540
rect 179676 96572 179732 96628
rect 180572 98476 180628 98532
rect 179676 91532 179732 91588
rect 179004 79772 179060 79828
rect 180348 83244 180404 83300
rect 180572 80556 180628 80612
rect 181692 93436 181748 93492
rect 182364 91644 182420 91700
rect 188412 98588 188468 98644
rect 185724 98364 185780 98420
rect 183708 95116 183764 95172
rect 184380 91756 184436 91812
rect 185052 80556 185108 80612
rect 187292 91868 187348 91924
rect 186396 89852 186452 89908
rect 187068 81452 187124 81508
rect 187292 80556 187348 80612
rect 187740 86492 187796 86548
rect 189084 96796 189140 96852
rect 189532 80556 189588 80612
rect 190428 80556 190484 80612
rect 199836 101500 199892 101556
rect 192444 100268 192500 100324
rect 191772 86604 191828 86660
rect 195804 96908 195860 96964
rect 195692 91980 195748 92036
rect 192668 89964 192724 90020
rect 195132 88172 195188 88228
rect 193788 86716 193844 86772
rect 192668 80556 192724 80612
rect 193116 80556 193172 80612
rect 194460 78204 194516 78260
rect 195692 80556 195748 80612
rect 198156 90188 198212 90244
rect 197820 81564 197876 81620
rect 197148 79996 197204 80052
rect 196476 78988 196532 79044
rect 198156 78988 198212 79044
rect 198492 90076 198548 90132
rect 199164 80332 199220 80388
rect 218652 101388 218708 101444
rect 203868 100380 203924 100436
rect 200508 98700 200564 98756
rect 201180 92092 201236 92148
rect 203196 90300 203252 90356
rect 201852 83356 201908 83412
rect 202524 80556 202580 80612
rect 205884 98812 205940 98868
rect 205212 90412 205268 90468
rect 204876 80556 204932 80612
rect 209916 97020 209972 97076
rect 209244 93660 209300 93716
rect 207900 93548 207956 93604
rect 207228 90524 207284 90580
rect 206556 80556 206612 80612
rect 208572 80444 208628 80500
rect 211260 95228 211316 95284
rect 210588 88284 210644 88340
rect 216748 88396 216804 88452
rect 212604 86828 212660 86884
rect 211932 84812 211988 84868
rect 215964 85036 216020 85092
rect 215292 84924 215348 84980
rect 213276 81676 213332 81732
rect 213948 80556 214004 80612
rect 214844 80556 214900 80612
rect 216636 83580 216692 83636
rect 218428 83692 218484 83748
rect 216748 80444 216804 80500
rect 217980 83468 218036 83524
rect 217308 80108 217364 80164
rect 218428 78988 218484 79044
rect 266252 100828 266308 100884
rect 246204 100604 246260 100660
rect 234332 100492 234388 100548
rect 221340 96684 221396 96740
rect 219996 95004 220052 95060
rect 219324 79884 219380 79940
rect 220668 80668 220724 80724
rect 223356 96572 223412 96628
rect 222684 85148 222740 85204
rect 222012 78988 222068 79044
rect 224700 87052 224756 87108
rect 224028 80108 224084 80164
rect 225148 85148 225204 85204
rect 230188 83804 230244 83860
rect 228620 83692 228676 83748
rect 226604 80556 226660 80612
rect 226044 80444 226100 80500
rect 225148 80220 225204 80276
rect 225372 80220 225428 80276
rect 228396 80556 228452 80612
rect 227388 78988 227444 79044
rect 229964 80556 230020 80612
rect 228620 80220 228676 80276
rect 228732 80444 228788 80500
rect 230188 80108 230244 80164
rect 232092 80556 232148 80612
rect 230076 79660 230132 79716
rect 231420 79548 231476 79604
rect 230748 79324 230804 79380
rect 233436 80556 233492 80612
rect 232764 79436 232820 79492
rect 234108 80556 234164 80612
rect 244860 99932 244916 99988
rect 235452 98252 235508 98308
rect 234332 79772 234388 79828
rect 234780 79772 234836 79828
rect 242844 96572 242900 96628
rect 238588 90636 238644 90692
rect 237692 86940 237748 86996
rect 236124 80556 236180 80612
rect 237468 80220 237524 80276
rect 236796 80108 236852 80164
rect 237692 79996 237748 80052
rect 238476 80556 238532 80612
rect 241836 80556 241892 80612
rect 238588 80332 238644 80388
rect 240828 80332 240884 80388
rect 239484 79996 239540 80052
rect 238812 79772 238868 79828
rect 240156 79884 240212 79940
rect 242172 80556 242228 80612
rect 243516 93212 243572 93268
rect 244188 80556 244244 80612
rect 245532 96684 245588 96740
rect 248892 97468 248948 97524
rect 248220 95788 248276 95844
rect 247548 94108 247604 94164
rect 246876 80556 246932 80612
rect 258300 95900 258356 95956
rect 256284 94556 256340 94612
rect 250236 92540 250292 92596
rect 249564 80556 249620 80612
rect 252252 92428 252308 92484
rect 251916 80556 251972 80612
rect 250908 77308 250964 77364
rect 255612 90748 255668 90804
rect 253484 80556 253540 80612
rect 252924 79660 252980 79716
rect 254268 80556 254324 80612
rect 254492 80444 254548 80500
rect 257628 94220 257684 94276
rect 256956 79660 257012 79716
rect 260988 94332 261044 94388
rect 260316 92652 260372 92708
rect 259644 80556 259700 80612
rect 258972 79100 259028 79156
rect 166348 60284 166404 60340
rect 166012 57260 166068 57316
rect 153692 31948 153748 32004
rect 163772 42700 163828 42756
rect 163772 19964 163828 20020
rect 163996 40908 164052 40964
rect 164556 39116 164612 39172
rect 164444 37324 164500 37380
rect 164220 35532 164276 35588
rect 164220 20076 164276 20132
rect 163996 19628 164052 19684
rect 164556 18508 164612 18564
rect 265244 18508 265300 18564
rect 164444 18284 164500 18340
rect 150332 17612 150388 17668
rect 4172 16716 4228 16772
rect 216860 16716 216916 16772
rect 217532 16716 217588 16772
rect 219100 16716 219156 16772
rect 221116 16716 221172 16772
rect 222460 16716 222516 16772
rect 222908 16716 222964 16772
rect 225820 16716 225876 16772
rect 226268 16716 226324 16772
rect 230748 16716 230804 16772
rect 231196 16716 231252 16772
rect 236572 16716 236628 16772
rect 239260 16716 239316 16772
rect 239932 16716 239988 16772
rect 240380 16716 240436 16772
rect 240604 16716 240660 16772
rect 243740 16716 243796 16772
rect 245084 16716 245140 16772
rect 223132 16604 223188 16660
rect 238588 16604 238644 16660
rect 245308 16268 245364 16324
rect 249564 16268 249620 16324
rect 216636 16156 216692 16212
rect 248556 16156 248612 16212
rect 114268 16044 114324 16100
rect 106540 14588 106596 14644
rect 69692 14476 69748 14532
rect 42812 14252 42868 14308
rect 37772 12572 37828 12628
rect 32508 10892 32564 10948
rect 24892 9212 24948 9268
rect 21084 7532 21140 7588
rect 17276 4172 17332 4228
rect 11564 3388 11620 3444
rect 13356 3388 13412 3444
rect 15372 2492 15428 2548
rect 19180 4172 19236 4228
rect 22988 4284 23044 4340
rect 30604 5852 30660 5908
rect 28700 4284 28756 4340
rect 26796 3388 26852 3444
rect 34412 6188 34468 6244
rect 36316 4060 36372 4116
rect 37772 4060 37828 4116
rect 42028 4060 42084 4116
rect 40124 3724 40180 3780
rect 53228 13468 53284 13524
rect 49644 11228 49700 11284
rect 47740 11004 47796 11060
rect 42812 4060 42868 4116
rect 43932 4396 43988 4452
rect 51548 6748 51604 6804
rect 38332 28 38388 84
rect 45948 140 46004 196
rect 54572 12684 54628 12740
rect 54572 6748 54628 6804
rect 61068 9324 61124 9380
rect 55356 3836 55412 3892
rect 57260 2604 57316 2660
rect 62972 7644 63028 7700
rect 66780 5964 66836 6020
rect 68684 4060 68740 4116
rect 104636 13692 104692 13748
rect 87500 13580 87556 13636
rect 81452 12908 81508 12964
rect 74172 12796 74228 12852
rect 72492 7532 72548 7588
rect 69692 4060 69748 4116
rect 70476 6076 70532 6132
rect 59276 252 59332 308
rect 65436 364 65492 420
rect 78204 11116 78260 11172
rect 76412 476 76468 532
rect 85820 8428 85876 8484
rect 83916 7756 83972 7812
rect 81452 7644 81508 7700
rect 82012 7644 82068 7700
rect 80108 4508 80164 4564
rect 92316 13020 92372 13076
rect 89628 9436 89684 9492
rect 92316 8428 92372 8484
rect 97244 9548 97300 9604
rect 91532 7868 91588 7924
rect 93436 4620 93492 4676
rect 95340 2716 95396 2772
rect 99036 2828 99092 2884
rect 102956 700 103012 756
rect 101052 588 101108 644
rect 112476 9660 112532 9716
rect 108668 7980 108724 8036
rect 110572 2940 110628 2996
rect 137004 15932 137060 15988
rect 117964 15148 118020 15204
rect 116732 13132 116788 13188
rect 116284 6300 116340 6356
rect 116732 6188 116788 6244
rect 133196 14700 133252 14756
rect 129612 11340 129668 11396
rect 127596 6524 127652 6580
rect 121996 6412 122052 6468
rect 120092 6188 120148 6244
rect 123900 3052 123956 3108
rect 125804 812 125860 868
rect 131516 8204 131572 8260
rect 135324 11452 135380 11508
rect 148428 15820 148484 15876
rect 142828 15260 142884 15316
rect 141036 11228 141092 11284
rect 139132 3164 139188 3220
rect 144620 14812 144676 14868
rect 146748 8092 146804 8148
rect 167468 14364 167524 14420
rect 154140 13244 154196 13300
rect 152460 9772 152516 9828
rect 150556 3276 150612 3332
rect 165564 12012 165620 12068
rect 158172 11564 158228 11620
rect 156156 4732 156212 4788
rect 160076 9884 160132 9940
rect 163884 6636 163940 6692
rect 161980 2380 162036 2436
rect 179116 12348 179172 12404
rect 175308 11676 175364 11732
rect 171500 10780 171556 10836
rect 169596 9996 169652 10052
rect 173404 8316 173460 8372
rect 177212 9100 177268 9156
rect 179116 8204 179172 8260
rect 184716 8204 184772 8260
rect 179116 7420 179172 7476
rect 181020 5740 181076 5796
rect 182924 4844 182980 4900
rect 185836 12962 185892 12964
rect 185836 12910 185838 12962
rect 185838 12910 185890 12962
rect 185890 12910 185892 12962
rect 185836 12908 185892 12910
rect 185948 12236 186004 12292
rect 186508 12962 186564 12964
rect 186508 12910 186510 12962
rect 186510 12910 186562 12962
rect 186562 12910 186564 12962
rect 186508 12908 186564 12910
rect 186396 12460 186452 12516
rect 186172 12236 186228 12292
rect 186844 13356 186900 13412
rect 187068 13356 187124 13412
rect 187516 12236 187572 12292
rect 187292 9212 187348 9268
rect 186620 4172 186676 4228
rect 186732 4956 186788 5012
rect 185724 2492 185780 2548
rect 186060 1036 186116 1092
rect 186060 700 186116 756
rect 188412 13132 188468 13188
rect 188636 12572 188692 12628
rect 188188 10892 188244 10948
rect 187964 5852 188020 5908
rect 188636 9212 188692 9268
rect 187740 4284 187796 4340
rect 189308 14252 189364 14308
rect 189084 12236 189140 12292
rect 189308 12124 189364 12180
rect 190204 13132 190260 13188
rect 190652 13356 190708 13412
rect 190428 12684 190484 12740
rect 190652 12684 190708 12740
rect 189980 11004 190036 11060
rect 189532 4396 189588 4452
rect 190540 10892 190596 10948
rect 189308 2604 189364 2660
rect 190876 12236 190932 12292
rect 191100 12124 191156 12180
rect 190652 10780 190708 10836
rect 189644 140 189700 196
rect 188860 28 188916 84
rect 191436 12236 191492 12292
rect 191772 12908 191828 12964
rect 191548 9324 191604 9380
rect 191436 6076 191492 6132
rect 192444 14476 192500 14532
rect 192556 12572 192612 12628
rect 192332 12460 192388 12516
rect 192332 7756 192388 7812
rect 192444 12124 192500 12180
rect 192220 5964 192276 6020
rect 192444 4508 192500 4564
rect 192668 12236 192724 12292
rect 193116 13132 193172 13188
rect 192892 7532 192948 7588
rect 191996 476 192052 532
rect 193452 12236 193508 12292
rect 193788 12124 193844 12180
rect 193564 11116 193620 11172
rect 194012 7644 194068 7700
rect 194124 12796 194180 12852
rect 193452 2716 193508 2772
rect 193340 700 193396 756
rect 191324 252 191380 308
rect 194684 13356 194740 13412
rect 194460 13020 194516 13076
rect 194236 12460 194292 12516
rect 194908 9436 194964 9492
rect 195132 7868 195188 7924
rect 195580 12236 195636 12292
rect 195804 9548 195860 9604
rect 195356 4620 195412 4676
rect 196140 11004 196196 11060
rect 196028 2828 196084 2884
rect 196364 1148 196420 1204
rect 196924 14588 196980 14644
rect 196700 13692 196756 13748
rect 197148 7980 197204 8036
rect 197372 2940 197428 2996
rect 197484 12236 197540 12292
rect 196476 1036 196532 1092
rect 197820 16044 197876 16100
rect 197596 9660 197652 9716
rect 198156 15148 198212 15204
rect 198044 6300 198100 6356
rect 198716 6412 198772 6468
rect 198492 6188 198548 6244
rect 197484 812 197540 868
rect 198156 4172 198212 4228
rect 199164 12236 199220 12292
rect 199500 11900 199556 11956
rect 200060 14700 200116 14756
rect 199836 12348 199892 12404
rect 200508 16044 200564 16100
rect 200284 11452 200340 11508
rect 199612 11340 199668 11396
rect 200396 9996 200452 10052
rect 199500 9772 199556 9828
rect 200060 9884 200116 9940
rect 199388 6524 199444 6580
rect 198940 3052 198996 3108
rect 200396 9660 200452 9716
rect 201180 15260 201236 15316
rect 201404 14812 201460 14868
rect 200956 11228 201012 11284
rect 201292 11676 201348 11732
rect 201852 15820 201908 15876
rect 201628 8092 201684 8148
rect 201964 9996 202020 10052
rect 201292 4732 201348 4788
rect 200732 3164 200788 3220
rect 202524 13244 202580 13300
rect 202300 11900 202356 11956
rect 202748 11676 202804 11732
rect 202972 11340 203028 11396
rect 203196 9772 203252 9828
rect 202076 3276 202132 3332
rect 204092 14364 204148 14420
rect 203868 12012 203924 12068
rect 204092 12236 204148 12292
rect 203644 6636 203700 6692
rect 203868 8428 203924 8484
rect 203420 2380 203476 2436
rect 204540 12684 204596 12740
rect 204316 9772 204372 9828
rect 204988 11452 205044 11508
rect 205436 12236 205492 12292
rect 205548 13244 205604 13300
rect 205212 9100 205268 9156
rect 204764 8316 204820 8372
rect 204092 7420 204148 7476
rect 205660 5740 205716 5796
rect 206108 8204 206164 8260
rect 207228 12796 207284 12852
rect 207004 12572 207060 12628
rect 207452 11004 207508 11060
rect 207564 13356 207620 13412
rect 206780 10892 206836 10948
rect 206556 9212 206612 9268
rect 206332 4956 206388 5012
rect 205884 4844 205940 4900
rect 208124 9996 208180 10052
rect 207900 9884 207956 9940
rect 208796 13356 208852 13412
rect 208572 13244 208628 13300
rect 208348 8428 208404 8484
rect 207676 4172 207732 4228
rect 209468 13356 209524 13412
rect 209692 13356 209748 13412
rect 209916 13356 209972 13412
rect 210140 13356 210196 13412
rect 209244 4396 209300 4452
rect 210588 6748 210644 6804
rect 211036 11564 211092 11620
rect 211260 9324 211316 9380
rect 211484 6412 211540 6468
rect 211932 12796 211988 12852
rect 212156 12684 212212 12740
rect 212380 11452 212436 11508
rect 212604 9212 212660 9268
rect 211708 6076 211764 6132
rect 210812 4284 210868 4340
rect 211260 4396 211316 4452
rect 210364 4172 210420 4228
rect 212828 4396 212884 4452
rect 213500 11676 213556 11732
rect 213276 8092 213332 8148
rect 213948 8204 214004 8260
rect 214172 7756 214228 7812
rect 213724 7532 213780 7588
rect 214620 15484 214676 15540
rect 214396 6300 214452 6356
rect 215292 15596 215348 15652
rect 215068 12012 215124 12068
rect 215964 15820 216020 15876
rect 215740 14252 215796 14308
rect 216412 13356 216468 13412
rect 217308 16044 217364 16100
rect 217084 13244 217140 13300
rect 216188 9660 216244 9716
rect 216748 11676 216804 11732
rect 215516 7644 215572 7700
rect 214844 5852 214900 5908
rect 215068 6748 215124 6804
rect 213052 4060 213108 4116
rect 213164 4172 213220 4228
rect 217756 11340 217812 11396
rect 218876 14476 218932 14532
rect 218652 13356 218708 13412
rect 218428 10780 218484 10836
rect 218876 11564 218932 11620
rect 218204 10108 218260 10164
rect 217980 6188 218036 6244
rect 216748 4620 216804 4676
rect 216972 4284 217028 4340
rect 219772 16044 219828 16100
rect 219996 14924 220052 14980
rect 220444 13132 220500 13188
rect 220668 12572 220724 12628
rect 221340 14924 221396 14980
rect 220892 12460 220948 12516
rect 221564 10892 221620 10948
rect 220220 10444 220276 10500
rect 219548 5964 219604 6020
rect 220780 9324 220836 9380
rect 219324 2604 219380 2660
rect 222236 14924 222292 14980
rect 222012 12908 222068 12964
rect 223356 12236 223412 12292
rect 222684 8316 222740 8372
rect 221788 3276 221844 3332
rect 222684 6412 222740 6468
rect 224028 12348 224084 12404
rect 223804 11116 223860 11172
rect 224476 13356 224532 13412
rect 224700 12236 224756 12292
rect 224252 9548 224308 9604
rect 224924 9436 224980 9492
rect 223580 2268 223636 2324
rect 224588 6076 224644 6132
rect 225372 12348 225428 12404
rect 226044 16044 226100 16100
rect 226492 15708 226548 15764
rect 225596 9324 225652 9380
rect 226492 12796 226548 12852
rect 225148 3164 225204 3220
rect 226828 15372 226884 15428
rect 226828 13132 226884 13188
rect 226716 12236 226772 12292
rect 227164 15148 227220 15204
rect 227388 12796 227444 12852
rect 226940 7980 226996 8036
rect 228060 12236 228116 12292
rect 228508 14364 228564 14420
rect 228284 12124 228340 12180
rect 228508 12684 228564 12740
rect 227836 11004 227892 11060
rect 227612 6076 227668 6132
rect 226828 5852 226884 5908
rect 226828 4508 226884 4564
rect 228620 7756 228676 7812
rect 229404 12236 229460 12292
rect 229180 11676 229236 11732
rect 228956 11228 229012 11284
rect 229628 7868 229684 7924
rect 228732 6636 228788 6692
rect 228620 3948 228676 4004
rect 230188 13580 230244 13636
rect 230188 13244 230244 13300
rect 230076 9996 230132 10052
rect 230188 11452 230244 11508
rect 230412 15260 230468 15316
rect 230412 13356 230468 13412
rect 230188 6300 230244 6356
rect 230188 4060 230244 4116
rect 229852 2380 229908 2436
rect 230188 3276 230244 3332
rect 230188 1036 230244 1092
rect 230412 7756 230468 7812
rect 231420 12684 231476 12740
rect 231644 12236 231700 12292
rect 232092 12684 232148 12740
rect 232204 9212 232260 9268
rect 230972 5852 231028 5908
rect 230524 1260 230580 1316
rect 232092 588 232148 644
rect 232540 12348 232596 12404
rect 232316 3052 232372 3108
rect 232988 12236 233044 12292
rect 233436 13804 233492 13860
rect 233436 12012 233492 12068
rect 233324 11676 233380 11732
rect 233436 7644 233492 7700
rect 233436 4396 233492 4452
rect 233212 2044 233268 2100
rect 232764 1596 232820 1652
rect 233884 14588 233940 14644
rect 233660 1484 233716 1540
rect 234108 4284 234164 4340
rect 234332 7644 234388 7700
rect 234220 2828 234276 2884
rect 234780 13132 234836 13188
rect 234892 12684 234948 12740
rect 234892 9212 234948 9268
rect 235228 13244 235284 13300
rect 235116 12348 235172 12404
rect 235116 9100 235172 9156
rect 235116 7532 235172 7588
rect 235116 4844 235172 4900
rect 235004 3276 235060 3332
rect 234556 1372 234612 1428
rect 235676 7532 235732 7588
rect 236124 13356 236180 13412
rect 235900 2716 235956 2772
rect 236012 4172 236068 4228
rect 235452 1148 235508 1204
rect 236796 12908 236852 12964
rect 237244 11788 237300 11844
rect 237020 11564 237076 11620
rect 236796 8204 236852 8260
rect 237468 6412 237524 6468
rect 236796 4172 236852 4228
rect 237916 12348 237972 12404
rect 237804 12236 237860 12292
rect 238364 12236 238420 12292
rect 238140 12012 238196 12068
rect 239036 12684 239092 12740
rect 238812 11788 238868 11844
rect 238476 9660 238532 9716
rect 237804 6524 237860 6580
rect 237916 8092 237972 8148
rect 237692 588 237748 644
rect 236348 476 236404 532
rect 240268 13692 240324 13748
rect 240268 12460 240324 12516
rect 240492 12908 240548 12964
rect 240828 12908 240884 12964
rect 240492 12460 240548 12516
rect 240156 12236 240212 12292
rect 239708 9884 239764 9940
rect 241500 13356 241556 13412
rect 241276 12236 241332 12292
rect 241724 9660 241780 9716
rect 241052 8204 241108 8260
rect 239484 4956 239540 5012
rect 238476 4732 238532 4788
rect 241724 4844 241780 4900
rect 239820 4620 239876 4676
rect 242396 12796 242452 12852
rect 242172 12348 242228 12404
rect 242620 11788 242676 11844
rect 241948 4844 242004 4900
rect 243068 14924 243124 14980
rect 243292 13356 243348 13412
rect 243292 12124 243348 12180
rect 244188 12796 244244 12852
rect 244412 12348 244468 12404
rect 244524 14588 244580 14644
rect 244412 12124 244468 12180
rect 244412 11900 244468 11956
rect 244860 14924 244916 14980
rect 244636 12124 244692 12180
rect 245532 12124 245588 12180
rect 245980 13356 246036 13412
rect 247772 15372 247828 15428
rect 245756 8092 245812 8148
rect 244524 6300 244580 6356
rect 243964 4732 244020 4788
rect 242844 4284 242900 4340
rect 243628 4172 243684 4228
rect 247436 4060 247492 4116
rect 245532 3948 245588 4004
rect 248556 11900 248612 11956
rect 249228 15484 249284 15540
rect 249452 13244 249508 13300
rect 249452 12460 249508 12516
rect 249340 11452 249396 11508
rect 249452 10108 249508 10164
rect 249452 9100 249508 9156
rect 249340 8876 249396 8932
rect 248556 3612 248612 3668
rect 248556 3164 248612 3220
rect 247772 924 247828 980
rect 248668 1260 248724 1316
rect 248668 364 248724 420
rect 260764 15820 260820 15876
rect 255052 15596 255108 15652
rect 253708 15372 253764 15428
rect 253708 15036 253764 15092
rect 253148 13804 253204 13860
rect 251916 11340 251972 11396
rect 249564 1148 249620 1204
rect 251244 4508 251300 4564
rect 251916 4060 251972 4116
rect 258860 14252 258916 14308
rect 257068 8876 257124 8932
rect 257068 4620 257124 4676
rect 257068 4396 257124 4452
rect 264572 13468 264628 13524
rect 264460 10108 264516 10164
rect 262668 4284 262724 4340
rect 264460 2940 264516 2996
rect 265468 15260 265524 15316
rect 265468 13356 265524 13412
rect 265692 15036 265748 15092
rect 265468 11116 265524 11172
rect 268156 96460 268212 96516
rect 266252 13132 266308 13188
rect 266364 94444 266420 94500
rect 265692 11116 265748 11172
rect 266700 90860 266756 90916
rect 266588 81004 266644 81060
rect 266364 9884 266420 9940
rect 266476 16044 266532 16100
rect 265468 8204 265524 8260
rect 265804 7980 265860 8036
rect 265468 5068 265524 5124
rect 265468 4732 265524 4788
rect 265692 4620 265748 4676
rect 265244 3052 265300 3108
rect 265580 3388 265636 3444
rect 265468 2492 265524 2548
rect 265580 2380 265636 2436
rect 265804 3052 265860 3108
rect 265692 2156 265748 2212
rect 265468 924 265524 980
rect 266924 85260 266980 85316
rect 266700 8316 266756 8372
rect 266812 76300 266868 76356
rect 269612 96012 269668 96068
rect 268156 83804 268212 83860
rect 268828 85708 268884 85764
rect 267932 83244 267988 83300
rect 267932 83020 267988 83076
rect 268268 80780 268324 80836
rect 268156 78876 268212 78932
rect 266924 14924 266980 14980
rect 267036 78316 267092 78372
rect 267932 78092 267988 78148
rect 267036 11564 267092 11620
rect 267820 13356 267876 13412
rect 266812 6412 266868 6468
rect 267820 4508 267876 4564
rect 266588 2828 266644 2884
rect 268044 77196 268100 77252
rect 268044 4844 268100 4900
rect 268604 78540 268660 78596
rect 268268 13244 268324 13300
rect 268380 17052 268436 17108
rect 268156 2716 268212 2772
rect 267932 1484 267988 1540
rect 268828 18396 268884 18452
rect 268940 82348 268996 82404
rect 268940 18284 268996 18340
rect 269500 17276 269556 17332
rect 268604 16828 268660 16884
rect 269388 17164 269444 17220
rect 269276 15932 269332 15988
rect 269164 15372 269220 15428
rect 268716 14588 268772 14644
rect 268492 13356 268548 13412
rect 268716 13244 268772 13300
rect 268716 12908 268772 12964
rect 268716 11676 268772 11732
rect 268940 10892 268996 10948
rect 269164 9100 269220 9156
rect 269388 9884 269444 9940
rect 269276 8092 269332 8148
rect 273084 305004 273140 305060
rect 273084 218428 273140 218484
rect 273084 96460 273140 96516
rect 273980 305228 274036 305284
rect 273532 94892 273588 94948
rect 273868 305116 273924 305172
rect 272972 93436 273028 93492
rect 273756 93436 273812 93492
rect 271292 91084 271348 91140
rect 269724 86044 269780 86100
rect 270620 84476 270676 84532
rect 269836 84252 269892 84308
rect 270284 84140 270340 84196
rect 271180 83244 271236 83300
rect 273868 93324 273924 93380
rect 273756 87052 273812 87108
rect 274652 230972 274708 231028
rect 274652 218428 274708 218484
rect 275324 101612 275380 101668
rect 275772 100492 275828 100548
rect 274876 98476 274932 98532
rect 276220 91532 276276 91588
rect 276332 90972 276388 91028
rect 276332 85260 276388 85316
rect 274428 83132 274484 83188
rect 274652 83804 274708 83860
rect 271292 78876 271348 78932
rect 271180 78540 271236 78596
rect 277116 101724 277172 101780
rect 277228 305452 277284 305508
rect 277564 305340 277620 305396
rect 277228 100156 277284 100212
rect 278348 304892 278404 304948
rect 278012 91644 278068 91700
rect 278124 304332 278180 304388
rect 276668 83132 276724 83188
rect 278460 101836 278516 101892
rect 278348 96796 278404 96852
rect 279020 245196 279076 245252
rect 279020 236796 279076 236852
rect 278908 95116 278964 95172
rect 280252 98364 280308 98420
rect 279804 91868 279860 91924
rect 279356 91756 279412 91812
rect 281148 304332 281204 304388
rect 281372 305116 281428 305172
rect 281372 101948 281428 102004
rect 280700 89852 280756 89908
rect 282604 305228 282660 305284
rect 283052 305340 283108 305396
rect 282492 304892 282548 304948
rect 282044 98588 282100 98644
rect 283052 96908 283108 96964
rect 283836 305116 283892 305172
rect 283388 89964 283444 90020
rect 284732 305452 284788 305508
rect 284732 305228 284788 305284
rect 284956 305116 285012 305172
rect 285628 305228 285684 305284
rect 285740 305452 285796 305508
rect 285292 304892 285348 304948
rect 285628 251916 285684 251972
rect 285628 245196 285684 245252
rect 286300 305228 286356 305284
rect 286972 305340 287028 305396
rect 286524 305116 286580 305172
rect 286412 250236 286468 250292
rect 286412 230972 286468 231028
rect 285740 100268 285796 100324
rect 285292 93660 285348 93716
rect 286412 96012 286468 96068
rect 285180 91980 285236 92036
rect 287420 90188 287476 90244
rect 286412 89852 286468 89908
rect 284956 88172 285012 88228
rect 284732 86716 284788 86772
rect 287308 87388 287364 87444
rect 284284 86604 284340 86660
rect 281596 86492 281652 86548
rect 282156 84364 282212 84420
rect 287868 86940 287924 86996
rect 287308 83916 287364 83972
rect 282156 83244 282212 83300
rect 278124 81452 278180 81508
rect 282156 82460 282212 82516
rect 289660 101500 289716 101556
rect 290108 98700 290164 98756
rect 290556 92092 290612 92148
rect 289212 90636 289268 90692
rect 288764 90076 288820 90132
rect 291452 305228 291508 305284
rect 291452 268716 291508 268772
rect 291676 268604 291732 268660
rect 291676 251916 291732 251972
rect 291452 250236 291508 250292
rect 292796 305228 292852 305284
rect 292348 100380 292404 100436
rect 294140 305228 294196 305284
rect 293692 98812 293748 98868
rect 295036 93548 295092 93604
rect 294588 90524 294644 90580
rect 293244 90412 293300 90468
rect 291900 90300 291956 90356
rect 295932 304892 295988 304948
rect 296380 97020 296436 97076
rect 295484 88396 295540 88452
rect 297388 273868 297444 273924
rect 297388 268604 297444 268660
rect 297276 95228 297332 95284
rect 296828 88284 296884 88340
rect 295596 88060 295652 88116
rect 291004 83356 291060 83412
rect 292236 86156 292292 86212
rect 288316 81564 288372 81620
rect 282156 79548 282212 79604
rect 287196 81452 287252 81508
rect 274652 78428 274708 78484
rect 298172 86828 298228 86884
rect 298284 305116 298340 305172
rect 297724 84812 297780 84868
rect 298284 83580 298340 83636
rect 295596 81788 295652 81844
rect 299068 305340 299124 305396
rect 299516 305228 299572 305284
rect 298956 91084 299012 91140
rect 299068 87388 299124 87444
rect 299068 85260 299124 85316
rect 299180 85708 299236 85764
rect 298956 84812 299012 84868
rect 300860 305116 300916 305172
rect 300748 271292 300804 271348
rect 300748 268716 300804 268772
rect 301532 291452 301588 291508
rect 301532 273868 301588 273924
rect 301308 85148 301364 85204
rect 300412 85036 300468 85092
rect 299964 84924 300020 84980
rect 302652 304892 302708 304948
rect 303996 303996 304052 304052
rect 304892 306684 304948 306740
rect 305340 306572 305396 306628
rect 304444 303660 304500 303716
rect 303548 303436 303604 303492
rect 305788 303212 305844 303268
rect 303100 301644 303156 301700
rect 306684 305228 306740 305284
rect 308476 305676 308532 305732
rect 308028 305452 308084 305508
rect 307580 305340 307636 305396
rect 307132 305116 307188 305172
rect 308924 304668 308980 304724
rect 306236 301532 306292 301588
rect 309820 301868 309876 301924
rect 309372 301308 309428 301364
rect 310716 306908 310772 306964
rect 311164 306796 311220 306852
rect 311612 303772 311668 303828
rect 311836 304220 311892 304276
rect 310268 299852 310324 299908
rect 311164 280588 311220 280644
rect 311164 271292 311220 271348
rect 302204 101388 302260 101444
rect 309148 94892 309204 94948
rect 309148 93436 309204 93492
rect 312508 303884 312564 303940
rect 312060 303548 312116 303604
rect 313404 305564 313460 305620
rect 312956 301756 313012 301812
rect 314300 304780 314356 304836
rect 315196 304556 315252 304612
rect 315084 304108 315140 304164
rect 314748 302204 314804 302260
rect 314972 302652 315028 302708
rect 313852 300412 313908 300468
rect 312508 296604 312564 296660
rect 312508 291452 312564 291508
rect 311836 89964 311892 90020
rect 316092 307356 316148 307412
rect 316540 306460 316596 306516
rect 315644 303324 315700 303380
rect 315084 91532 315140 91588
rect 315196 300972 315252 301028
rect 316988 300076 317044 300132
rect 317884 307132 317940 307188
rect 318332 303996 318388 304052
rect 318444 305788 318500 305844
rect 317436 298060 317492 298116
rect 318332 302540 318388 302596
rect 316652 296716 316708 296772
rect 316652 280588 316708 280644
rect 315196 87052 315252 87108
rect 315644 87948 315700 88004
rect 314972 86492 315028 86548
rect 318444 91644 318500 91700
rect 318556 302428 318612 302484
rect 319676 305228 319732 305284
rect 320124 305228 320180 305284
rect 319228 303324 319284 303380
rect 321020 302428 321076 302484
rect 322364 307244 322420 307300
rect 321916 307020 321972 307076
rect 321468 302092 321524 302148
rect 320572 301980 320628 302036
rect 318780 299964 318836 300020
rect 318892 300860 318948 300916
rect 318668 297948 318724 298004
rect 318668 90300 318724 90356
rect 318556 86940 318612 86996
rect 322812 300300 322868 300356
rect 323148 304892 323204 304948
rect 323260 303100 323316 303156
rect 323484 305228 323540 305284
rect 324156 305676 324212 305732
rect 324604 305676 324660 305732
rect 325052 304892 325108 304948
rect 325388 306684 325444 306740
rect 323708 304332 323764 304388
rect 324940 303660 324996 303716
rect 324044 303436 324100 303492
rect 323484 301420 323540 301476
rect 323596 301644 323652 301700
rect 324492 302764 324548 302820
rect 325500 304668 325556 304724
rect 325948 304220 326004 304276
rect 326284 306572 326340 306628
rect 325836 301308 325892 301364
rect 326396 304556 326452 304612
rect 326508 304444 326564 304500
rect 326508 300748 326564 300804
rect 326732 303212 326788 303268
rect 327740 306572 327796 306628
rect 327292 305676 327348 305732
rect 327180 305452 327236 305508
rect 327180 303660 327236 303716
rect 327740 304108 327796 304164
rect 328188 303436 328244 303492
rect 328524 303660 328580 303716
rect 326844 301644 326900 301700
rect 328076 302540 328132 302596
rect 327180 301532 327236 301588
rect 329084 305452 329140 305508
rect 328636 303212 328692 303268
rect 328972 300748 329028 300804
rect 329420 300748 329476 300804
rect 329980 306684 330036 306740
rect 330428 305676 330484 305732
rect 330876 304332 330932 304388
rect 331212 306908 331268 306964
rect 330316 301868 330372 301924
rect 329532 300188 329588 300244
rect 329868 300748 329924 300804
rect 330764 299852 330820 299908
rect 331324 305116 331380 305172
rect 331660 306796 331716 306852
rect 331772 305564 331828 305620
rect 332108 303772 332164 303828
rect 319116 298284 319172 298340
rect 332668 306796 332724 306852
rect 333004 303884 333060 303940
rect 332556 303548 332612 303604
rect 334012 303884 334068 303940
rect 333564 303548 333620 303604
rect 334908 306908 334964 306964
rect 335356 305676 335412 305732
rect 334460 302988 334516 303044
rect 334796 305004 334852 305060
rect 333116 299852 333172 299908
rect 333452 301756 333508 301812
rect 334348 300748 334404 300804
rect 333900 300412 333956 300468
rect 335020 305004 335076 305060
rect 335020 304220 335076 304276
rect 335692 303660 335748 303716
rect 335244 302204 335300 302260
rect 336252 305340 336308 305396
rect 336588 307356 336644 307412
rect 335804 301532 335860 301588
rect 336140 300860 336196 300916
rect 336700 304780 336756 304836
rect 337036 306460 337092 306516
rect 337148 301868 337204 301924
rect 338044 307356 338100 307412
rect 337596 301756 337652 301812
rect 338380 307132 338436 307188
rect 337484 300076 337540 300132
rect 338492 303660 338548 303716
rect 338828 303996 338884 304052
rect 339388 307132 339444 307188
rect 338940 303772 338996 303828
rect 339724 305228 339780 305284
rect 339276 299964 339332 300020
rect 339836 303884 339892 303940
rect 340172 303324 340228 303380
rect 340284 299964 340340 300020
rect 340620 301420 340676 301476
rect 322028 298284 322084 298340
rect 332332 298284 332388 298340
rect 337932 298284 337988 298340
rect 341180 305116 341236 305172
rect 342076 305116 342132 305172
rect 342412 307020 342468 307076
rect 341628 304444 341684 304500
rect 341516 302316 341572 302372
rect 341068 301980 341124 302036
rect 341964 302092 342020 302148
rect 342524 305676 342580 305732
rect 342860 307244 342916 307300
rect 342524 304668 342580 304724
rect 342524 300860 342580 300916
rect 343868 307244 343924 307300
rect 343420 307020 343476 307076
rect 342972 305676 343028 305732
rect 343756 303100 343812 303156
rect 343308 300300 343364 300356
rect 344204 302876 344260 302932
rect 344316 301980 344372 302036
rect 344652 304108 344708 304164
rect 344764 303996 344820 304052
rect 345660 306348 345716 306404
rect 345212 303324 345268 303380
rect 345996 304892 346052 304948
rect 345548 300860 345604 300916
rect 345100 300748 345156 300804
rect 346108 300076 346164 300132
rect 346444 305228 346500 305284
rect 347004 305564 347060 305620
rect 346556 304892 346612 304948
rect 347340 301644 347396 301700
rect 346892 301084 346948 301140
rect 347900 305228 347956 305284
rect 348236 306572 348292 306628
rect 347452 301420 347508 301476
rect 347788 305116 347844 305172
rect 347788 301196 347844 301252
rect 347788 300972 347844 301028
rect 348796 306572 348852 306628
rect 348348 301084 348404 301140
rect 348684 303436 348740 303492
rect 349132 303212 349188 303268
rect 349356 304332 349412 304388
rect 350140 306460 350196 306516
rect 350476 306684 350532 306740
rect 349692 303212 349748 303268
rect 349356 300972 349412 301028
rect 349580 302540 349636 302596
rect 349244 300300 349300 300356
rect 350028 300188 350084 300244
rect 351036 308028 351092 308084
rect 351148 304556 351204 304612
rect 350588 300188 350644 300244
rect 350924 300972 350980 301028
rect 351484 304556 351540 304612
rect 352380 305676 352436 305732
rect 351932 304220 351988 304276
rect 352828 301644 352884 301700
rect 353164 306796 353220 306852
rect 351148 300972 351204 301028
rect 351820 301308 351876 301364
rect 351372 300748 351428 300804
rect 352268 300860 352324 300916
rect 354172 306796 354228 306852
rect 354620 306684 354676 306740
rect 353724 305452 353780 305508
rect 353276 301980 353332 302036
rect 354060 303548 354116 303604
rect 353612 299852 353668 299908
rect 355068 303436 355124 303492
rect 355404 306908 355460 306964
rect 354956 302988 355012 303044
rect 354508 302876 354564 302932
rect 355964 305676 356020 305732
rect 356188 304892 356244 304948
rect 355516 303212 355572 303268
rect 355852 304108 355908 304164
rect 356412 304892 356468 304948
rect 356188 304108 356244 304164
rect 356300 304780 356356 304836
rect 356860 304668 356916 304724
rect 357756 302204 357812 302260
rect 357308 302092 357364 302148
rect 357644 301868 357700 301924
rect 356748 301532 356804 301588
rect 357196 300972 357252 301028
rect 358092 301756 358148 301812
rect 358204 301532 358260 301588
rect 358540 307356 358596 307412
rect 358652 306908 358708 306964
rect 358988 303660 359044 303716
rect 359100 303548 359156 303604
rect 359436 303772 359492 303828
rect 359996 307356 360052 307412
rect 359548 303660 359604 303716
rect 359884 307132 359940 307188
rect 360332 303884 360388 303940
rect 360892 305676 360948 305732
rect 361340 302876 361396 302932
rect 361676 305004 361732 305060
rect 361788 304444 361844 304500
rect 360444 300524 360500 300580
rect 361676 302540 361732 302596
rect 360780 299964 360836 300020
rect 363132 307132 363188 307188
rect 363580 306236 363636 306292
rect 363916 307020 363972 307076
rect 362684 305564 362740 305620
rect 362236 301756 362292 301812
rect 363468 302428 363524 302484
rect 363020 301308 363076 301364
rect 362572 301196 362628 301252
rect 364028 303772 364084 303828
rect 340844 298284 340900 298340
rect 352716 298284 352772 298340
rect 361228 298284 361284 298340
rect 364364 307244 364420 307300
rect 364924 302764 364980 302820
rect 365260 303996 365316 304052
rect 364812 300748 364868 300804
rect 365820 305228 365876 305284
rect 366156 306348 366212 306404
rect 365372 300412 365428 300468
rect 365708 303324 365764 303380
rect 366268 305340 366324 305396
rect 366716 305004 366772 305060
rect 366828 305452 366884 305508
rect 366604 300076 366660 300132
rect 367164 305452 367220 305508
rect 367500 304108 367556 304164
rect 367612 302316 367668 302372
rect 367948 301420 368004 301476
rect 368060 300076 368116 300132
rect 368396 304332 368452 304388
rect 368508 304108 368564 304164
rect 368956 303884 369012 303940
rect 369292 306572 369348 306628
rect 368844 301084 368900 301140
rect 369404 305676 369460 305732
rect 369740 300300 369796 300356
rect 370300 305564 370356 305620
rect 370636 306460 370692 306516
rect 369852 299964 369908 300020
rect 370188 302876 370244 302932
rect 370748 305004 370804 305060
rect 364140 298284 364196 298340
rect 371420 307916 371476 307972
rect 371196 304220 371252 304276
rect 371308 304108 371364 304164
rect 371308 302876 371364 302932
rect 372540 306572 372596 306628
rect 372092 306460 372148 306516
rect 371644 305228 371700 305284
rect 372988 304892 373044 304948
rect 371980 303996 372036 304052
rect 371196 300860 371252 300916
rect 371084 300188 371140 300244
rect 373884 304556 373940 304612
rect 374220 305116 374276 305172
rect 373436 303324 373492 303380
rect 373772 301980 373828 302036
rect 373324 301644 373380 301700
rect 372876 300860 372932 300916
rect 372428 300748 372484 300804
rect 374332 302092 374388 302148
rect 374668 306796 374724 306852
rect 374780 306348 374836 306404
rect 375116 306684 375172 306740
rect 375228 304780 375284 304836
rect 375676 303996 375732 304052
rect 375340 303212 375396 303268
rect 376012 303100 376068 303156
rect 376572 307020 376628 307076
rect 376236 304556 376292 304612
rect 376236 303436 376292 303492
rect 376460 304108 376516 304164
rect 376124 301644 376180 301700
rect 376908 300860 376964 300916
rect 377244 304444 377300 304500
rect 378812 307244 378868 307300
rect 377916 305676 377972 305732
rect 379148 306908 379204 306964
rect 377468 303212 377524 303268
rect 378252 302204 378308 302260
rect 377244 300860 377300 300916
rect 377804 301980 377860 302036
rect 377020 299852 377076 299908
rect 377356 300748 377412 300804
rect 378700 301532 378756 301588
rect 379260 301532 379316 301588
rect 379596 303548 379652 303604
rect 380156 304556 380212 304612
rect 380492 307356 380548 307412
rect 379708 301868 379764 301924
rect 380044 303660 380100 303716
rect 381500 306684 381556 306740
rect 381052 305676 381108 305732
rect 380604 303996 380660 304052
rect 382396 306796 382452 306852
rect 381948 303548 382004 303604
rect 381388 303100 381444 303156
rect 380940 300524 380996 300580
rect 382732 301756 382788 301812
rect 381836 301308 381892 301364
rect 382284 300860 382340 300916
rect 383292 307356 383348 307412
rect 383628 307132 383684 307188
rect 382844 300188 382900 300244
rect 383180 300748 383236 300804
rect 384076 306236 384132 306292
rect 383964 303996 384020 304052
rect 383964 302092 384020 302148
rect 383740 301756 383796 301812
rect 384188 304444 384244 304500
rect 384524 303772 384580 303828
rect 385084 308028 385140 308084
rect 385532 306908 385588 306964
rect 384636 301980 384692 302036
rect 385420 302988 385476 303044
rect 386428 303100 386484 303156
rect 386764 305340 386820 305396
rect 385980 300524 386036 300580
rect 386316 301420 386372 301476
rect 385868 300412 385924 300468
rect 386876 303772 386932 303828
rect 387324 302764 387380 302820
rect 387660 305116 387716 305172
rect 387212 302428 387268 302484
rect 387772 304780 387828 304836
rect 388108 305564 388164 305620
rect 388108 303996 388164 304052
rect 388108 300748 388164 300804
rect 389116 305116 389172 305172
rect 388668 304668 388724 304724
rect 389452 303884 389508 303940
rect 388220 300300 388276 300356
rect 389004 302876 389060 302932
rect 388556 300076 388612 300132
rect 390012 303772 390068 303828
rect 389564 302204 389620 302260
rect 389900 303100 389956 303156
rect 390460 300076 390516 300132
rect 390796 303996 390852 304052
rect 390348 299964 390404 300020
rect 390908 303884 390964 303940
rect 391244 305004 391300 305060
rect 392252 307132 392308 307188
rect 391804 306236 391860 306292
rect 392588 306460 392644 306516
rect 391356 304220 391412 304276
rect 392140 305228 392196 305284
rect 392700 305676 392756 305732
rect 393036 306572 393092 306628
rect 394044 305564 394100 305620
rect 393596 305452 393652 305508
rect 393148 305340 393204 305396
rect 394492 305228 394548 305284
rect 393484 304892 393540 304948
rect 394828 304780 394884 304836
rect 393820 304556 393876 304612
rect 393708 303324 393764 303380
rect 393932 304444 393988 304500
rect 393932 301420 393988 301476
rect 394380 303436 394436 303492
rect 393820 301308 393876 301364
rect 394940 303436 394996 303492
rect 395276 306348 395332 306404
rect 394828 302204 394884 302260
rect 394828 300748 394884 300804
rect 395836 305228 395892 305284
rect 395388 305004 395444 305060
rect 395724 303996 395780 304052
rect 395948 303996 396004 304052
rect 395948 303660 396004 303716
rect 396172 303660 396228 303716
rect 398860 308028 398916 308084
rect 396732 304892 396788 304948
rect 397068 307020 397124 307076
rect 396284 303324 396340 303380
rect 396172 302988 396228 303044
rect 396172 302316 396228 302372
rect 396620 301644 396676 301700
rect 397964 303212 398020 303268
rect 397516 299852 397572 299908
rect 398412 303100 398468 303156
rect 405580 307916 405636 307972
rect 403788 307356 403844 307412
rect 399308 307244 399364 307300
rect 402892 306796 402948 306852
rect 401996 306684 402052 306740
rect 401548 304108 401604 304164
rect 401100 302092 401156 302148
rect 400204 301868 400260 301924
rect 399756 301532 399812 301588
rect 400652 301308 400708 301364
rect 402332 304668 402388 304724
rect 402332 302428 402388 302484
rect 402444 303548 402500 303604
rect 403340 300188 403396 300244
rect 405132 301980 405188 302036
rect 404236 301756 404292 301812
rect 404684 301420 404740 301476
rect 411516 307468 411572 307524
rect 406028 306908 406084 306964
rect 409612 305116 409668 305172
rect 407372 303996 407428 304052
rect 406924 303660 406980 303716
rect 406476 300524 406532 300580
rect 407820 302988 407876 303044
rect 409164 302428 409220 302484
rect 408268 302204 408324 302260
rect 408716 300300 408772 300356
rect 418348 307468 418404 307524
rect 412748 307132 412804 307188
rect 411516 304108 411572 304164
rect 412300 306236 412356 306292
rect 411404 303884 411460 303940
rect 410508 303772 410564 303828
rect 410060 300748 410116 300804
rect 410956 300076 411012 300132
rect 411852 302876 411908 302932
rect 413196 305676 413252 305732
rect 414540 305564 414596 305620
rect 414092 305452 414148 305508
rect 413644 305340 413700 305396
rect 416332 305228 416388 305284
rect 415884 305004 415940 305060
rect 415436 303436 415492 303492
rect 414988 300748 415044 300804
rect 417228 304892 417284 304948
rect 416780 303324 416836 303380
rect 370860 298284 370916 298340
rect 384972 298284 385028 298340
rect 391692 298284 391748 298340
rect 319004 95004 319060 95060
rect 423276 320908 423332 320964
rect 423276 314188 423332 314244
rect 420140 299068 420196 299124
rect 420028 298060 420084 298116
rect 420140 285628 420196 285684
rect 420028 258636 420084 258692
rect 419132 94892 419188 94948
rect 421596 89852 421652 89908
rect 318892 86828 318948 86884
rect 351036 88060 351092 88116
rect 318332 86716 318388 86772
rect 319116 86156 319172 86212
rect 315644 84924 315700 84980
rect 315756 85260 315812 85316
rect 301756 83468 301812 83524
rect 314972 84476 315028 84532
rect 299180 83132 299236 83188
rect 298620 81676 298676 81732
rect 292236 80444 292292 80500
rect 295596 81228 295652 81284
rect 287196 78316 287252 78372
rect 295596 78204 295652 78260
rect 317324 84588 317380 84644
rect 317324 83804 317380 83860
rect 317436 84476 317492 84532
rect 319116 83916 319172 83972
rect 340956 86044 341012 86100
rect 317436 83692 317492 83748
rect 421596 87276 421652 87332
rect 414988 86044 415044 86100
rect 414988 83916 415044 83972
rect 422828 84252 422884 84308
rect 351036 83580 351092 83636
rect 340956 83468 341012 83524
rect 315756 83244 315812 83300
rect 419132 83244 419188 83300
rect 416668 82572 416724 82628
rect 416668 81452 416724 81508
rect 422828 82236 422884 82292
rect 427084 392588 427140 392644
rect 428428 392588 428484 392644
rect 428428 391356 428484 391412
rect 443212 391132 443268 391188
rect 439180 391020 439236 391076
rect 435148 390684 435204 390740
rect 446796 390460 446852 390516
rect 431116 387772 431172 387828
rect 442652 389340 442708 389396
rect 430892 383852 430948 383908
rect 429212 380492 429268 380548
rect 425852 373772 425908 373828
rect 424396 372092 424452 372148
rect 424956 340956 425012 341012
rect 424956 333452 425012 333508
rect 425068 324268 425124 324324
rect 425068 320908 425124 320964
rect 425180 84812 425236 84868
rect 425068 83132 425124 83188
rect 425068 80556 425124 80612
rect 425180 80444 425236 80500
rect 426748 368844 426804 368900
rect 426748 362796 426804 362852
rect 427532 368732 427588 368788
rect 427532 340956 427588 341012
rect 428764 92764 428820 92820
rect 425852 80332 425908 80388
rect 428204 82684 428260 82740
rect 424396 80220 424452 80276
rect 424172 80108 424228 80164
rect 419132 78428 419188 78484
rect 314972 78204 315028 78260
rect 270620 77084 270676 77140
rect 270284 23100 270340 23156
rect 269836 18508 269892 18564
rect 269724 16156 269780 16212
rect 270396 16716 270452 16772
rect 269948 15708 270004 15764
rect 269612 13356 269668 13412
rect 269724 13692 269780 13748
rect 269500 7980 269556 8036
rect 268940 6524 268996 6580
rect 269836 12572 269892 12628
rect 269948 10332 270004 10388
rect 270284 13580 270340 13636
rect 269724 6412 269780 6468
rect 269836 9884 269892 9940
rect 269948 5740 270004 5796
rect 270172 8204 270228 8260
rect 270172 4396 270228 4452
rect 269836 1596 269892 1652
rect 268492 1372 268548 1428
rect 270620 14476 270676 14532
rect 270396 4284 270452 4340
rect 270508 11116 270564 11172
rect 270508 3164 270564 3220
rect 275324 10444 275380 10500
rect 275212 9996 275268 10052
rect 275212 5292 275268 5348
rect 312396 10444 312452 10500
rect 287084 10332 287140 10388
rect 277228 9772 277284 9828
rect 275436 6972 275492 7028
rect 275436 5180 275492 5236
rect 275660 5292 275716 5348
rect 275324 4396 275380 4452
rect 275548 5068 275604 5124
rect 274092 4284 274148 4340
rect 270620 476 270676 532
rect 272188 4172 272244 4228
rect 275548 2492 275604 2548
rect 277564 9100 277620 9156
rect 277452 8764 277508 8820
rect 277340 8652 277396 8708
rect 277340 8316 277396 8372
rect 277228 4844 277284 4900
rect 275996 3948 276052 4004
rect 275772 3500 275828 3556
rect 275772 3164 275828 3220
rect 275660 2044 275716 2100
rect 277452 3052 277508 3108
rect 279132 8540 279188 8596
rect 278908 8428 278964 8484
rect 277564 2380 277620 2436
rect 277900 6188 277956 6244
rect 278908 3276 278964 3332
rect 283612 8204 283668 8260
rect 280812 6972 280868 7028
rect 280812 6300 280868 6356
rect 281708 6860 281764 6916
rect 279132 1372 279188 1428
rect 279804 4844 279860 4900
rect 280476 3612 280532 3668
rect 280364 2716 280420 2772
rect 280476 1596 280532 1652
rect 280364 1036 280420 1092
rect 282156 3724 282212 3780
rect 282156 1596 282212 1652
rect 285852 6972 285908 7028
rect 285628 6860 285684 6916
rect 285628 6412 285684 6468
rect 285740 5180 285796 5236
rect 285628 3724 285684 3780
rect 310716 10108 310772 10164
rect 290668 8764 290724 8820
rect 288988 8652 289044 8708
rect 288988 8316 289044 8372
rect 289100 8540 289156 8596
rect 289100 6636 289156 6692
rect 297164 8764 297220 8820
rect 290668 6636 290724 6692
rect 293132 8092 293188 8148
rect 287084 6300 287140 6356
rect 291228 5964 291284 6020
rect 287308 4844 287364 4900
rect 285740 3052 285796 3108
rect 286076 2604 286132 2660
rect 285628 2268 285684 2324
rect 287308 2156 287364 2212
rect 287420 3612 287476 3668
rect 285404 476 285460 532
rect 289324 2716 289380 2772
rect 295820 6972 295876 7028
rect 295820 6636 295876 6692
rect 304108 8652 304164 8708
rect 297164 6412 297220 6468
rect 302652 7084 302708 7140
rect 295372 6188 295428 6244
rect 294028 3164 294084 3220
rect 294028 1372 294084 1428
rect 295036 2380 295092 2436
rect 300748 5740 300804 5796
rect 295372 2380 295428 2436
rect 295484 5180 295540 5236
rect 296492 5068 296548 5124
rect 296492 4844 296548 4900
rect 298844 4844 298900 4900
rect 295484 2044 295540 2100
rect 296940 4396 296996 4452
rect 297388 3724 297444 3780
rect 297388 2828 297444 2884
rect 297612 3500 297668 3556
rect 297612 2716 297668 2772
rect 303996 6860 304052 6916
rect 303996 5068 304052 5124
rect 308364 6524 308420 6580
rect 304108 3276 304164 3332
rect 307356 5068 307412 5124
rect 307356 3164 307412 3220
rect 304556 2604 304612 2660
rect 308252 2604 308308 2660
rect 308252 2380 308308 2436
rect 305676 1932 305732 1988
rect 305676 1484 305732 1540
rect 306796 476 306852 532
rect 310716 5964 310772 6020
rect 310268 3724 310324 3780
rect 309148 3500 309204 3556
rect 309148 1932 309204 1988
rect 420700 10444 420756 10500
rect 413084 10332 413140 10388
rect 314188 9884 314244 9940
rect 365484 9660 365540 9716
rect 331212 9548 331268 9604
rect 319788 7980 319844 8036
rect 318108 4396 318164 4452
rect 315980 3388 316036 3444
rect 324268 5180 324324 5236
rect 320908 4732 320964 4788
rect 323820 3724 323876 3780
rect 320908 2828 320964 2884
rect 321692 3500 321748 3556
rect 324268 3164 324324 3220
rect 327404 4284 327460 4340
rect 325500 2716 325556 2772
rect 329532 4284 329588 4340
rect 336924 9436 336980 9492
rect 333116 4508 333172 4564
rect 335244 4508 335300 4564
rect 358092 9436 358148 9492
rect 342748 9324 342804 9380
rect 340956 6188 341012 6244
rect 338828 1708 338884 1764
rect 346668 9324 346724 9380
rect 344540 4620 344596 4676
rect 357196 8540 357252 8596
rect 357196 8204 357252 8260
rect 354060 6972 354116 7028
rect 348348 6412 348404 6468
rect 350252 6300 350308 6356
rect 352716 4172 352772 4228
rect 352380 4060 352436 4116
rect 352716 2716 352772 2772
rect 355964 3052 356020 3108
rect 361676 8204 361732 8260
rect 359772 6076 359828 6132
rect 363804 6972 363860 7028
rect 362796 6076 362852 6132
rect 362796 4060 362852 4116
rect 398188 9660 398244 9716
rect 370412 9548 370468 9604
rect 398076 7980 398132 8036
rect 370412 6972 370468 7028
rect 376908 7868 376964 7924
rect 373100 6860 373156 6916
rect 367388 4732 367444 4788
rect 369516 3388 369572 3444
rect 371308 3164 371364 3220
rect 375228 3612 375284 3668
rect 380940 7868 380996 7924
rect 378812 3500 378868 3556
rect 382620 7756 382676 7812
rect 386652 7756 386708 7812
rect 390460 6860 390516 6916
rect 384412 364 384468 420
rect 388332 5852 388388 5908
rect 394828 6412 394884 6468
rect 392364 5852 392420 5908
rect 394828 4396 394884 4452
rect 394044 3388 394100 3444
rect 397740 3388 397796 3444
rect 397740 476 397796 532
rect 398188 6860 398244 6916
rect 399868 9212 399924 9268
rect 398076 3612 398132 3668
rect 398076 1596 398132 1652
rect 408268 9212 408324 9268
rect 403788 8092 403844 8148
rect 401884 6300 401940 6356
rect 408268 6412 408324 6468
rect 411180 6748 411236 6804
rect 407596 4396 407652 4452
rect 406588 3388 406644 3444
rect 395836 252 395892 308
rect 405468 2940 405524 2996
rect 406588 1484 406644 1540
rect 409500 4172 409556 4228
rect 413196 8204 413252 8260
rect 419020 4844 419076 4900
rect 417116 4732 417172 4788
rect 413196 4508 413252 4564
rect 415212 4508 415268 4564
rect 416668 3724 416724 3780
rect 416668 3052 416724 3108
rect 428204 9660 428260 9716
rect 428428 7644 428484 7700
rect 425068 6748 425124 6804
rect 425068 4732 425124 4788
rect 420700 4396 420756 4452
rect 422604 4172 422660 4228
rect 420924 4060 420980 4116
rect 424508 4172 424564 4228
rect 426636 4172 426692 4228
rect 428988 84364 429044 84420
rect 428988 34412 429044 34468
rect 429100 82460 429156 82516
rect 429324 338604 429380 338660
rect 429324 324268 429380 324324
rect 430108 299292 430164 299348
rect 429660 89068 429716 89124
rect 429436 87836 429492 87892
rect 429212 79996 429268 80052
rect 429324 84588 429380 84644
rect 429100 14588 429156 14644
rect 428764 6748 428820 6804
rect 429436 7980 429492 8036
rect 429548 82572 429604 82628
rect 429660 22652 429716 22708
rect 429884 84924 429940 84980
rect 429996 80444 430052 80500
rect 429996 22764 430052 22820
rect 429884 14700 429940 14756
rect 429548 5852 429604 5908
rect 429324 4284 429380 4340
rect 430220 298396 430276 298452
rect 430220 4172 430276 4228
rect 430332 87276 430388 87332
rect 430108 4060 430164 4116
rect 434252 375452 434308 375508
rect 430892 79884 430948 79940
rect 431004 95900 431060 95956
rect 430892 78428 430948 78484
rect 432796 94556 432852 94612
rect 432572 94108 432628 94164
rect 431004 20076 431060 20132
rect 431116 92652 431172 92708
rect 431116 18396 431172 18452
rect 431228 86044 431284 86100
rect 430892 11228 430948 11284
rect 431452 83468 431508 83524
rect 432572 18172 432628 18228
rect 432684 87612 432740 87668
rect 432796 19516 432852 19572
rect 432908 92540 432964 92596
rect 434028 83580 434084 83636
rect 433020 80668 433076 80724
rect 433020 31948 433076 32004
rect 432908 17948 432964 18004
rect 432684 14812 432740 14868
rect 431452 11116 431508 11172
rect 431228 10892 431284 10948
rect 432124 4172 432180 4228
rect 435932 372988 435988 373044
rect 440188 372428 440244 372484
rect 436044 372316 436100 372372
rect 437612 372204 437668 372260
rect 437612 368844 437668 368900
rect 440188 368732 440244 368788
rect 436044 338604 436100 338660
rect 435932 93212 435988 93268
rect 437612 296940 437668 296996
rect 434252 79772 434308 79828
rect 435932 90748 435988 90804
rect 434476 79212 434532 79268
rect 434476 19628 434532 19684
rect 435932 17836 435988 17892
rect 436044 87500 436100 87556
rect 436716 85932 436772 85988
rect 436268 85820 436324 85876
rect 436044 16380 436100 16436
rect 436156 84476 436212 84532
rect 436716 16492 436772 16548
rect 436268 16268 436324 16324
rect 436156 13132 436212 13188
rect 435932 12572 435988 12628
rect 439740 100828 439796 100884
rect 439404 94220 439460 94276
rect 437724 92428 437780 92484
rect 439292 90860 439348 90916
rect 437724 19404 437780 19460
rect 437836 29372 437892 29428
rect 438508 17612 438564 17668
rect 438508 15036 438564 15092
rect 437836 14476 437892 14532
rect 439404 17724 439460 17780
rect 439516 80892 439572 80948
rect 439516 16604 439572 16660
rect 439292 7868 439348 7924
rect 437612 4508 437668 4564
rect 437836 4172 437892 4228
rect 446796 386316 446852 386372
rect 443212 386092 443268 386148
rect 442764 373212 442820 373268
rect 442876 371420 442932 371476
rect 443100 371308 443156 371364
rect 442876 100604 442932 100660
rect 442988 370636 443044 370692
rect 442764 96572 442820 96628
rect 442876 97468 442932 97524
rect 442652 93996 442708 94052
rect 442764 94332 442820 94388
rect 442652 88508 442708 88564
rect 442428 80780 442484 80836
rect 441644 34412 441700 34468
rect 439964 22764 440020 22820
rect 440076 22652 440132 22708
rect 440076 19180 440132 19236
rect 439964 15820 440020 15876
rect 441868 15036 441924 15092
rect 442428 13356 442484 13412
rect 442652 13020 442708 13076
rect 441868 11004 441924 11060
rect 451276 390460 451332 390516
rect 459340 389564 459396 389620
rect 463372 389452 463428 389508
rect 455308 386204 455364 386260
rect 447244 384188 447300 384244
rect 467404 384076 467460 384132
rect 479500 393036 479556 393092
rect 475468 392140 475524 392196
rect 483532 390908 483588 390964
rect 491596 387548 491652 387604
rect 487564 385980 487620 386036
rect 499660 389228 499716 389284
rect 495628 385868 495684 385924
rect 511756 392476 511812 392532
rect 507724 387436 507780 387492
rect 519820 392364 519876 392420
rect 523852 390796 523908 390852
rect 515788 387324 515844 387380
rect 503692 385756 503748 385812
rect 535948 392252 536004 392308
rect 531916 389116 531972 389172
rect 544012 392588 544068 392644
rect 539980 387212 540036 387268
rect 527884 385644 527940 385700
rect 471436 383964 471492 384020
rect 562604 380604 562660 380660
rect 587132 575372 587188 575428
rect 587244 535724 587300 535780
rect 590828 522508 590884 522564
rect 590492 469644 590548 469700
rect 587244 388892 587300 388948
rect 590380 403564 590436 403620
rect 587132 385532 587188 385588
rect 584668 378812 584724 378868
rect 544236 374556 544292 374612
rect 535052 373884 535108 373940
rect 535052 372428 535108 372484
rect 590380 373772 590436 373828
rect 544236 372316 544292 372372
rect 590716 456428 590772 456484
rect 590604 443212 590660 443268
rect 591052 496076 591108 496132
rect 590828 394268 590884 394324
rect 590940 430108 590996 430164
rect 590716 390684 590772 390740
rect 591276 482860 591332 482916
rect 591052 394156 591108 394212
rect 591164 416780 591220 416836
rect 591276 393932 591332 393988
rect 591164 383852 591220 383908
rect 590940 380492 590996 380548
rect 590604 375452 590660 375508
rect 591052 373212 591108 373268
rect 590492 372092 590548 372148
rect 590604 373100 590660 373156
rect 590492 370636 590548 370692
rect 590828 372988 590884 373044
rect 590604 337596 590660 337652
rect 590716 371420 590772 371476
rect 590492 311276 590548 311332
rect 590828 350924 590884 350980
rect 590940 371308 590996 371364
rect 591052 364140 591108 364196
rect 590940 324492 590996 324548
rect 590716 298060 590772 298116
rect 443212 296492 443268 296548
rect 443996 296828 444052 296884
rect 443100 99932 443156 99988
rect 442988 96684 443044 96740
rect 443212 97692 443268 97748
rect 442876 19292 442932 19348
rect 442988 89964 443044 90020
rect 443100 86268 443156 86324
rect 443100 12908 443156 12964
rect 442988 8092 443044 8148
rect 442764 7084 442820 7140
rect 444108 97580 444164 97636
rect 443436 94444 443492 94500
rect 443324 84028 443380 84084
rect 443324 12796 443380 12852
rect 443436 4396 443492 4452
rect 443548 90076 443604 90132
rect 443212 4172 443268 4228
rect 444108 7756 444164 7812
rect 587132 284620 587188 284676
rect 464492 19180 464548 19236
rect 460684 17500 460740 17556
rect 447356 15820 447412 15876
rect 444220 4620 444276 4676
rect 445452 7532 445508 7588
rect 458780 13356 458836 13412
rect 449260 8092 449316 8148
rect 456988 7980 457044 8036
rect 451164 5964 451220 6020
rect 454972 4844 455028 4900
rect 462588 5852 462644 5908
rect 587356 271404 587412 271460
rect 587244 178892 587300 178948
rect 587244 19404 587300 19460
rect 587580 218540 587636 218596
rect 587468 99596 587524 99652
rect 587468 19516 587524 19572
rect 587356 18172 587412 18228
rect 590828 165676 590884 165732
rect 587804 139244 587860 139300
rect 590492 112812 590548 112868
rect 590268 59948 590324 60004
rect 590044 46732 590100 46788
rect 589820 33628 589876 33684
rect 589820 19964 589876 20020
rect 590268 20076 590324 20132
rect 590044 19628 590100 19684
rect 587804 18060 587860 18116
rect 587580 17948 587636 18004
rect 590828 20860 590884 20916
rect 590940 152460 590996 152516
rect 591052 126028 591108 126084
rect 591276 86380 591332 86436
rect 591052 20972 591108 21028
rect 591164 73164 591220 73220
rect 590940 19852 590996 19908
rect 590492 17836 590548 17892
rect 591276 20636 591332 20692
rect 591276 20300 591332 20356
rect 591276 18396 591332 18452
rect 591164 17724 591220 17780
rect 587132 17612 587188 17668
rect 487340 16716 487396 16772
rect 472108 13244 472164 13300
rect 468300 11228 468356 11284
rect 466396 4732 466452 4788
rect 470204 588 470260 644
rect 481628 13132 481684 13188
rect 477820 4508 477876 4564
rect 475916 1708 475972 1764
rect 474012 588 474068 644
rect 479724 4060 479780 4116
rect 483532 4620 483588 4676
rect 485548 588 485604 644
rect 491148 16604 491204 16660
rect 489244 2828 489300 2884
rect 514108 16492 514164 16548
rect 508284 14812 508340 14868
rect 493052 13020 493108 13076
rect 498764 12908 498820 12964
rect 496860 4396 496916 4452
rect 494956 2604 495012 2660
rect 504476 12796 504532 12852
rect 500668 7868 500724 7924
rect 502572 2492 502628 2548
rect 506380 3388 506436 3444
rect 510188 12684 510244 12740
rect 512092 3388 512148 3444
rect 525420 16380 525476 16436
rect 519708 14700 519764 14756
rect 514220 8428 514276 8484
rect 514220 6748 514276 6804
rect 517804 3388 517860 3444
rect 515900 1708 515956 1764
rect 521612 6748 521668 6804
rect 523516 4284 523572 4340
rect 538748 16268 538804 16324
rect 529228 14588 529284 14644
rect 527324 588 527380 644
rect 531132 4284 531188 4340
rect 534940 3388 534996 3444
rect 533036 588 533092 644
rect 536844 2716 536900 2772
rect 565404 16156 565460 16212
rect 546812 14476 546868 14532
rect 544460 11116 544516 11172
rect 540652 3948 540708 4004
rect 542668 1708 542724 1764
rect 561596 11004 561652 11060
rect 552076 7756 552132 7812
rect 546812 4956 546868 5012
rect 550172 4956 550228 5012
rect 548268 4284 548324 4340
rect 546364 3836 546420 3892
rect 557788 3724 557844 3780
rect 555884 3388 555940 3444
rect 553980 588 554036 644
rect 559692 3388 559748 3444
rect 563500 10892 563556 10948
rect 567308 16044 567364 16100
rect 578732 15932 578788 15988
rect 569212 14364 569268 14420
rect 576828 14252 576884 14308
rect 574924 6748 574980 6804
rect 573020 4172 573076 4228
rect 571228 3388 571284 3444
rect 584444 12572 584500 12628
rect 580636 7644 580692 7700
rect 582540 4172 582596 4228
rect 452956 140 453012 196
<< metal3 >>
rect 540754 591052 540764 591108
rect 540820 591052 549388 591108
rect 549444 591052 549454 591108
rect 19170 590940 19180 590996
rect 19236 590940 33068 590996
rect 33124 590940 33134 590996
rect 518690 590940 518700 590996
rect 518756 590940 548044 590996
rect 548100 590940 548110 590996
rect 29474 590828 29484 590884
rect 29540 590828 55132 590884
rect 55188 590828 55198 590884
rect 496626 590828 496636 590884
rect 496692 590828 548156 590884
rect 548212 590828 548222 590884
rect 28354 590716 28364 590772
rect 28420 590716 77308 590772
rect 77364 590716 77374 590772
rect 474562 590716 474572 590772
rect 474628 590716 547708 590772
rect 547764 590716 547774 590772
rect 26786 590604 26796 590660
rect 26852 590604 99260 590660
rect 99316 590604 99326 590660
rect 452498 590604 452508 590660
rect 452564 590604 549612 590660
rect 549668 590604 549678 590660
rect 28466 590492 28476 590548
rect 28532 590492 143388 590548
rect 143444 590492 143454 590548
rect 242722 590492 242732 590548
rect 242788 590492 253708 590548
rect 253764 590492 253774 590548
rect 336802 590492 336812 590548
rect 336868 590492 341964 590548
rect 342020 590492 342030 590548
rect 364242 590492 364252 590548
rect 364308 590492 380492 590548
rect 380548 590492 380558 590548
rect 430434 590492 430444 590548
rect 430500 590492 548268 590548
rect 548324 590492 548334 590548
rect 162082 590156 162092 590212
rect 162148 590156 165452 590212
rect 165508 590156 165518 590212
rect 225922 590156 225932 590212
rect 225988 590156 231644 590212
rect 231700 590156 231710 590212
rect 317538 590156 317548 590212
rect 317604 590156 319900 590212
rect 319956 590156 319966 590212
rect 595560 588644 597000 588840
rect 590482 588588 590492 588644
rect 590548 588616 597000 588644
rect 590548 588588 595672 588616
rect 295586 587916 295596 587972
rect 295652 587916 297836 587972
rect 297892 587916 297902 587972
rect 314178 587916 314188 587972
rect 314244 587916 317548 587972
rect 317604 587916 317614 587972
rect -960 587188 480 587384
rect -960 587160 3388 587188
rect 392 587132 3388 587160
rect 3444 587132 3454 587188
rect 193218 583772 193228 583828
rect 193284 583772 209580 583828
rect 209636 583772 209646 583828
rect 268706 582988 268716 583044
rect 268772 582988 275772 583044
rect 275828 582988 275838 583044
rect 292226 581308 292236 581364
rect 292292 581308 295596 581364
rect 295652 581308 295662 581364
rect 386082 581308 386092 581364
rect 386148 581308 394828 581364
rect 394884 581308 394894 581364
rect 310818 579516 310828 579572
rect 310884 579516 314076 579572
rect 314132 579516 314142 579572
rect 188066 579292 188076 579348
rect 188132 579292 193228 579348
rect 193284 579292 193294 579348
rect 380482 577836 380492 577892
rect 380548 577836 383068 577892
rect 383124 577836 383134 577892
rect 29362 577276 29372 577332
rect 29428 577276 121324 577332
rect 121380 577276 121390 577332
rect 169698 577276 169708 577332
rect 169764 577276 187516 577332
rect 187572 577276 187582 577332
rect 29250 577164 29260 577220
rect 29316 577164 310828 577220
rect 310884 577164 310894 577220
rect 28466 577052 28476 577108
rect 28532 577052 336812 577108
rect 336868 577052 336878 577108
rect 223132 576268 225932 576324
rect 225988 576268 225998 576324
rect 28018 576044 28028 576100
rect 28084 576044 162092 576100
rect 162148 576044 162158 576100
rect 29250 575932 29260 575988
rect 29316 575932 169708 575988
rect 169764 575932 169774 575988
rect 29138 575820 29148 575876
rect 29204 575820 188076 575876
rect 188132 575820 188142 575876
rect 223132 575764 223188 576268
rect 28130 575708 28140 575764
rect 28196 575708 223188 575764
rect 29026 575596 29036 575652
rect 29092 575596 242732 575652
rect 242788 575596 242798 575652
rect 408258 575596 408268 575652
rect 408324 575596 547820 575652
rect 547876 575596 547886 575652
rect 28242 575484 28252 575540
rect 28308 575484 268716 575540
rect 268772 575484 268782 575540
rect 394818 575484 394828 575540
rect 394884 575484 549500 575540
rect 549556 575484 549566 575540
rect 595560 575428 597000 575624
rect 26450 575372 26460 575428
rect 26516 575372 292236 575428
rect 292292 575372 292302 575428
rect 383058 575372 383068 575428
rect 383124 575372 547932 575428
rect 547988 575372 547998 575428
rect 587122 575372 587132 575428
rect 587188 575400 597000 575428
rect 587188 575372 595672 575400
rect 26562 575036 26572 575092
rect 26628 575036 29260 575092
rect 29316 575036 29326 575092
rect 26674 574476 26684 574532
rect 26740 574476 28476 574532
rect 28532 574476 28542 574532
rect -960 573076 480 573272
rect -960 573048 12572 573076
rect 392 573020 12572 573048
rect 12628 573020 12638 573076
rect 595560 562212 597000 562408
rect 590594 562156 590604 562212
rect 590660 562184 597000 562212
rect 590660 562156 595672 562184
rect -960 558964 480 559160
rect -960 558936 3500 558964
rect 392 558908 3500 558936
rect 3556 558908 3566 558964
rect 595560 548996 597000 549192
rect 590706 548940 590716 548996
rect 590772 548968 597000 548996
rect 590772 548940 595672 548968
rect -960 544852 480 545048
rect -960 544824 4172 544852
rect 392 544796 4172 544824
rect 4228 544796 4238 544852
rect 595560 535780 597000 535976
rect 587234 535724 587244 535780
rect 587300 535752 597000 535780
rect 587300 535724 595672 535752
rect -960 530740 480 530936
rect -960 530712 14252 530740
rect 392 530684 14252 530712
rect 14308 530684 14318 530740
rect 595560 522564 597000 522760
rect 590818 522508 590828 522564
rect 590884 522536 597000 522564
rect 590884 522508 595672 522536
rect -960 516628 480 516824
rect -960 516600 4284 516628
rect 392 516572 4284 516600
rect 4340 516572 4350 516628
rect 595560 509348 597000 509544
rect 590818 509292 590828 509348
rect 590884 509320 597000 509348
rect 590884 509292 595672 509320
rect -960 502516 480 502712
rect -960 502488 4396 502516
rect 392 502460 4396 502488
rect 4452 502460 4462 502516
rect 595560 496132 597000 496328
rect 591042 496076 591052 496132
rect 591108 496104 597000 496132
rect 591108 496076 595672 496104
rect -960 488404 480 488600
rect -960 488376 4508 488404
rect 392 488348 4508 488376
rect 4564 488348 4574 488404
rect 595560 482916 597000 483112
rect 591266 482860 591276 482916
rect 591332 482888 597000 482916
rect 591332 482860 595672 482888
rect -960 474292 480 474488
rect -960 474264 4732 474292
rect 392 474236 4732 474264
rect 4788 474236 4798 474292
rect 595560 469700 597000 469896
rect 590482 469644 590492 469700
rect 590548 469672 597000 469700
rect 590548 469644 595672 469672
rect -960 460180 480 460376
rect -960 460152 4620 460180
rect 392 460124 4620 460152
rect 4676 460124 4686 460180
rect 595560 456484 597000 456680
rect 590706 456428 590716 456484
rect 590772 456456 597000 456484
rect 590772 456428 595672 456456
rect -960 446068 480 446264
rect -960 446040 17612 446068
rect 392 446012 17612 446040
rect 17668 446012 17678 446068
rect 595560 443268 597000 443464
rect 590594 443212 590604 443268
rect 590660 443240 597000 443268
rect 590660 443212 595672 443240
rect -960 431956 480 432152
rect -960 431928 4844 431956
rect 392 431900 4844 431928
rect 4900 431900 4910 431956
rect 595560 430164 597000 430248
rect 590930 430108 590940 430164
rect 590996 430108 597000 430164
rect 595560 430024 597000 430108
rect -960 417844 480 418040
rect -960 417816 3948 417844
rect 392 417788 3948 417816
rect 4004 417788 4014 417844
rect 595560 416836 597000 417032
rect 591154 416780 591164 416836
rect 591220 416808 597000 416836
rect 591220 416780 595672 416808
rect 3378 416668 3388 416724
rect 3444 416668 4844 416724
rect 4900 416668 4910 416724
rect -960 403732 480 403928
rect -960 403704 4956 403732
rect 392 403676 4956 403704
rect 5012 403676 5022 403732
rect 595560 403620 597000 403816
rect 590370 403564 590380 403620
rect 590436 403592 597000 403620
rect 590436 403564 595672 403592
rect 3490 403228 3500 403284
rect 3556 403228 4956 403284
rect 5012 403228 5022 403284
rect 28018 394492 28028 394548
rect 28084 394492 30268 394548
rect 30324 394492 30334 394548
rect 4834 394380 4844 394436
rect 4900 394380 152236 394436
rect 152292 394380 152302 394436
rect 4386 394268 4396 394324
rect 4452 394268 152012 394324
rect 152068 394268 152078 394324
rect 156930 394268 156940 394324
rect 156996 394268 235676 394324
rect 235732 394268 235742 394324
rect 442642 394268 442652 394324
rect 442708 394268 590828 394324
rect 590884 394268 590894 394324
rect 4834 394156 4844 394212
rect 4900 394156 162092 394212
rect 162148 394156 162158 394212
rect 437602 394156 437612 394212
rect 437668 394156 591052 394212
rect 591108 394156 591118 394212
rect 4162 394044 4172 394100
rect 4228 394044 162316 394100
rect 162372 394044 162382 394100
rect 427522 394044 427532 394100
rect 427588 394044 590604 394100
rect 590660 394044 590670 394100
rect 3938 393932 3948 393988
rect 4004 393932 166012 393988
rect 166068 393932 166078 393988
rect 424162 393932 424172 393988
rect 424228 393932 591276 393988
rect 591332 393932 591342 393988
rect 28130 393148 28140 393204
rect 28196 393148 30156 393204
rect 30212 393148 30222 393204
rect 130956 393148 208796 393204
rect 208852 393148 208862 393204
rect 130956 393092 131012 393148
rect 26450 393036 26460 393092
rect 26516 393036 28476 393092
rect 28532 393036 28542 393092
rect 96450 393036 96460 393092
rect 96516 393036 131012 393092
rect 381378 393036 381388 393092
rect 381444 393036 479500 393092
rect 479556 393036 479566 393092
rect 128706 392924 128716 392980
rect 128772 392924 186396 392980
rect 186452 392924 186462 392980
rect 443426 392924 443436 392980
rect 443492 392924 548268 392980
rect 548324 392924 548334 392980
rect 160962 392812 160972 392868
rect 161028 392812 237468 392868
rect 237524 392812 237534 392868
rect 442866 392812 442876 392868
rect 442932 392812 548156 392868
rect 548212 392812 548222 392868
rect 136770 392700 136780 392756
rect 136836 392700 223468 392756
rect 223524 392700 223534 392756
rect 229506 392700 229516 392756
rect 229572 392700 238588 392756
rect 238644 392700 238654 392756
rect 310930 392700 310940 392756
rect 310996 392700 326284 392756
rect 326340 392700 326350 392756
rect 334450 392700 334460 392756
rect 334516 392700 354508 392756
rect 354564 392700 354574 392756
rect 443202 392700 443212 392756
rect 443268 392700 549612 392756
rect 549668 392700 549678 392756
rect 52098 392588 52108 392644
rect 52164 392588 63868 392644
rect 63924 392588 63934 392644
rect 140802 392588 140812 392644
rect 140868 392588 228508 392644
rect 228564 392588 228574 392644
rect 237570 392588 237580 392644
rect 237636 392588 260316 392644
rect 260372 392588 260382 392644
rect 325266 392588 325276 392644
rect 325332 392588 358540 392644
rect 358596 392588 358606 392644
rect 359538 392588 359548 392644
rect 359604 392588 427084 392644
rect 427140 392588 427150 392644
rect 428418 392588 428428 392644
rect 428484 392588 544012 392644
rect 544068 392588 544078 392644
rect 30258 392476 30268 392532
rect 30324 392476 37772 392532
rect 37828 392476 37838 392532
rect 56130 392476 56140 392532
rect 56196 392476 70476 392532
rect 70532 392476 70542 392532
rect 100482 392476 100492 392532
rect 100548 392476 194908 392532
rect 194964 392476 194974 392532
rect 233538 392476 233548 392532
rect 233604 392476 263788 392532
rect 263844 392476 263854 392532
rect 314514 392476 314524 392532
rect 314580 392476 334348 392532
rect 334404 392476 334414 392532
rect 343522 392476 343532 392532
rect 343588 392476 382732 392532
rect 382788 392476 382798 392532
rect 393362 392476 393372 392532
rect 393428 392476 511756 392532
rect 511812 392476 511822 392532
rect 35970 392364 35980 392420
rect 36036 392364 57036 392420
rect 57092 392364 57102 392420
rect 60162 392364 60172 392420
rect 60228 392364 164556 392420
rect 164612 392364 164622 392420
rect 185154 392364 185164 392420
rect 185220 392364 241948 392420
rect 242004 392364 242014 392420
rect 245634 392364 245644 392420
rect 245700 392364 265468 392420
rect 265524 392364 265534 392420
rect 312722 392364 312732 392420
rect 312788 392364 330316 392420
rect 330372 392364 330382 392420
rect 334226 392364 334236 392420
rect 334292 392364 378700 392420
rect 378756 392364 378766 392420
rect 396946 392364 396956 392420
rect 397012 392364 519820 392420
rect 519876 392364 519886 392420
rect 31938 392252 31948 392308
rect 32004 392252 60396 392308
rect 60452 392252 60462 392308
rect 72258 392252 72268 392308
rect 72324 392252 188972 392308
rect 189028 392252 189038 392308
rect 189186 392252 189196 392308
rect 189252 392252 246988 392308
rect 247044 392252 247054 392308
rect 249666 392252 249676 392308
rect 249732 392252 270396 392308
rect 270452 392252 270462 392308
rect 273858 392252 273868 392308
rect 273924 392252 287644 392308
rect 287700 392252 287710 392308
rect 289986 392252 289996 392308
rect 290052 392252 294812 392308
rect 294868 392252 294878 392308
rect 318098 392252 318108 392308
rect 318164 392252 342412 392308
rect 342468 392252 342478 392308
rect 355282 392252 355292 392308
rect 355348 392252 402892 392308
rect 402948 392252 402958 392308
rect 404114 392252 404124 392308
rect 404180 392252 535948 392308
rect 536004 392252 536014 392308
rect 378690 392140 378700 392196
rect 378756 392140 475468 392196
rect 475524 392140 475534 392196
rect 164994 391580 165004 391636
rect 165060 391580 176316 391636
rect 176372 391580 176382 391636
rect 64194 391468 64204 391524
rect 64260 391468 65660 391524
rect 65716 391468 65726 391524
rect 132738 391468 132748 391524
rect 132804 391468 136108 391524
rect 136164 391468 136174 391524
rect 225474 391468 225484 391524
rect 225540 391468 231868 391524
rect 401426 391468 401436 391524
rect 401492 391468 406924 391524
rect 406980 391468 406990 391524
rect 231812 391412 231868 391468
rect 186386 391356 186396 391412
rect 186452 391356 223132 391412
rect 223188 391356 223198 391412
rect 231812 391356 243628 391412
rect 407698 391356 407708 391412
rect 407764 391356 428428 391412
rect 428484 391356 428494 391412
rect 152898 391244 152908 391300
rect 152964 391244 233884 391300
rect 233940 391244 233950 391300
rect 144834 391132 144844 391188
rect 144900 391132 230300 391188
rect 230356 391132 230366 391188
rect 112578 391020 112588 391076
rect 112644 391020 215964 391076
rect 216020 391020 216030 391076
rect 243572 390964 243628 391356
rect 348562 391244 348572 391300
rect 348628 391244 410956 391300
rect 411012 391244 411022 391300
rect 367938 391132 367948 391188
rect 368004 391132 443212 391188
rect 443268 391132 443278 391188
rect 362786 391020 362796 391076
rect 362852 391020 439180 391076
rect 439236 391020 439246 391076
rect 63858 390908 63868 390964
rect 63924 390908 187292 390964
rect 187348 390908 187358 390964
rect 243572 390908 266140 390964
rect 266196 390908 266206 390964
rect 336018 390908 336028 390964
rect 336084 390908 362572 390964
rect 362628 390908 362638 390964
rect 380818 390908 380828 390964
rect 380884 390908 483532 390964
rect 483588 390908 483598 390964
rect 57026 390796 57036 390852
rect 57092 390796 180124 390852
rect 180180 390796 180190 390852
rect 221442 390796 221452 390852
rect 221508 390796 264348 390852
rect 264404 390796 264414 390852
rect 337810 390796 337820 390852
rect 337876 390796 386764 390852
rect 386820 390796 386830 390852
rect 398738 390796 398748 390852
rect 398804 390796 523852 390852
rect 523908 390796 523918 390852
rect 4610 390684 4620 390740
rect 4676 390684 162204 390740
rect 162260 390684 162270 390740
rect 164546 390684 164556 390740
rect 164612 390684 192668 390740
rect 192724 390684 192734 390740
rect 193218 390684 193228 390740
rect 193284 390684 251804 390740
rect 251860 390684 251870 390740
rect 263778 390684 263788 390740
rect 263844 390684 269724 390740
rect 269780 390684 269790 390740
rect 301970 390684 301980 390740
rect 302036 390684 306124 390740
rect 306180 390684 306190 390740
rect 359314 390684 359324 390740
rect 359380 390684 435148 390740
rect 435204 390684 435214 390740
rect 436258 390684 436268 390740
rect 436324 390684 590716 390740
rect 590772 390684 590782 390740
rect 4274 390572 4284 390628
rect 4340 390572 165900 390628
rect 165956 390572 165966 390628
rect 169026 390572 169036 390628
rect 169092 390572 241052 390628
rect 241108 390572 241118 390628
rect 241602 390572 241612 390628
rect 241668 390572 273308 390628
rect 273364 390572 273374 390628
rect 305554 390572 305564 390628
rect 305620 390572 314188 390628
rect 314244 390572 314254 390628
rect 321682 390572 321692 390628
rect 321748 390572 350476 390628
rect 350532 390572 350542 390628
rect 351810 390572 351820 390628
rect 351876 390572 414988 390628
rect 415044 390572 415054 390628
rect 434242 390572 434252 390628
rect 434308 390572 590492 390628
rect 590548 390572 590558 390628
rect 446786 390460 446796 390516
rect 446852 390460 451276 390516
rect 451332 390460 451342 390516
rect 595560 390404 597000 390600
rect 188962 390348 188972 390404
rect 189028 390348 198044 390404
rect 198100 390348 198110 390404
rect 437714 390348 437724 390404
rect 437780 390376 597000 390404
rect 437780 390348 595672 390376
rect -960 389620 480 389816
rect 26562 389788 26572 389844
rect 26628 389788 27972 389844
rect 28466 389788 28476 389844
rect 28532 389788 31948 389844
rect 27916 389732 27972 389788
rect 31892 389732 31948 389788
rect 26674 389676 26684 389732
rect 26740 389676 27692 389732
rect 27748 389676 27758 389732
rect 27916 389676 28588 389732
rect 28644 389676 28654 389732
rect 29138 389676 29148 389732
rect 29204 389676 31052 389732
rect 31108 389676 31118 389732
rect 31892 389676 35084 389732
rect 35140 389676 35150 389732
rect 37762 389676 37772 389732
rect 37828 389676 40236 389732
rect 40292 389676 40302 389732
rect 303762 389676 303772 389732
rect 303828 389676 310156 389732
rect 310212 389676 310222 389732
rect -960 389592 169708 389620
rect 392 389564 169708 389592
rect 169764 389564 169774 389620
rect 370066 389564 370076 389620
rect 370132 389564 459340 389620
rect 459396 389564 459406 389620
rect 29026 389452 29036 389508
rect 29092 389452 35196 389508
rect 35252 389452 35262 389508
rect 371858 389452 371868 389508
rect 371924 389452 463372 389508
rect 463428 389452 463438 389508
rect 30258 389340 30268 389396
rect 30324 389340 34412 389396
rect 34468 389340 34478 389396
rect 177090 389340 177100 389396
rect 177156 389340 244636 389396
rect 244692 389340 244702 389396
rect 442642 389340 442652 389396
rect 442708 389340 549388 389396
rect 549444 389340 549454 389396
rect 120642 389228 120652 389284
rect 120708 389228 219548 389284
rect 219604 389228 219614 389284
rect 261762 389228 261772 389284
rect 261828 389228 282268 389284
rect 282324 389228 282334 389284
rect 387986 389228 387996 389284
rect 388052 389228 499660 389284
rect 499716 389228 499726 389284
rect 116610 389116 116620 389172
rect 116676 389116 217756 389172
rect 217812 389116 217822 389172
rect 253698 389116 253708 389172
rect 253764 389116 278684 389172
rect 278740 389116 278750 389172
rect 351026 389116 351036 389172
rect 351092 389116 370636 389172
rect 370692 389116 370702 389172
rect 402322 389116 402332 389172
rect 402388 389116 531916 389172
rect 531972 389116 531982 389172
rect 80322 389004 80332 389060
rect 80388 389004 201628 389060
rect 201684 389004 201694 389060
rect 238578 389004 238588 389060
rect 238644 389004 267932 389060
rect 267988 389004 267998 389060
rect 332434 389004 332444 389060
rect 332500 389004 374668 389060
rect 374724 389004 374734 389060
rect 440066 389004 440076 389060
rect 440132 389004 590716 389060
rect 590772 389004 590782 389060
rect 60386 388892 60396 388948
rect 60452 388892 189084 388948
rect 189140 388892 189150 388948
rect 197250 388892 197260 388948
rect 197316 388892 253596 388948
rect 253652 388892 253662 388948
rect 257730 388892 257740 388948
rect 257796 388892 280476 388948
rect 280532 388892 280542 388948
rect 352818 388892 352828 388948
rect 352884 388892 419020 388948
rect 419076 388892 419086 388948
rect 432674 388892 432684 388948
rect 432740 388892 587244 388948
rect 587300 388892 587310 388948
rect 340946 388220 340956 388276
rect 341012 388220 346444 388276
rect 346500 388220 346510 388276
rect 270386 387996 270396 388052
rect 270452 387996 276892 388052
rect 276948 387996 276958 388052
rect 300178 387996 300188 388052
rect 300244 387996 302092 388052
rect 302148 387996 302158 388052
rect 35074 387884 35084 387940
rect 35140 387884 41132 387940
rect 41188 387884 41198 387940
rect 173058 387884 173068 387940
rect 173124 387884 242844 387940
rect 242900 387884 242910 387940
rect 366146 387884 366156 387940
rect 366212 387884 398860 387940
rect 398916 387884 398926 387940
rect 148866 387772 148876 387828
rect 148932 387772 232092 387828
rect 232148 387772 232158 387828
rect 390562 387772 390572 387828
rect 390628 387772 431116 387828
rect 431172 387772 431182 387828
rect 88386 387660 88396 387716
rect 88452 387660 205212 387716
rect 205268 387660 205278 387716
rect 374546 387660 374556 387716
rect 374612 387660 423052 387716
rect 423108 387660 423118 387716
rect 84354 387548 84364 387604
rect 84420 387548 203420 387604
rect 203476 387548 203486 387604
rect 384402 387548 384412 387604
rect 384468 387548 491596 387604
rect 491652 387548 491662 387604
rect 70466 387436 70476 387492
rect 70532 387436 190876 387492
rect 190932 387436 190942 387492
rect 217410 387436 217420 387492
rect 217476 387436 262556 387492
rect 262612 387436 262622 387492
rect 328850 387436 328860 387492
rect 328916 387436 366604 387492
rect 366660 387436 366670 387492
rect 391570 387436 391580 387492
rect 391636 387436 507724 387492
rect 507780 387436 507790 387492
rect 44034 387324 44044 387380
rect 44100 387324 183708 387380
rect 183764 387324 183774 387380
rect 201282 387324 201292 387380
rect 201348 387324 255388 387380
rect 255444 387324 255454 387380
rect 323474 387324 323484 387380
rect 323540 387324 334460 387380
rect 334516 387324 334526 387380
rect 344530 387324 344540 387380
rect 344596 387324 390796 387380
rect 390852 387324 390862 387380
rect 395154 387324 395164 387380
rect 395220 387324 515788 387380
rect 515844 387324 515854 387380
rect 40002 387212 40012 387268
rect 40068 387212 181916 387268
rect 181972 387212 181982 387268
rect 184772 387212 246428 387268
rect 246484 387212 246494 387268
rect 265458 387212 265468 387268
rect 265524 387212 275100 387268
rect 275156 387212 275166 387268
rect 281922 387212 281932 387268
rect 281988 387212 291228 387268
rect 291284 387212 291294 387268
rect 316306 387212 316316 387268
rect 316372 387212 338380 387268
rect 338436 387212 338446 387268
rect 341394 387212 341404 387268
rect 341460 387212 394828 387268
rect 394884 387212 394894 387268
rect 405906 387212 405916 387268
rect 405972 387212 539980 387268
rect 540036 387212 540046 387268
rect 184772 387156 184828 387212
rect 181458 387100 181468 387156
rect 181524 387100 184828 387156
rect 285954 386428 285964 386484
rect 286020 386428 293020 386484
rect 293076 386428 293086 386484
rect 35186 386316 35196 386372
rect 35252 386316 39004 386372
rect 39060 386316 39070 386372
rect 194898 386316 194908 386372
rect 194964 386316 210588 386372
rect 210644 386316 210654 386372
rect 223458 386316 223468 386372
rect 223524 386316 226716 386372
rect 226772 386316 226782 386372
rect 246978 386316 246988 386372
rect 247044 386316 250012 386372
rect 250068 386316 250078 386372
rect 294018 386316 294028 386372
rect 294084 386316 296604 386372
rect 296660 386316 296670 386372
rect 327058 386316 327068 386372
rect 327124 386316 336028 386372
rect 336084 386316 336094 386372
rect 350354 386316 350364 386372
rect 350420 386316 351820 386372
rect 351876 386316 351886 386372
rect 355730 386316 355740 386372
rect 355796 386316 359548 386372
rect 359604 386316 359614 386372
rect 366482 386316 366492 386372
rect 366548 386316 446796 386372
rect 446852 386316 446862 386372
rect 176306 386204 176316 386260
rect 176372 386204 239260 386260
rect 239316 386204 239326 386260
rect 362898 386204 362908 386260
rect 362964 386204 367948 386260
rect 368004 386204 368014 386260
rect 368274 386204 368284 386260
rect 368340 386204 455308 386260
rect 455364 386204 455374 386260
rect 136098 386092 136108 386148
rect 136164 386092 224924 386148
rect 224980 386092 224990 386148
rect 377234 386092 377244 386148
rect 377300 386092 378700 386148
rect 378756 386092 378766 386148
rect 379026 386092 379036 386148
rect 379092 386092 381388 386148
rect 381444 386092 381454 386148
rect 443202 386092 443212 386148
rect 443268 386092 547708 386148
rect 547764 386092 547774 386148
rect 108546 385980 108556 386036
rect 108612 385980 214172 386036
rect 214228 385980 214238 386036
rect 339602 385980 339612 386036
rect 339668 385980 344540 386036
rect 344596 385980 344606 386036
rect 344978 385980 344988 386036
rect 345044 385980 355292 386036
rect 355348 385980 355358 386036
rect 382610 385980 382620 386036
rect 382676 385980 487564 386036
rect 487620 385980 487630 386036
rect 104514 385868 104524 385924
rect 104580 385868 212380 385924
rect 212436 385868 212446 385924
rect 241938 385868 241948 385924
rect 242004 385868 248220 385924
rect 248276 385868 248286 385924
rect 260306 385868 260316 385924
rect 260372 385868 271516 385924
rect 271572 385868 271582 385924
rect 336018 385868 336028 385924
rect 336084 385868 343532 385924
rect 343588 385868 343598 385924
rect 353938 385868 353948 385924
rect 354004 385868 374556 385924
rect 374612 385868 374622 385924
rect 386194 385868 386204 385924
rect 386260 385868 495628 385924
rect 495684 385868 495694 385924
rect 76290 385756 76300 385812
rect 76356 385756 199836 385812
rect 199892 385756 199902 385812
rect 213378 385756 213388 385812
rect 213444 385756 260764 385812
rect 260820 385756 260830 385812
rect 277890 385756 277900 385812
rect 277956 385756 289436 385812
rect 289492 385756 289502 385812
rect 343186 385756 343196 385812
rect 343252 385756 366156 385812
rect 366212 385756 366222 385812
rect 389778 385756 389788 385812
rect 389844 385756 503692 385812
rect 503748 385756 503758 385812
rect 68226 385644 68236 385700
rect 68292 385644 196252 385700
rect 196308 385644 196318 385700
rect 210018 385644 210028 385700
rect 210084 385644 258972 385700
rect 259028 385644 259038 385700
rect 269826 385644 269836 385700
rect 269892 385644 285852 385700
rect 285908 385644 285918 385700
rect 309138 385644 309148 385700
rect 309204 385644 322252 385700
rect 322308 385644 322318 385700
rect 330642 385644 330652 385700
rect 330708 385644 351036 385700
rect 351092 385644 351102 385700
rect 357522 385644 357532 385700
rect 357588 385644 390572 385700
rect 390628 385644 390638 385700
rect 400530 385644 400540 385700
rect 400596 385644 527884 385700
rect 527940 385644 527950 385700
rect 40338 385532 40348 385588
rect 40404 385532 47852 385588
rect 47908 385532 47918 385588
rect 65650 385532 65660 385588
rect 65716 385532 194460 385588
rect 194516 385532 194526 385588
rect 205314 385532 205324 385588
rect 205380 385532 257180 385588
rect 257236 385532 257246 385588
rect 265794 385532 265804 385588
rect 265860 385532 284060 385588
rect 284116 385532 284126 385588
rect 307346 385532 307356 385588
rect 307412 385532 318220 385588
rect 318276 385532 318286 385588
rect 319890 385532 319900 385588
rect 319956 385532 340956 385588
rect 341012 385532 341022 385588
rect 346770 385532 346780 385588
rect 346836 385532 401436 385588
rect 401492 385532 401502 385588
rect 432562 385532 432572 385588
rect 432628 385532 587132 385588
rect 587188 385532 587198 385588
rect 28578 384748 28588 384804
rect 28644 384748 30324 384804
rect 361106 384748 361116 384804
rect 361172 384748 362796 384804
rect 362852 384748 362862 384804
rect 30268 384692 30324 384748
rect 30268 384636 33404 384692
rect 33460 384636 33470 384692
rect 124674 384300 124684 384356
rect 124740 384300 221340 384356
rect 221396 384300 221406 384356
rect 92418 384188 92428 384244
rect 92484 384188 207004 384244
rect 207060 384188 207070 384244
rect 364690 384188 364700 384244
rect 364756 384188 447244 384244
rect 447300 384188 447310 384244
rect 31042 384076 31052 384132
rect 31108 384076 36764 384132
rect 36820 384076 36830 384132
rect 48066 384076 48076 384132
rect 48132 384076 185500 384132
rect 185556 384076 185566 384132
rect 373650 384076 373660 384132
rect 373716 384076 467404 384132
rect 467460 384076 467470 384132
rect 4722 383964 4732 384020
rect 4788 383964 152124 384020
rect 152180 383964 152190 384020
rect 375442 383964 375452 384020
rect 375508 383964 471436 384020
rect 471492 383964 471502 384020
rect 4498 383852 4508 383908
rect 4564 383852 165788 383908
rect 165844 383852 165854 383908
rect 430882 383852 430892 383908
rect 430948 383852 591164 383908
rect 591220 383852 591230 383908
rect 29250 382956 29260 383012
rect 29316 382956 33516 383012
rect 33572 382956 33582 383012
rect 41122 382172 41132 382228
rect 41188 382172 48636 382228
rect 48692 382172 48702 382228
rect 33394 381836 33404 381892
rect 33460 381836 37772 381892
rect 37828 381836 37838 381892
rect 34402 381388 34412 381444
rect 34468 381388 36876 381444
rect 36932 381388 36942 381444
rect 38994 381388 39004 381444
rect 39060 381388 42812 381444
rect 42868 381388 42878 381444
rect 48626 381276 48636 381332
rect 48692 381276 50428 381332
rect 50484 381276 50494 381332
rect 434466 380604 434476 380660
rect 434532 380604 562604 380660
rect 562660 380604 562670 380660
rect 19170 380492 19180 380548
rect 19236 380492 163772 380548
rect 163828 380492 163838 380548
rect 429202 380492 429212 380548
rect 429268 380492 590940 380548
rect 590996 380492 591006 380548
rect 33506 379708 33516 379764
rect 33572 379708 37044 379764
rect 36988 379652 37044 379708
rect 36988 379596 43708 379652
rect 36866 379484 36876 379540
rect 36932 379484 42028 379540
rect 42084 379484 42094 379540
rect 43652 379316 43708 379596
rect 43652 379260 46956 379316
rect 47012 379260 47022 379316
rect 27906 378924 27916 378980
rect 27972 378924 172172 378980
rect 172228 378924 172238 378980
rect 10994 378812 11004 378868
rect 11060 378812 166348 378868
rect 166404 378812 166414 378868
rect 425842 378812 425852 378868
rect 425908 378812 584668 378868
rect 584724 378812 584734 378868
rect 50418 378028 50428 378084
rect 50484 378028 52164 378084
rect 52108 377972 52164 378028
rect 27682 377916 27692 377972
rect 27748 377916 28700 377972
rect 28756 377916 28766 377972
rect 52108 377916 57036 377972
rect 57092 377916 57102 377972
rect 28242 377356 28252 377412
rect 28308 377356 36876 377412
rect 36932 377356 36942 377412
rect 42018 377356 42028 377412
rect 42084 377356 48636 377412
rect 48692 377356 48702 377412
rect 12562 377244 12572 377300
rect 12628 377244 163996 377300
rect 164052 377244 164062 377300
rect 595560 377188 597000 377384
rect 4946 377132 4956 377188
rect 5012 377132 166012 377188
rect 166068 377132 166078 377188
rect 424162 377132 424172 377188
rect 424228 377160 597000 377188
rect 424228 377132 595672 377160
rect 46946 376236 46956 376292
rect 47012 376236 50428 376292
rect 50484 376236 50494 376292
rect 47842 376124 47852 376180
rect 47908 376124 62188 376180
rect 62244 376124 62254 376180
rect 57026 376012 57036 376068
rect 57092 376012 154588 376068
rect 154644 376012 154654 376068
rect 36866 375900 36876 375956
rect 36932 375900 151004 375956
rect 151060 375900 151070 375956
rect 37762 375788 37772 375844
rect 37828 375788 152908 375844
rect 152964 375788 152974 375844
rect -960 375508 480 375704
rect 28690 375676 28700 375732
rect 28756 375676 154252 375732
rect 154308 375676 154318 375732
rect 29474 375564 29484 375620
rect 29540 375564 163996 375620
rect 164052 375564 164062 375620
rect -960 375480 152236 375508
rect 392 375452 152236 375480
rect 152292 375452 152302 375508
rect 165442 375452 165452 375508
rect 165508 375452 174104 375508
rect 413756 375284 413812 375480
rect 434242 375452 434252 375508
rect 434308 375452 590604 375508
rect 590660 375452 590670 375508
rect 419972 375340 441196 375396
rect 441252 375340 441262 375396
rect 419972 375284 420028 375340
rect 413756 375228 420028 375284
rect 153794 374780 153804 374836
rect 153860 374780 174104 374836
rect 413896 374780 420924 374836
rect 420980 374780 420990 374836
rect 29362 374556 29372 374612
rect 29428 374556 164556 374612
rect 164612 374556 164622 374612
rect 544226 374556 544236 374612
rect 544292 374556 547932 374612
rect 547988 374556 547998 374612
rect 62178 374444 62188 374500
rect 62244 374444 151116 374500
rect 151172 374444 151182 374500
rect 154578 374444 154588 374500
rect 154644 374444 157948 374500
rect 158004 374444 158014 374500
rect 48626 374332 48636 374388
rect 48692 374332 149324 374388
rect 149380 374332 149390 374388
rect 150994 374332 151004 374388
rect 151060 374332 154364 374388
rect 154420 374332 154430 374388
rect 36978 374220 36988 374276
rect 37044 374220 156156 374276
rect 156212 374220 156222 374276
rect 160738 374108 160748 374164
rect 160804 374108 174104 374164
rect 413896 374108 422604 374164
rect 422660 374108 422670 374164
rect 28354 373996 28364 374052
rect 28420 373996 164332 374052
rect 164388 373996 164398 374052
rect 26786 373884 26796 373940
rect 26852 373884 164108 373940
rect 164164 373884 164174 373940
rect 535042 373884 535052 373940
rect 535108 373884 549500 373940
rect 549556 373884 549566 373940
rect 14242 373772 14252 373828
rect 14308 373772 163884 373828
rect 163940 373772 163950 373828
rect 425842 373772 425852 373828
rect 425908 373772 590380 373828
rect 590436 373772 590446 373828
rect 160514 373436 160524 373492
rect 160580 373436 174104 373492
rect 413896 373436 417564 373492
rect 417620 373436 417630 373492
rect 442754 373212 442764 373268
rect 442820 373212 591052 373268
rect 591108 373212 591118 373268
rect 437938 373100 437948 373156
rect 438004 373100 590604 373156
rect 590660 373100 590670 373156
rect 50418 372988 50428 373044
rect 50484 372988 58828 373044
rect 152898 372988 152908 373044
rect 152964 372988 156324 373044
rect 435922 372988 435932 373044
rect 435988 372988 590828 373044
rect 590884 372988 590894 373044
rect 58772 372820 58828 372988
rect 156268 372932 156324 372988
rect 156268 372876 159516 372932
rect 159572 372876 159582 372932
rect 58772 372764 67228 372820
rect 153682 372764 153692 372820
rect 153748 372764 174104 372820
rect 413896 372764 432908 372820
rect 432964 372764 432974 372820
rect 67172 372596 67228 372764
rect 67172 372540 151116 372596
rect 151172 372540 151182 372596
rect 42802 372428 42812 372484
rect 42868 372428 152796 372484
rect 152852 372428 152862 372484
rect 440178 372428 440188 372484
rect 440244 372428 535052 372484
rect 535108 372428 535118 372484
rect 28466 372316 28476 372372
rect 28532 372316 164220 372372
rect 164276 372316 164286 372372
rect 436034 372316 436044 372372
rect 436100 372316 544236 372372
rect 544292 372316 544302 372372
rect 4946 372204 4956 372260
rect 5012 372204 150780 372260
rect 150836 372204 150846 372260
rect 437602 372204 437612 372260
rect 437668 372204 547820 372260
rect 547876 372204 547886 372260
rect 17602 372092 17612 372148
rect 17668 372092 163772 372148
rect 163828 372092 163838 372148
rect 168802 372092 168812 372148
rect 168868 372092 174104 372148
rect 413896 372092 417676 372148
rect 417732 372092 417742 372148
rect 424386 372092 424396 372148
rect 424452 372092 590492 372148
rect 590548 372092 590558 372148
rect 4274 371420 4284 371476
rect 4340 371420 150332 371476
rect 150388 371420 150398 371476
rect 157154 371420 157164 371476
rect 157220 371420 174104 371476
rect 413896 371420 417900 371476
rect 417956 371420 417966 371476
rect 442866 371420 442876 371476
rect 442932 371420 590716 371476
rect 590772 371420 590782 371476
rect 4162 371308 4172 371364
rect 4228 371308 150556 371364
rect 150612 371308 150622 371364
rect 157938 371308 157948 371364
rect 158004 371308 161308 371364
rect 443090 371308 443100 371364
rect 443156 371308 590940 371364
rect 590996 371308 591006 371364
rect 161252 371140 161308 371308
rect 161252 371084 162876 371140
rect 162932 371084 162942 371140
rect 160402 370748 160412 370804
rect 160468 370748 174104 370804
rect 413896 370748 421036 370804
rect 421092 370748 421102 370804
rect 149538 370636 149548 370692
rect 149604 370636 151452 370692
rect 151508 370636 151518 370692
rect 442978 370636 442988 370692
rect 443044 370636 590492 370692
rect 590548 370636 590558 370692
rect 169810 370076 169820 370132
rect 169876 370076 174104 370132
rect 413896 370076 425964 370132
rect 426020 370076 426030 370132
rect 151218 369628 151228 369684
rect 151284 369628 153020 369684
rect 153076 369628 153086 369684
rect 156370 369628 156380 369684
rect 156436 369628 158452 369684
rect 158396 369572 158452 369628
rect 158396 369516 160524 369572
rect 160580 369516 160590 369572
rect 155026 369404 155036 369460
rect 155092 369404 174104 369460
rect 413896 369404 427980 369460
rect 428036 369404 428046 369460
rect 154802 369180 154812 369236
rect 154868 369180 159516 369236
rect 159572 369180 159582 369236
rect 159618 368844 159628 368900
rect 159684 368844 166796 368900
rect 166852 368844 166862 368900
rect 426738 368844 426748 368900
rect 426804 368844 437612 368900
rect 437668 368844 437678 368900
rect 155586 368732 155596 368788
rect 155652 368732 174104 368788
rect 413896 368732 418348 368788
rect 418404 368732 418414 368788
rect 427522 368732 427532 368788
rect 427588 368732 440188 368788
rect 440244 368732 440254 368788
rect 155362 368060 155372 368116
rect 155428 368060 174104 368116
rect 413896 368060 440972 368116
rect 441028 368060 441038 368116
rect 151442 367948 151452 368004
rect 151508 367948 154532 368004
rect 154690 367948 154700 368004
rect 154756 367948 157052 368004
rect 157108 367948 157118 368004
rect 154476 367892 154532 367948
rect 154476 367836 160412 367892
rect 160468 367836 160478 367892
rect 156818 367388 156828 367444
rect 156884 367388 174104 367444
rect 413896 367388 429436 367444
rect 429492 367388 429502 367444
rect 157042 367052 157052 367108
rect 157108 367052 169820 367108
rect 169876 367052 169886 367108
rect 155138 366716 155148 366772
rect 155204 366716 174104 366772
rect 413896 366716 432796 366772
rect 432852 366716 432862 366772
rect 166786 366156 166796 366212
rect 166852 366156 172396 366212
rect 172452 366156 172462 366212
rect 157826 366044 157836 366100
rect 157892 366044 174104 366100
rect 413896 366044 419020 366100
rect 419076 366044 419086 366100
rect 418338 365484 418348 365540
rect 418404 365484 441084 365540
rect 441140 365484 441150 365540
rect 159618 365372 159628 365428
rect 159684 365372 167244 365428
rect 167300 365372 167310 365428
rect 170818 365372 170828 365428
rect 170884 365372 174104 365428
rect 413896 365372 419916 365428
rect 419972 365372 419982 365428
rect 153906 364700 153916 364756
rect 153972 364700 174104 364756
rect 413896 364700 416108 364756
rect 416164 364700 416174 364756
rect 151218 364476 151228 364532
rect 151284 364476 154476 364532
rect 154532 364476 154542 364532
rect 162866 364476 162876 364532
rect 162932 364476 167580 364532
rect 167636 364476 167646 364532
rect 152898 364364 152908 364420
rect 152964 364364 154588 364420
rect 154644 364364 154654 364420
rect 591042 364140 591052 364196
rect 591108 364168 595672 364196
rect 591108 364140 597000 364168
rect 169810 364028 169820 364084
rect 169876 364028 174104 364084
rect 413896 364028 420812 364084
rect 420868 364028 420878 364084
rect 595560 363944 597000 364140
rect 170482 363356 170492 363412
rect 170548 363356 174104 363412
rect 413896 363356 437388 363412
rect 437444 363356 437454 363412
rect 153010 363020 153020 363076
rect 153076 363020 162092 363076
rect 162148 363020 162158 363076
rect 154354 362796 154364 362852
rect 154420 362796 160748 362852
rect 160804 362796 160814 362852
rect 420914 362796 420924 362852
rect 420980 362796 426748 362852
rect 426804 362796 426814 362852
rect 154578 362684 154588 362740
rect 154644 362684 158060 362740
rect 158116 362684 158126 362740
rect 172610 362684 172620 362740
rect 172676 362684 174104 362740
rect 413896 362684 438396 362740
rect 438452 362684 438462 362740
rect 160290 362124 160300 362180
rect 160356 362124 169820 362180
rect 169876 362124 169886 362180
rect 167458 362012 167468 362068
rect 167524 362012 174104 362068
rect 413896 362012 422492 362068
rect 422548 362012 422558 362068
rect 149912 361676 165452 361732
rect 165508 361676 165518 361732
rect 441186 361676 441196 361732
rect 441252 361676 444136 361732
rect 392 361592 4172 361620
rect -960 361564 4172 361592
rect 4228 361564 4238 361620
rect -960 361368 480 361564
rect 161186 361340 161196 361396
rect 161252 361340 174104 361396
rect 413896 361340 420700 361396
rect 420756 361340 420766 361396
rect 170258 360668 170268 360724
rect 170324 360668 174104 360724
rect 413896 360668 419804 360724
rect 419860 360668 419870 360724
rect 156930 360332 156940 360388
rect 156996 360332 170828 360388
rect 170884 360332 170894 360388
rect 421026 360332 421036 360388
rect 421092 360332 441196 360388
rect 441252 360332 441262 360388
rect 169250 359996 169260 360052
rect 169316 359996 174104 360052
rect 413896 359996 434924 360052
rect 434980 359996 434990 360052
rect 167234 359548 167244 359604
rect 167300 359548 168084 359604
rect 168028 359492 168084 359548
rect 168028 359436 171388 359492
rect 171444 359436 171454 359492
rect 166114 359324 166124 359380
rect 166180 359324 174104 359380
rect 413896 359324 417452 359380
rect 417508 359324 417518 359380
rect 158050 358764 158060 358820
rect 158116 358764 162204 358820
rect 162260 358764 162270 358820
rect 157714 358652 157724 358708
rect 157780 358652 174104 358708
rect 413896 358652 442540 358708
rect 442596 358652 442606 358708
rect 149912 358092 153804 358148
rect 153860 358092 153870 358148
rect 420914 358092 420924 358148
rect 420980 358092 444136 358148
rect 154466 357868 154476 357924
rect 154532 357868 160524 357924
rect 160580 357868 160590 357924
rect 174076 357588 174132 358008
rect 413896 357980 419692 358036
rect 419748 357980 419758 358036
rect 173170 357532 173180 357588
rect 173236 357532 174132 357588
rect 171042 357308 171052 357364
rect 171108 357308 174104 357364
rect 413896 357308 431228 357364
rect 431284 357308 431294 357364
rect 422594 356972 422604 357028
rect 422660 356972 440188 357028
rect 440244 356972 440254 357028
rect 169362 356636 169372 356692
rect 169428 356636 174104 356692
rect 413896 356636 417788 356692
rect 417844 356636 417854 356692
rect 158498 355964 158508 356020
rect 158564 355964 174104 356020
rect 413896 355964 421596 356020
rect 421652 355964 421662 356020
rect 169810 355292 169820 355348
rect 169876 355292 174104 355348
rect 413896 355292 436604 355348
rect 436660 355292 436670 355348
rect 167570 355068 167580 355124
rect 167636 355068 170268 355124
rect 170324 355068 170334 355124
rect 172498 354620 172508 354676
rect 172564 354620 174104 354676
rect 413896 354620 433244 354676
rect 433300 354620 433310 354676
rect 149912 354508 154364 354564
rect 154420 354508 154430 354564
rect 154690 354508 154700 354564
rect 154756 354508 156324 354564
rect 440178 354508 440188 354564
rect 440244 354508 444136 354564
rect 156268 354452 156324 354508
rect 156268 354396 158844 354452
rect 158900 354396 158910 354452
rect 167570 354396 167580 354452
rect 167636 354396 170492 354452
rect 170548 354396 170558 354452
rect 156146 353948 156156 354004
rect 156212 353948 174104 354004
rect 413896 353948 415772 354004
rect 415828 353948 415838 354004
rect 150882 353612 150892 353668
rect 150948 353612 169820 353668
rect 169876 353612 169886 353668
rect 417666 353612 417676 353668
rect 417732 353612 441308 353668
rect 441364 353612 441374 353668
rect 158610 353276 158620 353332
rect 158676 353276 174104 353332
rect 413896 353276 418012 353332
rect 418068 353276 418078 353332
rect 157042 352716 157052 352772
rect 157108 352716 160860 352772
rect 160916 352716 160926 352772
rect 171266 352604 171276 352660
rect 171332 352604 174104 352660
rect 413896 352604 429212 352660
rect 429268 352604 429278 352660
rect 170818 351932 170828 351988
rect 170884 351932 174104 351988
rect 413896 351932 427868 351988
rect 427924 351932 427934 351988
rect 173012 351260 174104 351316
rect 413896 351260 420924 351316
rect 420980 351260 420990 351316
rect 173012 351204 173068 351260
rect 169708 351148 173068 351204
rect 169708 351092 169764 351148
rect 162530 351036 162540 351092
rect 162596 351036 169764 351092
rect 149912 350924 154476 350980
rect 154532 350924 154542 350980
rect 417554 350924 417564 350980
rect 417620 350924 444136 350980
rect 590818 350924 590828 350980
rect 590884 350952 595672 350980
rect 590884 350924 597000 350952
rect 595560 350728 597000 350924
rect 170930 350588 170940 350644
rect 170996 350588 174104 350644
rect 413896 350588 418236 350644
rect 418292 350588 418302 350644
rect 169138 349916 169148 349972
rect 169204 349916 174104 349972
rect 413896 349916 438956 349972
rect 439012 349916 439022 349972
rect 171378 349468 171388 349524
rect 171444 349468 173852 349524
rect 173908 349468 173918 349524
rect 169026 349244 169036 349300
rect 169092 349244 174104 349300
rect 413896 349244 426412 349300
rect 426468 349244 426478 349300
rect 160850 348684 160860 348740
rect 160916 348684 167132 348740
rect 167188 348684 167198 348740
rect 417890 348684 417900 348740
rect 417956 348684 440188 348740
rect 440244 348684 440254 348740
rect 154354 348572 154364 348628
rect 154420 348572 174104 348628
rect 413896 348572 417564 348628
rect 417620 348572 417630 348628
rect 418226 348572 418236 348628
rect 418292 348572 443324 348628
rect 443380 348572 443390 348628
rect 165666 347900 165676 347956
rect 165732 347900 174104 347956
rect 413896 347900 416668 347956
rect 416724 347900 416734 347956
rect 158834 347788 158844 347844
rect 158900 347788 161308 347844
rect 161252 347732 161308 347788
rect 161252 347676 162316 347732
rect 162372 347676 162382 347732
rect 392 347480 4172 347508
rect -960 347452 4172 347480
rect 4228 347452 4238 347508
rect -960 347256 480 347452
rect 149912 347340 153692 347396
rect 153748 347340 153758 347396
rect 432898 347340 432908 347396
rect 432964 347340 444136 347396
rect 173730 347228 173740 347284
rect 173796 347228 174104 347284
rect 413896 347228 416780 347284
rect 416836 347228 416846 347284
rect 416658 346892 416668 346948
rect 416724 346892 433132 346948
rect 433188 346892 433198 346948
rect 174066 346556 174076 346612
rect 174132 346556 174142 346612
rect 413896 346556 426300 346612
rect 426356 346556 426366 346612
rect 167122 346108 167132 346164
rect 167188 346108 169876 346164
rect 169820 345828 169876 346108
rect 170594 345884 170604 345940
rect 170660 345884 174104 345940
rect 413896 345884 417676 345940
rect 417732 345884 417742 345940
rect 169820 345772 173068 345828
rect 173012 345716 173068 345772
rect 173012 345660 173964 345716
rect 174020 345660 174030 345716
rect 418002 345324 418012 345380
rect 418068 345324 429324 345380
rect 429380 345324 429390 345380
rect 161074 345212 161084 345268
rect 161140 345212 174104 345268
rect 413896 345212 418236 345268
rect 418292 345212 418302 345268
rect 172386 344540 172396 344596
rect 172452 344540 174104 344596
rect 413896 344540 424396 344596
rect 424452 344540 424462 344596
rect 156034 343868 156044 343924
rect 156100 343868 174104 343924
rect 413896 343868 427756 343924
rect 427812 343868 427822 343924
rect 149912 343756 168812 343812
rect 168868 343756 168878 343812
rect 441298 343756 441308 343812
rect 441364 343756 444136 343812
rect 416770 343532 416780 343588
rect 416836 343532 438172 343588
rect 438228 343532 438238 343588
rect 154242 343196 154252 343252
rect 154308 343196 174104 343252
rect 413896 343196 423276 343252
rect 423332 343196 423342 343252
rect 170706 342524 170716 342580
rect 170772 342524 174104 342580
rect 413896 342524 434812 342580
rect 434868 342524 434878 342580
rect 150994 341852 151004 341908
rect 151060 341852 174104 341908
rect 413896 341852 416668 341908
rect 416724 341852 416734 341908
rect 425954 341852 425964 341908
rect 426020 341852 441644 341908
rect 441700 341852 441710 341908
rect 155922 341180 155932 341236
rect 155988 341180 174104 341236
rect 413896 341180 424284 341236
rect 424340 341180 424350 341236
rect 424946 340956 424956 341012
rect 425012 340956 427532 341012
rect 427588 340956 427598 341012
rect 165554 340508 165564 340564
rect 165620 340508 174104 340564
rect 413896 340508 423164 340564
rect 423220 340508 423230 340564
rect 152338 340284 152348 340340
rect 152404 340284 170940 340340
rect 170996 340284 171006 340340
rect 427970 340284 427980 340340
rect 428036 340284 440300 340340
rect 440356 340284 440366 340340
rect 149912 340172 157164 340228
rect 157220 340172 157230 340228
rect 416658 340172 416668 340228
rect 416724 340172 439068 340228
rect 439124 340172 439134 340228
rect 440178 340172 440188 340228
rect 440244 340172 444136 340228
rect 160850 339836 160860 339892
rect 160916 339836 174104 339892
rect 413896 339836 415996 339892
rect 416052 339836 416062 339892
rect 157602 339164 157612 339220
rect 157668 339164 174104 339220
rect 413896 339164 426188 339220
rect 426244 339164 426254 339220
rect 429314 338604 429324 338660
rect 429380 338604 436044 338660
rect 436100 338604 436110 338660
rect 155810 338492 155820 338548
rect 155876 338492 174104 338548
rect 413896 338492 433020 338548
rect 433076 338492 433086 338548
rect 154130 337820 154140 337876
rect 154196 337820 174104 337876
rect 413896 337820 423052 337876
rect 423108 337820 423118 337876
rect 414082 337708 414092 337764
rect 414148 337708 420924 337764
rect 420980 337708 420990 337764
rect 595560 337652 597000 337736
rect 590594 337596 590604 337652
rect 590660 337596 597000 337652
rect 595560 337512 597000 337596
rect 174066 337148 174076 337204
rect 174132 337148 174142 337204
rect 413896 337148 421484 337204
rect 421540 337148 421550 337204
rect 420914 336812 420924 336868
rect 420980 336812 441532 336868
rect 441588 336812 441598 336868
rect 149912 336588 160412 336644
rect 160468 336588 160478 336644
rect 441186 336588 441196 336644
rect 441252 336588 444136 336644
rect 157490 336476 157500 336532
rect 157556 336476 174104 336532
rect 413896 336476 432908 336532
rect 432964 336476 432974 336532
rect 169810 335804 169820 335860
rect 169876 335804 174104 335860
rect 413896 335804 431004 335860
rect 431060 335804 431070 335860
rect 167346 335132 167356 335188
rect 167412 335132 174104 335188
rect 413896 335132 438284 335188
rect 438340 335132 438350 335188
rect 160738 334460 160748 334516
rect 160804 334460 174104 334516
rect 413896 334460 421372 334516
rect 421428 334460 421438 334516
rect 164210 334348 164220 334404
rect 164276 334348 170492 334404
rect 170548 334348 170558 334404
rect 432786 334348 432796 334404
rect 432852 334348 441308 334404
rect 441364 334348 441374 334404
rect 157378 333788 157388 333844
rect 157444 333788 174104 333844
rect 413896 333788 419468 333844
rect 419524 333788 419534 333844
rect 419122 333452 419132 333508
rect 419188 333452 424956 333508
rect 425012 333452 425022 333508
rect -960 333172 480 333368
rect -960 333144 7532 333172
rect 392 333116 7532 333144
rect 7588 333116 7598 333172
rect 170482 333116 170492 333172
rect 170548 333116 174104 333172
rect 413896 333116 434700 333172
rect 434756 333116 434766 333172
rect 149912 333004 157052 333060
rect 157108 333004 157118 333060
rect 441634 333004 441644 333060
rect 441700 333004 444136 333060
rect 154018 332444 154028 332500
rect 154084 332444 174104 332500
rect 413896 332444 422940 332500
rect 422996 332444 423006 332500
rect 420802 331884 420812 331940
rect 420868 331884 440748 331940
rect 440804 331884 440814 331940
rect 158834 331772 158844 331828
rect 158900 331772 174104 331828
rect 413896 331772 421260 331828
rect 421316 331772 421326 331828
rect 157266 331100 157276 331156
rect 157332 331100 174104 331156
rect 413896 331100 434588 331156
rect 434644 331100 434654 331156
rect 167234 330428 167244 330484
rect 167300 330428 174104 330484
rect 413896 330428 436492 330484
rect 436548 330428 436558 330484
rect 155698 330092 155708 330148
rect 155764 330092 169820 330148
rect 169876 330092 169886 330148
rect 422482 330092 422492 330148
rect 422548 330092 440860 330148
rect 440916 330092 440926 330148
rect 168914 329756 168924 329812
rect 168980 329756 174104 329812
rect 413896 329756 422716 329812
rect 422772 329756 422782 329812
rect 149912 329420 155036 329476
rect 155092 329420 155102 329476
rect 440178 329420 440188 329476
rect 440244 329420 444136 329476
rect 164098 329196 164108 329252
rect 164164 329196 170716 329252
rect 170772 329196 170782 329252
rect 160626 329084 160636 329140
rect 160692 329084 174104 329140
rect 413896 329084 424508 329140
rect 424564 329084 424574 329140
rect 169810 328412 169820 328468
rect 169876 328412 174104 328468
rect 413896 328412 419356 328468
rect 419412 328412 419422 328468
rect 174076 327348 174132 327768
rect 413896 327740 427644 327796
rect 427700 327740 427710 327796
rect 173058 327292 173068 327348
rect 173124 327292 174132 327348
rect 162418 327068 162428 327124
rect 162484 327068 174104 327124
rect 413896 327068 422604 327124
rect 422660 327068 422670 327124
rect 153794 326396 153804 326452
rect 153860 326396 174104 326452
rect 413896 326396 422828 326452
rect 422884 326396 422894 326452
rect 149912 325836 155596 325892
rect 155652 325836 155662 325892
rect 441074 325836 441084 325892
rect 441140 325836 444136 325892
rect 151106 325724 151116 325780
rect 151172 325724 174104 325780
rect 413896 325724 421036 325780
rect 421092 325724 421102 325780
rect 157154 325276 157164 325332
rect 157220 325276 169820 325332
rect 169876 325276 169886 325332
rect 169810 325052 169820 325108
rect 169876 325052 174104 325108
rect 413896 325052 419244 325108
rect 419300 325052 419310 325108
rect 170482 324604 170492 324660
rect 170548 324604 173964 324660
rect 174020 324604 174030 324660
rect 590930 324492 590940 324548
rect 590996 324520 595672 324548
rect 590996 324492 597000 324520
rect 172274 324380 172284 324436
rect 172340 324380 174104 324436
rect 413896 324380 425964 324436
rect 426020 324380 426030 324436
rect 425058 324268 425068 324324
rect 425124 324268 429324 324324
rect 429380 324268 429390 324324
rect 595560 324296 597000 324492
rect 153682 323708 153692 323764
rect 153748 323708 174104 323764
rect 413896 323708 416668 323764
rect 416724 323708 416734 323764
rect 418226 323484 418236 323540
rect 418292 323484 431116 323540
rect 431172 323484 431182 323540
rect 417778 323372 417788 323428
rect 417844 323372 441196 323428
rect 441252 323372 441262 323428
rect 160402 323036 160412 323092
rect 160468 323036 174104 323092
rect 413896 323036 418012 323092
rect 418068 323036 418078 323092
rect 158722 322364 158732 322420
rect 158788 322364 174104 322420
rect 413896 322364 419580 322420
rect 419636 322364 419646 322420
rect 149912 322252 155372 322308
rect 155428 322252 155438 322308
rect 440962 322252 440972 322308
rect 441028 322252 444136 322308
rect 169922 321692 169932 321748
rect 169988 321692 174104 321748
rect 413896 321692 419132 321748
rect 419188 321692 419198 321748
rect 172162 321020 172172 321076
rect 172228 321020 174104 321076
rect 413896 321020 417788 321076
rect 417844 321020 417854 321076
rect 423266 320908 423276 320964
rect 423332 320908 425068 320964
rect 425124 320908 425134 320964
rect 165442 320348 165452 320404
rect 165508 320348 174104 320404
rect 413896 320348 422492 320404
rect 422548 320348 422558 320404
rect 429426 320124 429436 320180
rect 429492 320124 440188 320180
rect 440244 320124 440254 320180
rect 155474 320012 155484 320068
rect 155540 320012 170492 320068
rect 170548 320012 170558 320068
rect 416658 320012 416668 320068
rect 416724 320012 441084 320068
rect 441140 320012 441150 320068
rect 161970 319676 161980 319732
rect 162036 319676 174104 319732
rect 413896 319676 438844 319732
rect 438900 319676 438910 319732
rect -960 319060 480 319256
rect -960 319032 3388 319060
rect 392 319004 3388 319032
rect 3444 319004 3454 319060
rect 171154 319004 171164 319060
rect 171220 319004 174104 319060
rect 413896 319004 429436 319060
rect 429492 319004 429502 319060
rect 149912 318668 156828 318724
rect 156884 318668 156894 318724
rect 440178 318668 440188 318724
rect 440244 318668 444136 318724
rect 157042 318444 157052 318500
rect 157108 318444 169820 318500
rect 169876 318444 169886 318500
rect 160962 318332 160972 318388
rect 161028 318332 174104 318388
rect 413896 318332 426076 318388
rect 426132 318332 426142 318388
rect 167122 317660 167132 317716
rect 167188 317660 174104 317716
rect 413896 317660 420812 317716
rect 420868 317660 420878 317716
rect 168802 316988 168812 317044
rect 168868 316988 174104 317044
rect 413896 316988 427980 317044
rect 428036 316988 428046 317044
rect 169810 316316 169820 316372
rect 169876 316316 174104 316372
rect 413896 316316 436380 316372
rect 436436 316316 436446 316372
rect 170706 315644 170716 315700
rect 170772 315644 174104 315700
rect 413896 315644 420924 315700
rect 420980 315644 420990 315700
rect 149912 315084 155148 315140
rect 155204 315084 155214 315140
rect 155586 315084 155596 315140
rect 155652 315084 169932 315140
rect 169988 315084 169998 315140
rect 441298 315084 441308 315140
rect 441364 315084 444136 315140
rect 155362 314972 155372 315028
rect 155428 314972 169820 315028
rect 169876 314972 169886 315028
rect 170930 314972 170940 315028
rect 170996 314972 174104 315028
rect 413896 314972 430892 315028
rect 430948 314972 430958 315028
rect 170482 314300 170492 314356
rect 170548 314300 174104 314356
rect 413896 314300 432796 314356
rect 432852 314300 432862 314356
rect 418338 314188 418348 314244
rect 418404 314188 423276 314244
rect 423332 314188 423342 314244
rect 417554 313292 417564 313348
rect 417620 313292 441644 313348
rect 441700 313292 441710 313348
rect 149912 311500 157836 311556
rect 157892 311500 157902 311556
rect 419010 311500 419020 311556
rect 419076 311500 444136 311556
rect 590482 311276 590492 311332
rect 590548 311304 595672 311332
rect 590548 311276 597000 311304
rect 595560 311080 597000 311276
rect 378354 308252 378364 308308
rect 378420 308252 396508 308308
rect 396452 308084 396508 308252
rect 351026 308028 351036 308084
rect 351092 308028 356188 308084
rect 385074 308028 385084 308084
rect 385140 308028 385150 308084
rect 396452 308028 398860 308084
rect 398916 308028 398926 308084
rect 356132 307972 356188 308028
rect 385084 307972 385140 308028
rect 149912 307916 156940 307972
rect 156996 307916 157006 307972
rect 356132 307916 371420 307972
rect 371476 307916 371486 307972
rect 385084 307916 405580 307972
rect 405636 307916 405646 307972
rect 419906 307916 419916 307972
rect 419972 307916 444136 307972
rect 411506 307468 411516 307524
rect 411572 307468 418348 307524
rect 418404 307468 418414 307524
rect 316082 307356 316092 307412
rect 316148 307356 336588 307412
rect 336644 307356 336654 307412
rect 338034 307356 338044 307412
rect 338100 307356 358540 307412
rect 358596 307356 358606 307412
rect 359986 307356 359996 307412
rect 360052 307356 380492 307412
rect 380548 307356 380558 307412
rect 383282 307356 383292 307412
rect 383348 307356 403788 307412
rect 403844 307356 403854 307412
rect 322354 307244 322364 307300
rect 322420 307244 342860 307300
rect 342916 307244 342926 307300
rect 343858 307244 343868 307300
rect 343924 307244 364364 307300
rect 364420 307244 364430 307300
rect 378802 307244 378812 307300
rect 378868 307244 399308 307300
rect 399364 307244 399374 307300
rect 317874 307132 317884 307188
rect 317940 307132 338380 307188
rect 338436 307132 338446 307188
rect 339378 307132 339388 307188
rect 339444 307132 359884 307188
rect 359940 307132 359950 307188
rect 363122 307132 363132 307188
rect 363188 307132 383628 307188
rect 383684 307132 383694 307188
rect 392242 307132 392252 307188
rect 392308 307132 412748 307188
rect 412804 307132 412814 307188
rect 321906 307020 321916 307076
rect 321972 307020 342412 307076
rect 342468 307020 342478 307076
rect 343410 307020 343420 307076
rect 343476 307020 363916 307076
rect 363972 307020 363982 307076
rect 376562 307020 376572 307076
rect 376628 307020 397068 307076
rect 397124 307020 397134 307076
rect 310706 306908 310716 306964
rect 310772 306908 331212 306964
rect 331268 306908 331278 306964
rect 334898 306908 334908 306964
rect 334964 306908 355404 306964
rect 355460 306908 355470 306964
rect 358642 306908 358652 306964
rect 358708 306908 379148 306964
rect 379204 306908 379214 306964
rect 385522 306908 385532 306964
rect 385588 306908 406028 306964
rect 406084 306908 406094 306964
rect 311154 306796 311164 306852
rect 311220 306796 331660 306852
rect 331716 306796 331726 306852
rect 332658 306796 332668 306852
rect 332724 306796 353164 306852
rect 353220 306796 353230 306852
rect 354162 306796 354172 306852
rect 354228 306796 374668 306852
rect 374724 306796 374734 306852
rect 382386 306796 382396 306852
rect 382452 306796 402892 306852
rect 402948 306796 402958 306852
rect 304882 306684 304892 306740
rect 304948 306684 325388 306740
rect 325444 306684 325454 306740
rect 329970 306684 329980 306740
rect 330036 306684 350476 306740
rect 350532 306684 350542 306740
rect 354610 306684 354620 306740
rect 354676 306684 375116 306740
rect 375172 306684 375182 306740
rect 381490 306684 381500 306740
rect 381556 306684 401996 306740
rect 402052 306684 402062 306740
rect 305330 306572 305340 306628
rect 305396 306572 326284 306628
rect 326340 306572 326350 306628
rect 327730 306572 327740 306628
rect 327796 306572 348236 306628
rect 348292 306572 348302 306628
rect 348786 306572 348796 306628
rect 348852 306572 369292 306628
rect 369348 306572 369358 306628
rect 372530 306572 372540 306628
rect 372596 306572 393036 306628
rect 393092 306572 393102 306628
rect 316530 306460 316540 306516
rect 316596 306460 337036 306516
rect 337092 306460 337102 306516
rect 350130 306460 350140 306516
rect 350196 306460 370636 306516
rect 370692 306460 370702 306516
rect 372082 306460 372092 306516
rect 372148 306460 392588 306516
rect 392644 306460 392654 306516
rect 345650 306348 345660 306404
rect 345716 306348 366156 306404
rect 366212 306348 366222 306404
rect 374770 306348 374780 306404
rect 374836 306348 395276 306404
rect 395332 306348 395342 306404
rect 363570 306236 363580 306292
rect 363636 306236 384076 306292
rect 384132 306236 384142 306292
rect 391794 306236 391804 306292
rect 391860 306236 412300 306292
rect 412356 306236 412366 306292
rect 223682 305788 223692 305844
rect 223748 305788 318444 305844
rect 318500 305788 318510 305844
rect 189298 305676 189308 305732
rect 189364 305676 202300 305732
rect 202356 305676 202366 305732
rect 206546 305676 206556 305732
rect 206612 305676 216636 305732
rect 216692 305676 216702 305732
rect 272150 305676 272188 305732
rect 272244 305676 272254 305732
rect 308466 305676 308476 305732
rect 308532 305676 320684 305732
rect 320740 305676 320750 305732
rect 324118 305676 324156 305732
rect 324212 305676 324222 305732
rect 324566 305676 324604 305732
rect 324660 305676 324670 305732
rect 327254 305676 327292 305732
rect 327348 305676 327358 305732
rect 330390 305676 330428 305732
rect 330484 305676 330494 305732
rect 335346 305676 335356 305732
rect 335412 305676 336476 305732
rect 336532 305676 336542 305732
rect 342486 305676 342524 305732
rect 342580 305676 342590 305732
rect 342934 305676 342972 305732
rect 343028 305676 343038 305732
rect 352342 305676 352380 305732
rect 352436 305676 352446 305732
rect 355954 305676 355964 305732
rect 356020 305676 357756 305732
rect 357812 305676 357822 305732
rect 360854 305676 360892 305732
rect 360948 305676 360958 305732
rect 369366 305676 369404 305732
rect 369460 305676 369470 305732
rect 377906 305676 377916 305732
rect 377972 305676 379596 305732
rect 379652 305676 379662 305732
rect 381014 305676 381052 305732
rect 381108 305676 381118 305732
rect 392690 305676 392700 305732
rect 392756 305676 413196 305732
rect 413252 305676 413262 305732
rect 185714 305564 185724 305620
rect 185780 305564 198716 305620
rect 198772 305564 198782 305620
rect 206098 305564 206108 305620
rect 206164 305564 216188 305620
rect 216244 305564 216254 305620
rect 232978 305564 232988 305620
rect 233044 305564 238588 305620
rect 238644 305564 238654 305620
rect 313394 305564 313404 305620
rect 313460 305564 331548 305620
rect 331604 305564 331614 305620
rect 331762 305564 331772 305620
rect 331828 305564 337708 305620
rect 346994 305564 347004 305620
rect 347060 305564 356188 305620
rect 362646 305564 362684 305620
rect 362740 305564 362750 305620
rect 370290 305564 370300 305620
rect 370356 305564 388108 305620
rect 388164 305564 388174 305620
rect 394034 305564 394044 305620
rect 394100 305564 414540 305620
rect 414596 305564 414606 305620
rect 337652 305508 337708 305564
rect 356132 305508 356188 305564
rect 187954 305452 187964 305508
rect 188020 305452 201404 305508
rect 201460 305452 201470 305508
rect 203074 305452 203084 305508
rect 203140 305452 213500 305508
rect 213556 305452 213566 305508
rect 215506 305452 215516 305508
rect 215572 305452 223804 305508
rect 223860 305452 223870 305508
rect 234322 305452 234332 305508
rect 234388 305452 239036 305508
rect 239092 305452 239102 305508
rect 271730 305452 271740 305508
rect 271796 305452 277228 305508
rect 277284 305452 277294 305508
rect 284722 305452 284732 305508
rect 284788 305452 285740 305508
rect 285796 305452 285806 305508
rect 308018 305452 308028 305508
rect 308084 305452 320012 305508
rect 320068 305452 320078 305508
rect 325892 305452 327180 305508
rect 327236 305452 327246 305508
rect 329074 305452 329084 305508
rect 329140 305452 330876 305508
rect 330932 305452 330942 305508
rect 331772 305452 334964 305508
rect 337652 305452 349580 305508
rect 349636 305452 349646 305508
rect 353714 305452 353724 305508
rect 353780 305452 353790 305508
rect 356132 305452 366828 305508
rect 366884 305452 366894 305508
rect 367154 305452 367164 305508
rect 367220 305452 378812 305508
rect 378868 305452 378878 305508
rect 393586 305452 393596 305508
rect 393652 305452 414092 305508
rect 414148 305452 414158 305508
rect 325892 305396 325948 305452
rect 183474 305340 183484 305396
rect 183540 305340 196924 305396
rect 196980 305340 196990 305396
rect 198482 305340 198492 305396
rect 198548 305340 209468 305396
rect 209524 305340 209534 305396
rect 209794 305340 209804 305396
rect 209860 305340 219324 305396
rect 219380 305340 219390 305396
rect 231634 305340 231644 305396
rect 231700 305340 237244 305396
rect 237300 305340 237310 305396
rect 272962 305340 272972 305396
rect 273028 305340 277564 305396
rect 277620 305340 277630 305396
rect 283042 305340 283052 305396
rect 283108 305340 286972 305396
rect 287028 305340 287038 305396
rect 296482 305340 296492 305396
rect 296548 305340 299068 305396
rect 299124 305340 299134 305396
rect 307570 305340 307580 305396
rect 307636 305340 325948 305396
rect 331772 305284 331828 305452
rect 183026 305228 183036 305284
rect 183092 305228 196476 305284
rect 196532 305228 196542 305284
rect 201394 305228 201404 305284
rect 201460 305228 212604 305284
rect 212660 305228 212670 305284
rect 224466 305228 224476 305284
rect 224532 305228 230972 305284
rect 231028 305228 231038 305284
rect 236562 305228 236572 305284
rect 236628 305228 241276 305284
rect 241332 305228 241342 305284
rect 273942 305228 273980 305284
rect 274036 305228 274046 305284
rect 282566 305228 282604 305284
rect 282660 305228 282670 305284
rect 284722 305228 284732 305284
rect 284788 305228 285628 305284
rect 285684 305228 285694 305284
rect 286262 305228 286300 305284
rect 286356 305228 286366 305284
rect 290658 305228 290668 305284
rect 290724 305228 291452 305284
rect 291508 305228 291518 305284
rect 292338 305228 292348 305284
rect 292404 305228 292796 305284
rect 292852 305228 292862 305284
rect 294102 305228 294140 305284
rect 294196 305228 294206 305284
rect 299058 305228 299068 305284
rect 299124 305228 299516 305284
rect 299572 305228 299582 305284
rect 306674 305228 306684 305284
rect 306740 305228 310828 305284
rect 310884 305228 310894 305284
rect 319666 305228 319676 305284
rect 319732 305228 319742 305284
rect 320114 305228 320124 305284
rect 320180 305228 323484 305284
rect 323540 305228 323550 305284
rect 325892 305228 331828 305284
rect 334908 305284 334964 305452
rect 353724 305396 353780 305452
rect 336242 305340 336252 305396
rect 336308 305340 352828 305396
rect 352884 305340 352894 305396
rect 353724 305340 362068 305396
rect 366258 305340 366268 305396
rect 366324 305340 386764 305396
rect 386820 305340 386830 305396
rect 393138 305340 393148 305396
rect 393204 305340 413644 305396
rect 413700 305340 413710 305396
rect 334908 305228 339724 305284
rect 339780 305228 339790 305284
rect 340956 305228 346444 305284
rect 346500 305228 346510 305284
rect 347890 305228 347900 305284
rect 347956 305228 361956 305284
rect 319676 305172 319732 305228
rect 325892 305172 325948 305228
rect -960 304948 480 305144
rect 182578 305116 182588 305172
rect 182644 305116 196028 305172
rect 196084 305116 196094 305172
rect 198706 305116 198716 305172
rect 198772 305116 209916 305172
rect 209972 305116 209982 305172
rect 222002 305116 222012 305172
rect 222068 305116 229628 305172
rect 229684 305116 229694 305172
rect 234770 305116 234780 305172
rect 234836 305116 239484 305172
rect 239540 305116 239550 305172
rect 272626 305116 272636 305172
rect 272692 305116 273868 305172
rect 273924 305116 273934 305172
rect 281362 305116 281372 305172
rect 281428 305116 283836 305172
rect 283892 305116 283902 305172
rect 284946 305116 284956 305172
rect 285012 305116 286524 305172
rect 286580 305116 286590 305172
rect 298274 305116 298284 305172
rect 298340 305116 300860 305172
rect 300916 305116 300926 305172
rect 307122 305116 307132 305172
rect 307188 305116 314188 305172
rect 319676 305116 325948 305172
rect 331314 305116 331324 305172
rect 331380 305116 334236 305172
rect 334292 305116 334302 305172
rect 314132 305060 314188 305116
rect 340956 305060 341012 305228
rect 341170 305116 341180 305172
rect 341236 305116 341246 305172
rect 342066 305116 342076 305172
rect 342132 305116 347788 305172
rect 347844 305116 347854 305172
rect 349412 305116 355348 305172
rect 177202 305004 177212 305060
rect 177268 305004 191100 305060
rect 191156 305004 191166 305060
rect 199714 305004 199724 305060
rect 199780 305004 211260 305060
rect 211316 305004 211326 305060
rect 215954 305004 215964 305060
rect 216020 305004 224700 305060
rect 224756 305004 224766 305060
rect 228386 305004 228396 305060
rect 228452 305004 273084 305060
rect 273140 305004 273150 305060
rect 314132 305004 322588 305060
rect 322644 305004 322654 305060
rect 323372 305004 334796 305060
rect 334852 305004 334862 305060
rect 335010 305004 335020 305060
rect 335076 305004 341012 305060
rect 341180 305060 341236 305116
rect 349412 305060 349468 305116
rect 341180 305004 349468 305060
rect 355292 305060 355348 305116
rect 361900 305060 361956 305228
rect 362012 305172 362068 305340
rect 365810 305228 365820 305284
rect 365876 305228 371084 305284
rect 371140 305228 371150 305284
rect 371634 305228 371644 305284
rect 371700 305228 392140 305284
rect 392196 305228 392206 305284
rect 394454 305228 394492 305284
rect 394548 305228 394558 305284
rect 395826 305228 395836 305284
rect 395892 305228 416332 305284
rect 416388 305228 416398 305284
rect 362012 305116 374220 305172
rect 374276 305116 374286 305172
rect 378802 305116 378812 305172
rect 378868 305116 387660 305172
rect 387716 305116 387726 305172
rect 389106 305116 389116 305172
rect 389172 305116 409612 305172
rect 409668 305116 409678 305172
rect 355292 305004 361676 305060
rect 361732 305004 361742 305060
rect 361890 305004 361900 305060
rect 361956 305004 361966 305060
rect 366706 305004 366716 305060
rect 366772 305004 369908 305060
rect 370738 305004 370748 305060
rect 370804 305004 391244 305060
rect 391300 305004 391310 305060
rect 395378 305004 395388 305060
rect 395444 305004 415884 305060
rect 415940 305004 415950 305060
rect -960 304920 9212 304948
rect 392 304892 9212 304920
rect 9268 304892 9278 304948
rect 154466 304892 154476 304948
rect 154532 304892 169372 304948
rect 169428 304892 169438 304948
rect 178994 304892 179004 304948
rect 179060 304892 192892 304948
rect 192948 304892 192958 304948
rect 204754 304892 204764 304948
rect 204820 304892 271292 304948
rect 271348 304892 271358 304948
rect 278338 304892 278348 304948
rect 278404 304892 282492 304948
rect 282548 304892 282558 304948
rect 285282 304892 285292 304948
rect 285348 304892 295932 304948
rect 295988 304892 295998 304948
rect 302642 304892 302652 304948
rect 302708 304892 323148 304948
rect 323204 304892 323214 304948
rect 323372 304836 323428 305004
rect 325042 304892 325052 304948
rect 325108 304892 345996 304948
rect 346052 304892 346062 304948
rect 346546 304892 346556 304948
rect 346612 304892 356188 304948
rect 356244 304892 356254 304948
rect 356402 304892 356412 304948
rect 356468 304892 364588 304948
rect 364644 304892 364654 304948
rect 189746 304780 189756 304836
rect 189812 304780 202748 304836
rect 202804 304780 202814 304836
rect 209458 304780 209468 304836
rect 209524 304780 218876 304836
rect 218932 304780 218942 304836
rect 230738 304780 230748 304836
rect 230804 304780 236348 304836
rect 236404 304780 236414 304836
rect 241826 304780 241836 304836
rect 241892 304780 245756 304836
rect 245812 304780 245822 304836
rect 314290 304780 314300 304836
rect 314356 304780 323428 304836
rect 323484 304780 330988 304836
rect 331044 304780 331054 304836
rect 336690 304780 336700 304836
rect 336756 304780 349468 304836
rect 352818 304780 352828 304836
rect 352884 304780 356300 304836
rect 356356 304780 356366 304836
rect 192882 304668 192892 304724
rect 192948 304668 204988 304724
rect 205044 304668 205054 304724
rect 209122 304668 209132 304724
rect 209188 304668 218428 304724
rect 218484 304668 218494 304724
rect 241266 304668 241276 304724
rect 241332 304668 245308 304724
rect 245364 304668 245374 304724
rect 308914 304668 308924 304724
rect 308980 304668 320796 304724
rect 320852 304668 320862 304724
rect 323484 304612 323540 304780
rect 325490 304668 325500 304724
rect 325556 304668 342524 304724
rect 342580 304668 342590 304724
rect 349412 304612 349468 304780
rect 369852 304724 369908 305004
rect 372978 304892 372988 304948
rect 373044 304892 393484 304948
rect 393540 304892 393550 304948
rect 396722 304892 396732 304948
rect 396788 304892 417228 304948
rect 417284 304892 417294 304948
rect 375218 304780 375228 304836
rect 375284 304780 384748 304836
rect 387762 304780 387772 304836
rect 387828 304780 394828 304836
rect 394884 304780 394894 304836
rect 384692 304724 384748 304780
rect 356850 304668 356860 304724
rect 356916 304668 367948 304724
rect 369852 304668 383068 304724
rect 383124 304668 383134 304724
rect 384692 304668 388444 304724
rect 388500 304668 388510 304724
rect 388658 304668 388668 304724
rect 388724 304668 402332 304724
rect 402388 304668 402398 304724
rect 367892 304612 367948 304668
rect 196018 304556 196028 304612
rect 196084 304556 208124 304612
rect 208180 304556 208190 304612
rect 211250 304556 211260 304612
rect 211316 304556 220668 304612
rect 220724 304556 220734 304612
rect 226706 304556 226716 304612
rect 226772 304556 233660 304612
rect 233716 304556 233726 304612
rect 240146 304556 240156 304612
rect 240212 304556 243964 304612
rect 244020 304556 244030 304612
rect 315186 304556 315196 304612
rect 315252 304556 323540 304612
rect 326386 304556 326396 304612
rect 326452 304556 341404 304612
rect 341460 304556 341470 304612
rect 349412 304556 351148 304612
rect 351204 304556 351214 304612
rect 351474 304556 351484 304612
rect 351540 304556 366268 304612
rect 366324 304556 366334 304612
rect 367892 304556 372988 304612
rect 373044 304556 373054 304612
rect 373874 304556 373884 304612
rect 373940 304556 376236 304612
rect 376292 304556 376302 304612
rect 380146 304556 380156 304612
rect 380212 304556 393820 304612
rect 393876 304556 393886 304612
rect 191762 304444 191772 304500
rect 191828 304444 200060 304500
rect 200116 304444 200126 304500
rect 226258 304444 226268 304500
rect 226324 304444 232764 304500
rect 232820 304444 232830 304500
rect 244402 304444 244412 304500
rect 244468 304444 247548 304500
rect 247604 304444 247614 304500
rect 320002 304444 320012 304500
rect 320068 304444 326508 304500
rect 326564 304444 326574 304500
rect 341618 304444 341628 304500
rect 341684 304444 354396 304500
rect 354452 304444 354462 304500
rect 361778 304444 361788 304500
rect 361844 304444 377244 304500
rect 377300 304444 377310 304500
rect 384178 304444 384188 304500
rect 384244 304444 393932 304500
rect 393988 304444 393998 304500
rect 149912 304332 153916 304388
rect 153972 304332 153982 304388
rect 225810 304332 225820 304388
rect 225876 304332 232316 304388
rect 232372 304332 232382 304388
rect 243954 304332 243964 304388
rect 244020 304332 247100 304388
rect 247156 304332 247166 304388
rect 278114 304332 278124 304388
rect 278180 304332 281148 304388
rect 281204 304332 281214 304388
rect 323698 304332 323708 304388
rect 323764 304332 329196 304388
rect 329252 304332 329262 304388
rect 330866 304332 330876 304388
rect 330932 304332 349356 304388
rect 349412 304332 349422 304388
rect 361890 304332 361900 304388
rect 361956 304332 368396 304388
rect 368452 304332 368462 304388
rect 416098 304332 416108 304388
rect 416164 304332 444136 304388
rect 214610 304220 214620 304276
rect 214676 304220 222908 304276
rect 222964 304220 222974 304276
rect 225362 304220 225372 304276
rect 225428 304220 231868 304276
rect 231924 304220 231934 304276
rect 233202 304220 233212 304276
rect 233268 304220 311836 304276
rect 311892 304220 311902 304276
rect 325938 304220 325948 304276
rect 326004 304220 335020 304276
rect 335076 304220 335086 304276
rect 351922 304220 351932 304276
rect 351988 304220 371196 304276
rect 371252 304220 371262 304276
rect 391346 304220 391356 304276
rect 391412 304220 398076 304276
rect 398132 304220 398142 304276
rect 214162 304108 214172 304164
rect 214228 304108 222460 304164
rect 222516 304108 222526 304164
rect 233650 304108 233660 304164
rect 233716 304108 315084 304164
rect 315140 304108 315150 304164
rect 327702 304108 327740 304164
rect 327796 304108 327806 304164
rect 344614 304108 344652 304164
rect 344708 304108 344718 304164
rect 355814 304108 355852 304164
rect 355908 304108 355918 304164
rect 356178 304108 356188 304164
rect 356244 304108 367500 304164
rect 367556 304108 367566 304164
rect 368498 304108 368508 304164
rect 368564 304108 371308 304164
rect 371364 304108 371374 304164
rect 376422 304108 376460 304164
rect 376516 304108 376526 304164
rect 388434 304108 388444 304164
rect 388500 304108 393204 304164
rect 401510 304108 401548 304164
rect 401604 304108 401614 304164
rect 405234 304108 405244 304164
rect 405300 304108 411516 304164
rect 411572 304108 411582 304164
rect 393148 304052 393204 304108
rect 186610 303996 186620 304052
rect 186676 303996 199612 304052
rect 199668 303996 199678 304052
rect 202738 303996 202748 304052
rect 202804 303996 213052 304052
rect 213108 303996 213118 304052
rect 219314 303996 219324 304052
rect 219380 303996 226940 304052
rect 226996 303996 227006 304052
rect 235890 303996 235900 304052
rect 235956 303996 240828 304052
rect 240884 303996 240894 304052
rect 249666 303996 249676 304052
rect 249732 303996 251580 304052
rect 251636 303996 251646 304052
rect 252466 303996 252476 304052
rect 252532 303996 253820 304052
rect 253876 303996 253886 304052
rect 303986 303996 303996 304052
rect 304052 303996 309148 304052
rect 309204 303996 309214 304052
rect 318322 303996 318332 304052
rect 318388 303996 338828 304052
rect 338884 303996 338894 304052
rect 344754 303996 344764 304052
rect 344820 303996 365260 304052
rect 365316 303996 365326 304052
rect 366258 303996 366268 304052
rect 366324 303996 371980 304052
rect 372036 303996 372046 304052
rect 375666 303996 375676 304052
rect 375732 303996 377580 304052
rect 377636 303996 377646 304052
rect 380594 303996 380604 304052
rect 380660 303996 383964 304052
rect 384020 303996 384030 304052
rect 388098 303996 388108 304052
rect 388164 303996 390796 304052
rect 390852 303996 390862 304052
rect 393148 303996 395724 304052
rect 395780 303996 395790 304052
rect 395938 303996 395948 304052
rect 396004 303996 407372 304052
rect 407428 303996 407438 304052
rect 180338 303884 180348 303940
rect 180404 303884 193788 303940
rect 193844 303884 193854 303940
rect 204306 303884 204316 303940
rect 204372 303884 214396 303940
rect 214452 303884 214462 303940
rect 216178 303884 216188 303940
rect 216244 303884 224252 303940
rect 224308 303884 224318 303940
rect 224690 303884 224700 303940
rect 224756 303884 231420 303940
rect 231476 303884 231486 303940
rect 236674 303884 236684 303940
rect 236740 303884 241724 303940
rect 241780 303884 241790 303940
rect 250898 303884 250908 303940
rect 250964 303884 252588 303940
rect 252644 303884 252654 303940
rect 252914 303884 252924 303940
rect 252980 303884 254268 303940
rect 254324 303884 254334 303940
rect 312498 303884 312508 303940
rect 312564 303884 333004 303940
rect 333060 303884 333070 303940
rect 334002 303884 334012 303940
rect 334068 303884 336028 303940
rect 336084 303884 336094 303940
rect 339826 303884 339836 303940
rect 339892 303884 360332 303940
rect 360388 303884 360398 303940
rect 368946 303884 368956 303940
rect 369012 303884 389452 303940
rect 389508 303884 389518 303940
rect 390898 303884 390908 303940
rect 390964 303884 411404 303940
rect 411460 303884 411470 303940
rect 180786 303772 180796 303828
rect 180852 303772 194236 303828
rect 194292 303772 194302 303828
rect 200050 303772 200060 303828
rect 200116 303772 210812 303828
rect 210868 303772 210878 303828
rect 216626 303772 216636 303828
rect 216692 303772 225148 303828
rect 225204 303772 225214 303828
rect 234994 303772 235004 303828
rect 235060 303772 239932 303828
rect 239988 303772 239998 303828
rect 249218 303772 249228 303828
rect 249284 303772 251132 303828
rect 251188 303772 251198 303828
rect 253362 303772 253372 303828
rect 253428 303772 254716 303828
rect 254772 303772 254782 303828
rect 311602 303772 311612 303828
rect 311668 303772 332108 303828
rect 332164 303772 332174 303828
rect 338930 303772 338940 303828
rect 338996 303772 359436 303828
rect 359492 303772 359502 303828
rect 364018 303772 364028 303828
rect 364084 303772 384524 303828
rect 384580 303772 384590 303828
rect 386866 303772 386876 303828
rect 386932 303772 386942 303828
rect 390002 303772 390012 303828
rect 390068 303772 410508 303828
rect 410564 303772 410574 303828
rect 386876 303716 386932 303772
rect 181234 303660 181244 303716
rect 181300 303660 194684 303716
rect 194740 303660 194750 303716
rect 197922 303660 197932 303716
rect 197988 303660 209020 303716
rect 209076 303660 209086 303716
rect 229618 303660 229628 303716
rect 229684 303660 235452 303716
rect 235508 303660 235518 303716
rect 304434 303660 304444 303716
rect 304500 303660 324940 303716
rect 324996 303660 325006 303716
rect 327170 303660 327180 303716
rect 327236 303660 328524 303716
rect 328580 303660 328590 303716
rect 330978 303660 330988 303716
rect 331044 303660 335692 303716
rect 335748 303660 335758 303716
rect 338482 303660 338492 303716
rect 338548 303660 358988 303716
rect 359044 303660 359054 303716
rect 359538 303660 359548 303716
rect 359604 303660 380044 303716
rect 380100 303660 380110 303716
rect 386876 303660 395948 303716
rect 396004 303660 396014 303716
rect 396162 303660 396172 303716
rect 396228 303660 406924 303716
rect 406980 303660 406990 303716
rect 178098 303548 178108 303604
rect 178164 303548 191996 303604
rect 192052 303548 192062 303604
rect 193554 303548 193564 303604
rect 193620 303548 205436 303604
rect 205492 303548 205502 303604
rect 212370 303548 212380 303604
rect 212436 303548 221564 303604
rect 221620 303548 221630 303604
rect 229954 303548 229964 303604
rect 230020 303548 235564 303604
rect 235620 303548 235630 303604
rect 312050 303548 312060 303604
rect 312116 303548 332556 303604
rect 332612 303548 332622 303604
rect 333554 303548 333564 303604
rect 333620 303548 354060 303604
rect 354116 303548 354126 303604
rect 359090 303548 359100 303604
rect 359156 303548 379596 303604
rect 379652 303548 379662 303604
rect 381938 303548 381948 303604
rect 382004 303548 402444 303604
rect 402500 303548 402510 303604
rect 178546 303436 178556 303492
rect 178612 303436 192444 303492
rect 192500 303436 192510 303492
rect 193778 303436 193788 303492
rect 193844 303436 206332 303492
rect 206388 303436 206398 303492
rect 210466 303436 210476 303492
rect 210532 303436 220220 303492
rect 220276 303436 220286 303492
rect 222450 303436 222460 303492
rect 222516 303436 230076 303492
rect 230132 303436 230142 303492
rect 235442 303436 235452 303492
rect 235508 303436 240380 303492
rect 240436 303436 240446 303492
rect 303538 303436 303548 303492
rect 303604 303436 324044 303492
rect 324100 303436 324110 303492
rect 328178 303436 328188 303492
rect 328244 303436 348684 303492
rect 348740 303436 348750 303492
rect 355058 303436 355068 303492
rect 355124 303436 372988 303492
rect 376226 303436 376236 303492
rect 376292 303436 394380 303492
rect 394436 303436 394446 303492
rect 394930 303436 394940 303492
rect 394996 303436 415436 303492
rect 415492 303436 415502 303492
rect 184370 303324 184380 303380
rect 184436 303324 198268 303380
rect 198324 303324 198334 303380
rect 204978 303324 204988 303380
rect 205044 303324 215740 303380
rect 215796 303324 215806 303380
rect 217746 303324 217756 303380
rect 217812 303324 226044 303380
rect 226100 303324 226110 303380
rect 232306 303324 232316 303380
rect 232372 303324 238140 303380
rect 238196 303324 238206 303380
rect 315634 303324 315644 303380
rect 315700 303324 319004 303380
rect 319060 303324 319070 303380
rect 319218 303324 319228 303380
rect 319284 303324 340172 303380
rect 340228 303324 340238 303380
rect 345202 303324 345212 303380
rect 345268 303324 365708 303380
rect 365764 303324 365774 303380
rect 372932 303268 372988 303436
rect 373426 303324 373436 303380
rect 373492 303324 393708 303380
rect 393764 303324 393774 303380
rect 396274 303324 396284 303380
rect 396340 303324 416780 303380
rect 416836 303324 416846 303380
rect 160514 303212 160524 303268
rect 160580 303212 171164 303268
rect 171220 303212 171230 303268
rect 179890 303212 179900 303268
rect 179956 303212 197820 303268
rect 197876 303212 197886 303268
rect 199154 303212 199164 303268
rect 199220 303212 210364 303268
rect 210420 303212 210430 303268
rect 210802 303212 210812 303268
rect 210868 303212 219772 303268
rect 219828 303212 219838 303268
rect 221554 303212 221564 303268
rect 221620 303212 228732 303268
rect 228788 303212 228798 303268
rect 243506 303212 243516 303268
rect 243572 303212 246652 303268
rect 246708 303212 246718 303268
rect 247986 303212 247996 303268
rect 248052 303212 250236 303268
rect 250292 303212 250302 303268
rect 305778 303212 305788 303268
rect 305844 303212 326732 303268
rect 326788 303212 326798 303268
rect 328626 303212 328636 303268
rect 328692 303212 349132 303268
rect 349188 303212 349198 303268
rect 349682 303212 349692 303268
rect 349748 303212 355348 303268
rect 355506 303212 355516 303268
rect 355572 303212 364588 303268
rect 372932 303212 375340 303268
rect 375396 303212 375406 303268
rect 377458 303212 377468 303268
rect 377524 303212 397964 303268
rect 398020 303212 398030 303268
rect 429426 303212 429436 303268
rect 429492 303212 440972 303268
rect 441028 303212 441038 303268
rect 187058 303100 187068 303156
rect 187124 303100 191772 303156
rect 191828 303100 191838 303156
rect 192434 303100 192444 303156
rect 192500 303100 204540 303156
rect 204596 303100 204606 303156
rect 205426 303100 205436 303156
rect 205492 303100 215292 303156
rect 215348 303100 215358 303156
rect 243058 303100 243068 303156
rect 243124 303100 246204 303156
rect 246260 303100 246270 303156
rect 247538 303100 247548 303156
rect 247604 303100 249788 303156
rect 249844 303100 249854 303156
rect 323250 303100 323260 303156
rect 323316 303100 343756 303156
rect 343812 303100 343822 303156
rect 355292 303044 355348 303212
rect 364532 303156 364588 303212
rect 364532 303100 376012 303156
rect 376068 303100 376078 303156
rect 381350 303100 381388 303156
rect 381444 303100 381454 303156
rect 386418 303100 386428 303156
rect 386484 303100 386494 303156
rect 389862 303100 389900 303156
rect 389956 303100 389966 303156
rect 398374 303100 398412 303156
rect 398468 303100 398478 303156
rect 386428 303044 386484 303100
rect 191986 302988 191996 303044
rect 192052 302988 204092 303044
rect 204148 302988 204158 303044
rect 245298 302988 245308 303044
rect 245364 302988 248444 303044
rect 248500 302988 248510 303044
rect 334450 302988 334460 303044
rect 334516 302988 354956 303044
rect 355012 302988 355022 303044
rect 355292 302988 370244 303044
rect 370188 302932 370244 302988
rect 370412 302988 385420 303044
rect 385476 302988 385486 303044
rect 386428 302988 396172 303044
rect 396228 302988 396238 303044
rect 396452 302988 407820 303044
rect 407876 302988 407886 303044
rect 191762 302876 191772 302932
rect 191828 302876 203644 302932
rect 203700 302876 203710 302932
rect 204530 302876 204540 302932
rect 204596 302876 214844 302932
rect 214900 302876 214910 302932
rect 255154 302876 255164 302932
rect 255220 302876 256508 302932
rect 256564 302876 256574 302932
rect 329186 302876 329196 302932
rect 329252 302876 344204 302932
rect 344260 302876 344270 302932
rect 351026 302876 351036 302932
rect 351092 302876 354508 302932
rect 354564 302876 354574 302932
rect 361330 302876 361340 302932
rect 361396 302876 369516 302932
rect 369572 302876 369582 302932
rect 370178 302876 370188 302932
rect 370244 302876 370254 302932
rect 370412 302820 370468 302988
rect 371298 302876 371308 302932
rect 371364 302876 389004 302932
rect 389060 302876 389070 302932
rect 396452 302820 396508 302988
rect 398066 302876 398076 302932
rect 398132 302876 411852 302932
rect 411908 302876 411918 302932
rect 238130 302764 238140 302820
rect 238196 302764 238588 302820
rect 254706 302764 254716 302820
rect 254772 302764 256060 302820
rect 256116 302764 256126 302820
rect 324454 302764 324492 302820
rect 324548 302764 324558 302820
rect 364914 302764 364924 302820
rect 364980 302764 370468 302820
rect 387314 302764 387324 302820
rect 387380 302764 396508 302820
rect 203634 302652 203644 302708
rect 203700 302652 213948 302708
rect 214004 302652 214014 302708
rect 211922 302540 211932 302596
rect 211988 302540 221116 302596
rect 221172 302540 221182 302596
rect 238532 302484 238588 302764
rect 254258 302652 254268 302708
rect 254324 302652 255612 302708
rect 255668 302652 255678 302708
rect 256274 302652 256284 302708
rect 256340 302652 314972 302708
rect 315028 302652 315038 302708
rect 242946 302540 242956 302596
rect 243012 302540 318332 302596
rect 318388 302540 318398 302596
rect 322578 302540 322588 302596
rect 322644 302540 328076 302596
rect 328132 302540 328142 302596
rect 347778 302540 347788 302596
rect 347844 302540 349580 302596
rect 349636 302540 349646 302596
rect 354386 302540 354396 302596
rect 354452 302540 361676 302596
rect 361732 302540 361742 302596
rect 213490 302428 213500 302484
rect 213556 302428 221788 302484
rect 221844 302428 221854 302484
rect 226930 302428 226940 302484
rect 226996 302428 232876 302484
rect 232932 302428 232942 302484
rect 238532 302428 318556 302484
rect 318612 302428 318622 302484
rect 321010 302428 321020 302484
rect 321076 302428 322644 302484
rect 363430 302428 363468 302484
rect 363524 302428 363534 302484
rect 383058 302428 383068 302484
rect 383124 302428 387212 302484
rect 387268 302428 387278 302484
rect 402322 302428 402332 302484
rect 402388 302428 409164 302484
rect 409220 302428 409230 302484
rect 322588 302372 322644 302428
rect 188850 302316 188860 302372
rect 188916 302316 201852 302372
rect 201908 302316 201918 302372
rect 238578 302316 238588 302372
rect 238644 302316 242620 302372
rect 242676 302316 242686 302372
rect 244850 302316 244860 302372
rect 244916 302316 247660 302372
rect 247716 302316 247726 302372
rect 322588 302316 341516 302372
rect 341572 302316 341582 302372
rect 367574 302316 367612 302372
rect 367668 302316 367678 302372
rect 377570 302316 377580 302372
rect 377636 302316 396172 302372
rect 396228 302316 396238 302372
rect 186162 302204 186172 302260
rect 186228 302204 199052 302260
rect 199108 302204 199118 302260
rect 218866 302204 218876 302260
rect 218932 302204 226492 302260
rect 226548 302204 226558 302260
rect 239026 302204 239036 302260
rect 239092 302204 242732 302260
rect 242788 302204 242798 302260
rect 245746 302204 245756 302260
rect 245812 302204 248892 302260
rect 248948 302204 248958 302260
rect 314738 302204 314748 302260
rect 314804 302204 335244 302260
rect 335300 302204 335310 302260
rect 357746 302204 357756 302260
rect 357812 302204 378252 302260
rect 378308 302204 378318 302260
rect 389554 302204 389564 302260
rect 389620 302204 393148 302260
rect 393204 302204 393214 302260
rect 394818 302204 394828 302260
rect 394884 302204 408268 302260
rect 408324 302204 408334 302260
rect 190194 302092 190204 302148
rect 190260 302092 203196 302148
rect 203252 302092 203262 302148
rect 206770 302092 206780 302148
rect 206836 302092 217084 302148
rect 217140 302092 217150 302148
rect 220658 302092 220668 302148
rect 220724 302092 228284 302148
rect 228340 302092 228350 302148
rect 239474 302092 239484 302148
rect 239540 302092 243180 302148
rect 243236 302092 243246 302148
rect 246194 302092 246204 302148
rect 246260 302092 249340 302148
rect 249396 302092 249406 302148
rect 321458 302092 321468 302148
rect 321524 302092 341964 302148
rect 342020 302092 342030 302148
rect 357298 302092 357308 302148
rect 357364 302092 374164 302148
rect 374294 302092 374332 302148
rect 374388 302092 374398 302148
rect 383954 302092 383964 302148
rect 384020 302092 401100 302148
rect 401156 302092 401166 302148
rect 374108 302036 374164 302092
rect 182130 301980 182140 302036
rect 182196 301980 195580 302036
rect 195636 301980 195646 302036
rect 197362 301980 197372 302036
rect 197428 301980 208572 302036
rect 208628 301980 208638 302036
rect 220210 301980 220220 302036
rect 220276 301980 227836 302036
rect 227892 301980 227902 302036
rect 230962 301980 230972 302036
rect 231028 301980 236796 302036
rect 236852 301980 236862 302036
rect 240370 301980 240380 302036
rect 240436 301980 244076 302036
rect 244132 301980 244142 302036
rect 320562 301980 320572 302036
rect 320628 301980 341068 302036
rect 341124 301980 341134 302036
rect 344278 301980 344316 302036
rect 344372 301980 344382 302036
rect 353266 301980 353276 302036
rect 353332 301980 373772 302036
rect 373828 301980 373838 302036
rect 374108 301980 377804 302036
rect 377860 301980 377870 302036
rect 384626 301980 384636 302036
rect 384692 301980 405132 302036
rect 405188 301980 405198 302036
rect 181682 301868 181692 301924
rect 181748 301868 195132 301924
rect 195188 301868 195198 301924
rect 201282 301868 201292 301924
rect 201348 301868 212156 301924
rect 212212 301868 212222 301924
rect 214834 301868 214844 301924
rect 214900 301868 223356 301924
rect 223412 301868 223422 301924
rect 228274 301868 228284 301924
rect 228340 301868 234892 301924
rect 234948 301868 234958 301924
rect 240818 301868 240828 301924
rect 240884 301868 244524 301924
rect 244580 301868 244590 301924
rect 309810 301868 309820 301924
rect 309876 301868 330316 301924
rect 330372 301868 330382 301924
rect 337138 301868 337148 301924
rect 337204 301868 357644 301924
rect 357700 301868 357710 301924
rect 379698 301868 379708 301924
rect 379764 301868 400204 301924
rect 400260 301868 400270 301924
rect 417442 301868 417452 301924
rect 417508 301868 424620 301924
rect 424676 301868 424686 301924
rect 183922 301756 183932 301812
rect 183988 301756 197260 301812
rect 197316 301756 197326 301812
rect 200834 301756 200844 301812
rect 200900 301756 211708 301812
rect 211764 301756 211774 301812
rect 217074 301756 217084 301812
rect 217140 301756 225596 301812
rect 225652 301756 225662 301812
rect 227826 301756 227836 301812
rect 227892 301756 234556 301812
rect 234612 301756 234622 301812
rect 312946 301756 312956 301812
rect 313012 301756 333452 301812
rect 333508 301756 333518 301812
rect 337586 301756 337596 301812
rect 337652 301756 358092 301812
rect 358148 301756 358158 301812
rect 362226 301756 362236 301812
rect 362292 301756 382732 301812
rect 382788 301756 382798 301812
rect 383730 301756 383740 301812
rect 383796 301756 404236 301812
rect 404292 301756 404302 301812
rect 417666 301756 417676 301812
rect 417732 301756 436716 301812
rect 436772 301756 436782 301812
rect 179442 301644 179452 301700
rect 179508 301644 193340 301700
rect 193396 301644 193406 301700
rect 195570 301644 195580 301700
rect 195636 301644 207676 301700
rect 207732 301644 207742 301700
rect 208114 301644 208124 301700
rect 208180 301644 217532 301700
rect 217588 301644 217598 301700
rect 219762 301644 219772 301700
rect 219828 301644 227388 301700
rect 227444 301644 227454 301700
rect 303090 301644 303100 301700
rect 303156 301644 323596 301700
rect 323652 301644 323662 301700
rect 326834 301644 326844 301700
rect 326900 301644 347340 301700
rect 347396 301644 347406 301700
rect 352818 301644 352828 301700
rect 352884 301644 373324 301700
rect 373380 301644 373390 301700
rect 376114 301644 376124 301700
rect 376180 301644 396620 301700
rect 396676 301644 396686 301700
rect 415986 301644 415996 301700
rect 416052 301644 441420 301700
rect 441476 301644 441486 301700
rect 177650 301532 177660 301588
rect 177716 301532 191548 301588
rect 191604 301532 191614 301588
rect 194674 301532 194684 301588
rect 194740 301532 206668 301588
rect 206724 301532 206734 301588
rect 306226 301532 306236 301588
rect 306292 301532 327180 301588
rect 327236 301532 327246 301588
rect 335794 301532 335804 301588
rect 335860 301532 356748 301588
rect 356804 301532 356814 301588
rect 358194 301532 358204 301588
rect 358260 301532 378700 301588
rect 378756 301532 378766 301588
rect 379250 301532 379260 301588
rect 379316 301532 399756 301588
rect 399812 301532 399822 301588
rect 415762 301532 415772 301588
rect 415828 301532 441756 301588
rect 441812 301532 441822 301588
rect 188402 301420 188412 301476
rect 188468 301420 200956 301476
rect 201012 301420 201022 301476
rect 202290 301420 202300 301476
rect 202356 301420 321692 301476
rect 321748 301420 321758 301476
rect 323474 301420 323484 301476
rect 323540 301420 340620 301476
rect 340676 301420 340686 301476
rect 347442 301420 347452 301476
rect 347508 301420 367948 301476
rect 368004 301420 368014 301476
rect 371074 301420 371084 301476
rect 371140 301420 386316 301476
rect 386372 301420 386382 301476
rect 393922 301420 393932 301476
rect 393988 301420 404684 301476
rect 404740 301420 404750 301476
rect 195122 301308 195132 301364
rect 195188 301308 207228 301364
rect 207284 301308 207294 301364
rect 227378 301308 227388 301364
rect 227444 301308 234108 301364
rect 234164 301308 234174 301364
rect 309362 301308 309372 301364
rect 309428 301308 325836 301364
rect 325892 301308 325902 301364
rect 334226 301308 334236 301364
rect 334292 301308 351820 301364
rect 351876 301308 351886 301364
rect 357746 301308 357756 301364
rect 357812 301308 363020 301364
rect 363076 301308 363086 301364
rect 369506 301308 369516 301364
rect 369572 301308 381836 301364
rect 381892 301308 381902 301364
rect 393810 301308 393820 301364
rect 393876 301308 400652 301364
rect 400708 301308 400718 301364
rect 194226 301196 194236 301252
rect 194292 301196 205884 301252
rect 205940 301196 205950 301252
rect 237234 301196 237244 301252
rect 237300 301196 242172 301252
rect 242228 301196 242238 301252
rect 247090 301196 247100 301252
rect 247156 301196 252588 301252
rect 252644 301196 252654 301252
rect 347778 301196 347788 301252
rect 347844 301196 362572 301252
rect 362628 301196 362638 301252
rect 251122 301084 251132 301140
rect 251188 301084 310828 301140
rect 310884 301084 310894 301140
rect 341394 301084 341404 301140
rect 341460 301084 346892 301140
rect 346948 301084 346958 301140
rect 348338 301084 348348 301140
rect 348404 301084 368844 301140
rect 368900 301084 368910 301140
rect 221106 300972 221116 301028
rect 221172 300972 229180 301028
rect 229236 300972 229246 301028
rect 248434 300972 248444 301028
rect 248500 300972 250684 301028
rect 250740 300972 250750 301028
rect 251570 300972 251580 301028
rect 251636 300972 315196 301028
rect 315252 300972 315262 301028
rect 344418 300972 344428 301028
rect 344484 300972 347788 301028
rect 347844 300972 347854 301028
rect 349346 300972 349356 301028
rect 349412 300972 350924 301028
rect 350980 300972 350990 301028
rect 351138 300972 351148 301028
rect 351204 300972 357196 301028
rect 357252 300972 357262 301028
rect 222898 300860 222908 300916
rect 222964 300860 230524 300916
rect 230580 300860 230590 300916
rect 250226 300860 250236 300916
rect 250292 300860 252364 300916
rect 252420 300860 252430 300916
rect 252578 300860 252588 300916
rect 252644 300860 318892 300916
rect 318948 300860 318958 300916
rect 332546 300860 332556 300916
rect 332612 300860 336140 300916
rect 336196 300860 336206 300916
rect 342514 300860 342524 300916
rect 342580 300860 345548 300916
rect 345604 300860 345614 300916
rect 349570 300860 349580 300916
rect 349636 300860 352268 300916
rect 352324 300860 352334 300916
rect 371186 300860 371196 300916
rect 371252 300860 372876 300916
rect 372932 300860 372942 300916
rect 374546 300860 374556 300916
rect 374612 300860 376908 300916
rect 376964 300860 376974 300916
rect 377234 300860 377244 300916
rect 377300 300860 382284 300916
rect 382340 300860 382350 300916
rect 149912 300748 160300 300804
rect 160356 300748 160366 300804
rect 208562 300748 208572 300804
rect 208628 300748 217980 300804
rect 218036 300748 218046 300804
rect 218390 300748 218428 300804
rect 218484 300748 218494 300804
rect 228694 300748 228732 300804
rect 228788 300748 228798 300804
rect 229142 300748 229180 300804
rect 229236 300748 229246 300804
rect 231858 300748 231868 300804
rect 231924 300748 237692 300804
rect 237748 300748 237758 300804
rect 242134 300748 242172 300804
rect 242228 300748 242238 300804
rect 249778 300748 249788 300804
rect 249844 300748 252028 300804
rect 252084 300748 252094 300804
rect 260502 300748 260540 300804
rect 260596 300748 260606 300804
rect 326498 300748 326508 300804
rect 326564 300748 328972 300804
rect 329028 300748 329038 300804
rect 329382 300748 329420 300804
rect 329476 300748 329486 300804
rect 329830 300748 329868 300804
rect 329924 300748 329934 300804
rect 331538 300748 331548 300804
rect 331604 300748 334348 300804
rect 334404 300748 334414 300804
rect 342626 300748 342636 300804
rect 342692 300748 345100 300804
rect 345156 300748 345166 300804
rect 351334 300748 351372 300804
rect 351428 300748 351438 300804
rect 364774 300748 364812 300804
rect 364868 300748 364878 300804
rect 372390 300748 372428 300804
rect 372484 300748 372494 300804
rect 372978 300748 372988 300804
rect 373044 300748 377356 300804
rect 377412 300748 377422 300804
rect 379698 300748 379708 300804
rect 379764 300748 383180 300804
rect 383236 300748 383246 300804
rect 388070 300748 388108 300804
rect 388164 300748 388174 300804
rect 394790 300748 394828 300804
rect 394884 300748 394894 300804
rect 399746 300748 399756 300804
rect 399812 300748 410060 300804
rect 410116 300748 410126 300804
rect 414950 300748 414988 300804
rect 415044 300748 415054 300804
rect 440738 300748 440748 300804
rect 440804 300748 444136 300804
rect 171602 300636 171612 300692
rect 171668 300636 176204 300692
rect 176260 300636 176270 300692
rect 360434 300524 360444 300580
rect 360500 300524 380940 300580
rect 380996 300524 381006 300580
rect 385970 300524 385980 300580
rect 386036 300524 406476 300580
rect 406532 300524 406542 300580
rect 313842 300412 313852 300468
rect 313908 300412 333900 300468
rect 333956 300412 333966 300468
rect 365362 300412 365372 300468
rect 365428 300412 385868 300468
rect 385924 300412 385934 300468
rect 322802 300300 322812 300356
rect 322868 300300 343308 300356
rect 343364 300300 343374 300356
rect 349234 300300 349244 300356
rect 349300 300300 369740 300356
rect 369796 300300 369806 300356
rect 388210 300300 388220 300356
rect 388276 300300 408716 300356
rect 408772 300300 408782 300356
rect 329522 300188 329532 300244
rect 329588 300188 350028 300244
rect 350084 300188 350094 300244
rect 350578 300188 350588 300244
rect 350644 300188 371084 300244
rect 371140 300188 371150 300244
rect 382834 300188 382844 300244
rect 382900 300188 403340 300244
rect 403396 300188 403406 300244
rect 316978 300076 316988 300132
rect 317044 300076 337484 300132
rect 337540 300076 337550 300132
rect 346098 300076 346108 300132
rect 346164 300076 366604 300132
rect 366660 300076 366670 300132
rect 368050 300076 368060 300132
rect 368116 300076 388556 300132
rect 388612 300076 388622 300132
rect 390450 300076 390460 300132
rect 390516 300076 410956 300132
rect 411012 300076 411022 300132
rect 187506 299964 187516 300020
rect 187572 299964 200508 300020
rect 200564 299964 200574 300020
rect 318770 299964 318780 300020
rect 318836 299964 339276 300020
rect 339332 299964 339342 300020
rect 340274 299964 340284 300020
rect 340340 299964 360780 300020
rect 360836 299964 360846 300020
rect 369842 299964 369852 300020
rect 369908 299964 390348 300020
rect 390404 299964 390414 300020
rect 174290 299852 174300 299908
rect 174356 299852 228396 299908
rect 228452 299852 228462 299908
rect 310258 299852 310268 299908
rect 310324 299852 330764 299908
rect 330820 299852 330830 299908
rect 333106 299852 333116 299908
rect 333172 299852 353612 299908
rect 353668 299852 353678 299908
rect 377010 299852 377020 299908
rect 377076 299852 397516 299908
rect 397572 299852 397582 299908
rect 212594 299516 212604 299572
rect 212660 299516 220108 299572
rect 223318 299516 223356 299572
rect 223412 299516 223422 299572
rect 237654 299516 237692 299572
rect 237748 299516 237758 299572
rect 220052 299460 220108 299516
rect 217942 299404 217980 299460
rect 218036 299404 218046 299460
rect 220052 299404 428540 299460
rect 428596 299404 428606 299460
rect 207218 299292 207228 299348
rect 207284 299292 430108 299348
rect 430164 299292 430174 299348
rect 201842 299180 201852 299236
rect 201908 299180 428428 299236
rect 428484 299180 428494 299236
rect 191090 299068 191100 299124
rect 191156 299068 420140 299124
rect 420196 299068 420206 299124
rect 196532 298956 204764 299012
rect 204820 298956 204830 299012
rect 246866 298956 246876 299012
rect 246932 298956 442988 299012
rect 443044 298956 443054 299012
rect 196532 298788 196588 298956
rect 213042 298844 213052 298900
rect 213108 298844 423724 298900
rect 423780 298844 423790 298900
rect 172274 298732 172284 298788
rect 172340 298732 196588 298788
rect 207666 298732 207676 298788
rect 207732 298732 414092 298788
rect 414148 298732 414158 298788
rect 418002 298732 418012 298788
rect 418068 298732 421148 298788
rect 421204 298732 421214 298788
rect 196914 298620 196924 298676
rect 196980 298620 426748 298676
rect 426804 298620 426814 298676
rect 190642 298508 190652 298564
rect 190708 298508 423612 298564
rect 423668 298508 423678 298564
rect 196466 298396 196476 298452
rect 196532 298396 430220 298452
rect 430276 298396 430286 298452
rect 184818 298284 184828 298340
rect 184884 298284 184894 298340
rect 185266 298284 185276 298340
rect 185332 298284 238588 298340
rect 255574 298284 255612 298340
rect 255668 298284 255678 298340
rect 260054 298284 260092 298340
rect 260148 298284 260158 298340
rect 267092 298284 314188 298340
rect 319106 298284 319116 298340
rect 319172 298284 322028 298340
rect 322084 298284 322094 298340
rect 332294 298284 332332 298340
rect 332388 298284 332398 298340
rect 337922 298284 337932 298340
rect 337988 298284 338212 298340
rect 340834 298284 340844 298340
rect 340900 298284 341124 298340
rect 352678 298284 352716 298340
rect 352772 298284 352782 298340
rect 358652 298284 361228 298340
rect 361284 298284 361294 298340
rect 364130 298284 364140 298340
rect 364196 298284 367948 298340
rect 184828 298004 184884 298284
rect 238532 298228 238588 298284
rect 267092 298228 267148 298284
rect 238532 298172 267148 298228
rect 314132 298228 314188 298284
rect 314132 298172 337708 298228
rect 337764 298172 337774 298228
rect 338156 298116 338212 298284
rect 317426 298060 317436 298116
rect 317492 298060 338212 298116
rect 341068 298116 341124 298284
rect 343522 298172 343532 298228
rect 343588 298172 356188 298228
rect 356244 298172 356254 298228
rect 358652 298116 358708 298284
rect 341068 298060 358708 298116
rect 367892 298004 367948 298284
rect 370636 298284 370860 298340
rect 370916 298284 370926 298340
rect 384934 298284 384972 298340
rect 385028 298284 385038 298340
rect 387996 298284 391692 298340
rect 391748 298284 391758 298340
rect 396452 298284 423388 298340
rect 423444 298284 423454 298340
rect 370636 298116 370692 298284
rect 371074 298172 371084 298228
rect 371140 298172 384860 298228
rect 384916 298172 384926 298228
rect 387996 298116 388052 298284
rect 370636 298060 388052 298116
rect 184828 297948 318668 298004
rect 318724 297948 318734 298004
rect 332322 297948 332332 298004
rect 332388 297948 352716 298004
rect 352772 297948 352782 298004
rect 367892 297948 384972 298004
rect 385028 297948 385038 298004
rect 396452 297892 396508 298284
rect 414082 298060 414092 298116
rect 414148 298060 420028 298116
rect 420084 298060 420094 298116
rect 590706 298060 590716 298116
rect 590772 298088 595672 298116
rect 590772 298060 597000 298088
rect 337698 297836 337708 297892
rect 337764 297836 343532 297892
rect 343588 297836 343598 297892
rect 356178 297836 356188 297892
rect 356244 297836 371084 297892
rect 371140 297836 371150 297892
rect 384850 297836 384860 297892
rect 384916 297836 396508 297892
rect 595560 297864 597000 298060
rect 149912 297164 164220 297220
rect 164276 297164 164286 297220
rect 437378 297164 437388 297220
rect 437444 297164 444136 297220
rect 255602 296940 255612 296996
rect 255668 296940 437612 296996
rect 437668 296940 437678 296996
rect 260082 296828 260092 296884
rect 260148 296828 443996 296884
rect 444052 296828 444062 296884
rect 316642 296716 316652 296772
rect 316708 296716 405244 296772
rect 405300 296716 405310 296772
rect 312498 296604 312508 296660
rect 312564 296604 413980 296660
rect 414036 296604 414046 296660
rect 417778 296604 417788 296660
rect 417844 296604 438060 296660
rect 438116 296604 438126 296660
rect 314962 296492 314972 296548
rect 315028 296492 443212 296548
rect 443268 296492 443278 296548
rect 424498 294812 424508 294868
rect 424564 294812 441308 294868
rect 441364 294812 441374 294868
rect 149912 293580 172620 293636
rect 172676 293580 172686 293636
rect 438386 293580 438396 293636
rect 438452 293580 444136 293636
rect 301522 291452 301532 291508
rect 301588 291452 312508 291508
rect 312564 291452 312574 291508
rect -960 290836 480 291032
rect -960 290808 3500 290836
rect 392 290780 3500 290808
rect 3556 290780 3566 290836
rect 149912 289996 167468 290052
rect 167524 289996 167534 290052
rect 440850 289996 440860 290052
rect 440916 289996 444136 290052
rect 167682 288988 167692 289044
rect 167748 288988 171052 289044
rect 171108 288988 171118 289044
rect 149912 286412 161196 286468
rect 161252 286412 161262 286468
rect 420690 286412 420700 286468
rect 420756 286412 444136 286468
rect 420130 285628 420140 285684
rect 420196 285628 420476 285684
rect 420532 285628 420542 285684
rect 595560 284676 597000 284872
rect 587122 284620 587132 284676
rect 587188 284648 597000 284676
rect 587188 284620 595672 284648
rect 149912 282828 167580 282884
rect 167636 282828 167646 282884
rect 419794 282828 419804 282884
rect 419860 282828 444136 282884
rect 311154 280588 311164 280644
rect 311220 280588 316652 280644
rect 316708 280588 316718 280644
rect 149912 279244 169260 279300
rect 169316 279244 169326 279300
rect 434914 279244 434924 279300
rect 434980 279244 444136 279300
rect -960 276724 480 276920
rect -960 276696 2492 276724
rect 392 276668 2492 276696
rect 2548 276668 2558 276724
rect 149912 275660 166124 275716
rect 166180 275660 166190 275716
rect 424610 275660 424620 275716
rect 424676 275660 444136 275716
rect 297378 273868 297388 273924
rect 297444 273868 301532 273924
rect 301588 273868 301598 273924
rect 149912 272076 157724 272132
rect 157780 272076 157790 272132
rect 442530 272076 442540 272132
rect 442596 272076 444136 272132
rect 595560 271460 597000 271656
rect 587346 271404 587356 271460
rect 587412 271432 597000 271460
rect 587412 271404 595672 271432
rect 300738 271292 300748 271348
rect 300804 271292 311164 271348
rect 311220 271292 311230 271348
rect 291442 268716 291452 268772
rect 291508 268716 300748 268772
rect 300804 268716 300814 268772
rect 291666 268604 291676 268660
rect 291732 268604 297388 268660
rect 297444 268604 297454 268660
rect 149912 268492 173180 268548
rect 173236 268492 173246 268548
rect 419682 268492 419692 268548
rect 419748 268492 444136 268548
rect 153906 265468 153916 265524
rect 153972 265468 161980 265524
rect 162036 265468 162046 265524
rect 149912 264908 167692 264964
rect 167748 264908 167758 264964
rect 431218 264908 431228 264964
rect 431284 264908 444136 264964
rect -960 262612 480 262808
rect -960 262584 4172 262612
rect 392 262556 4172 262584
rect 4228 262556 4238 262612
rect 149912 261324 154476 261380
rect 154532 261324 154542 261380
rect 441186 261324 441196 261380
rect 441252 261324 444136 261380
rect 420018 258636 420028 258692
rect 420084 258636 420588 258692
rect 420644 258636 420654 258692
rect 595560 258244 597000 258440
rect 587122 258188 587132 258244
rect 587188 258216 597000 258244
rect 587188 258188 595672 258216
rect 149912 257740 158508 257796
rect 158564 257740 158574 257796
rect 421586 257740 421596 257796
rect 421652 257740 444136 257796
rect 160514 257068 160524 257124
rect 160580 257068 162428 257124
rect 162484 257068 162494 257124
rect 149912 254156 150892 254212
rect 150948 254156 150958 254212
rect 436594 254156 436604 254212
rect 436660 254156 444136 254212
rect 285618 251916 285628 251972
rect 285684 251916 291676 251972
rect 291732 251916 291742 251972
rect 149912 250572 172508 250628
rect 172564 250572 172574 250628
rect 433234 250572 433244 250628
rect 433300 250572 444136 250628
rect 286402 250236 286412 250292
rect 286468 250236 291452 250292
rect 291508 250236 291518 250292
rect -960 248500 480 248696
rect 438834 248556 438844 248612
rect 438900 248556 441196 248612
rect 441252 248556 441262 248612
rect -960 248472 9884 248500
rect 392 248444 9884 248472
rect 9940 248444 9950 248500
rect 149912 246988 156156 247044
rect 156212 246988 156222 247044
rect 441746 246988 441756 247044
rect 441812 246988 444136 247044
rect 279010 245196 279020 245252
rect 279076 245196 285628 245252
rect 285684 245196 285694 245252
rect 595560 245028 597000 245224
rect 590482 244972 590492 245028
rect 590548 245000 597000 245028
rect 590548 244972 595672 245000
rect 172386 243628 172396 243684
rect 172452 243628 174188 243684
rect 174244 243628 174254 243684
rect 149912 243404 158620 243460
rect 158676 243404 158686 243460
rect 429314 243404 429324 243460
rect 429380 243404 444136 243460
rect 149912 239820 171388 239876
rect 171444 239820 171454 239876
rect 429202 239820 429212 239876
rect 429268 239820 444136 239876
rect 272962 236796 272972 236852
rect 273028 236796 279020 236852
rect 279076 236796 279086 236852
rect 149912 236236 170828 236292
rect 170884 236236 170894 236292
rect 427858 236236 427868 236292
rect 427924 236236 444136 236292
rect -960 234388 480 234584
rect -960 234360 4284 234388
rect 392 234332 4284 234360
rect 4340 234332 4350 234388
rect 438274 233436 438284 233492
rect 438340 233436 441756 233492
rect 441812 233436 441822 233492
rect 149912 232652 162540 232708
rect 162596 232652 162606 232708
rect 441522 232652 441532 232708
rect 441588 232652 444136 232708
rect 595560 231924 597000 232008
rect 590706 231868 590716 231924
rect 590772 231868 597000 231924
rect 595560 231784 597000 231868
rect 274642 230972 274652 231028
rect 274708 230972 286412 231028
rect 286468 230972 286478 231028
rect 160402 230188 160412 230244
rect 160468 230188 162652 230244
rect 162708 230188 162718 230244
rect 149912 229068 152348 229124
rect 152404 229068 152414 229124
rect 443314 229068 443324 229124
rect 443380 229068 444136 229124
rect 149912 225484 169148 225540
rect 169204 225484 169214 225540
rect 438946 225484 438956 225540
rect 439012 225484 444136 225540
rect 149912 221900 169036 221956
rect 169092 221900 169102 221956
rect 426402 221900 426412 221956
rect 426468 221900 444136 221956
rect -960 220276 480 220472
rect -960 220248 7756 220276
rect 392 220220 7756 220248
rect 7812 220220 7822 220276
rect 595560 218596 597000 218792
rect 587570 218540 587580 218596
rect 587636 218568 597000 218596
rect 587636 218540 595672 218568
rect 273074 218428 273084 218484
rect 273140 218428 274652 218484
rect 274708 218428 274718 218484
rect 149912 218316 154364 218372
rect 154420 218316 154430 218372
rect 441634 218316 441644 218372
rect 441700 218316 444136 218372
rect 149912 214732 165676 214788
rect 165732 214732 165742 214788
rect 433122 214732 433132 214788
rect 433188 214732 444136 214788
rect 149912 211148 173740 211204
rect 173796 211148 173806 211204
rect 438162 211148 438172 211204
rect 438228 211148 444136 211204
rect 149912 207564 173964 207620
rect 174020 207564 174030 207620
rect 426290 207564 426300 207620
rect 426356 207564 444136 207620
rect -960 206164 480 206360
rect -960 206136 7980 206164
rect 392 206108 7980 206136
rect 8036 206108 8046 206164
rect 595560 205380 597000 205576
rect 590594 205324 590604 205380
rect 590660 205352 597000 205380
rect 590660 205324 595672 205352
rect 434802 204988 434812 205044
rect 434868 204988 441532 205044
rect 441588 204988 441598 205044
rect 149912 203980 170604 204036
rect 170660 203980 170670 204036
rect 436706 203980 436716 204036
rect 436772 203980 444136 204036
rect 149912 200396 161084 200452
rect 161140 200396 161150 200452
rect 431106 200396 431116 200452
rect 431172 200396 444136 200452
rect 149912 196812 172396 196868
rect 172452 196812 172462 196868
rect 424386 196812 424396 196868
rect 424452 196812 444136 196868
rect 149912 193228 156044 193284
rect 156100 193228 156110 193284
rect 427746 193228 427756 193284
rect 427812 193228 444136 193284
rect -960 192052 480 192248
rect 595560 192164 597000 192360
rect 590818 192108 590828 192164
rect 590884 192136 597000 192164
rect 590884 192108 595672 192136
rect -960 192024 6188 192052
rect 392 191996 6188 192024
rect 6244 191996 6254 192052
rect 149912 189644 154252 189700
rect 154308 189644 154318 189700
rect 423266 189644 423276 189700
rect 423332 189644 444136 189700
rect 149912 186060 164108 186116
rect 164164 186060 164174 186116
rect 441522 186060 441532 186116
rect 441588 186060 444136 186116
rect 149912 182476 151004 182532
rect 151060 182476 151070 182532
rect 439058 182476 439068 182532
rect 439124 182476 444136 182532
rect 595560 178948 597000 179144
rect 149912 178892 155932 178948
rect 155988 178892 155998 178948
rect 424274 178892 424284 178948
rect 424340 178892 444136 178948
rect 587234 178892 587244 178948
rect 587300 178920 597000 178948
rect 587300 178892 595672 178920
rect -960 177940 480 178136
rect -960 177912 4396 177940
rect 392 177884 4396 177912
rect 4452 177884 4462 177940
rect 149912 175308 165564 175364
rect 165620 175308 165630 175364
rect 423154 175308 423164 175364
rect 423220 175308 444136 175364
rect 421474 173852 421484 173908
rect 421540 173852 441532 173908
rect 441588 173852 441598 173908
rect 149912 171724 160860 171780
rect 160916 171724 160926 171780
rect 441410 171724 441420 171780
rect 441476 171724 444136 171780
rect 419570 170492 419580 170548
rect 419636 170492 441420 170548
rect 441476 170492 441486 170548
rect 149912 168140 157612 168196
rect 157668 168140 157678 168196
rect 426178 168140 426188 168196
rect 426244 168140 444136 168196
rect 595560 165732 597000 165928
rect 590818 165676 590828 165732
rect 590884 165704 597000 165732
rect 590884 165676 595672 165704
rect 149912 164556 155820 164612
rect 155876 164556 155886 164612
rect 433010 164556 433020 164612
rect 433076 164556 444136 164612
rect -960 163828 480 164024
rect -960 163800 9436 163828
rect 392 163772 9436 163800
rect 9492 163772 9502 163828
rect 156034 163772 156044 163828
rect 156100 163772 170940 163828
rect 170996 163772 171006 163828
rect 149912 160972 154140 161028
rect 154196 160972 154206 161028
rect 423042 160972 423052 161028
rect 423108 160972 444136 161028
rect 154354 160412 154364 160468
rect 154420 160412 167356 160468
rect 167412 160412 167422 160468
rect 154130 157948 154140 158004
rect 154196 157948 160972 158004
rect 161028 157948 161038 158004
rect 149912 157388 174076 157444
rect 174132 157388 174142 157444
rect 441522 157388 441532 157444
rect 441588 157388 444136 157444
rect 149912 153804 157500 153860
rect 157556 153804 157566 153860
rect 432898 153804 432908 153860
rect 432964 153804 444136 153860
rect 595560 152516 597000 152712
rect 590930 152460 590940 152516
rect 590996 152488 597000 152516
rect 590996 152460 595672 152488
rect 149912 150220 155708 150276
rect 155764 150220 155774 150276
rect 430994 150220 431004 150276
rect 431060 150220 444136 150276
rect -960 149716 480 149912
rect -960 149688 4508 149716
rect 392 149660 4508 149688
rect 4564 149660 4574 149716
rect 149912 146636 154364 146692
rect 154420 146636 154430 146692
rect 441746 146636 441756 146692
rect 441812 146636 444136 146692
rect 149912 143052 160748 143108
rect 160804 143052 160814 143108
rect 421362 143052 421372 143108
rect 421428 143052 444136 143108
rect 149912 139468 157388 139524
rect 157444 139468 157454 139524
rect 419458 139468 419468 139524
rect 419524 139468 444136 139524
rect 595560 139300 597000 139496
rect 587794 139244 587804 139300
rect 587860 139272 597000 139300
rect 587860 139244 595672 139272
rect 149912 135884 155484 135940
rect 155540 135884 155550 135940
rect 434690 135884 434700 135940
rect 434756 135884 444136 135940
rect -960 135604 480 135800
rect -960 135576 4620 135604
rect 392 135548 4620 135576
rect 4676 135548 4686 135604
rect 154242 132412 154252 132468
rect 154308 132412 158844 132468
rect 158900 132412 158910 132468
rect 149912 132300 154028 132356
rect 154084 132300 154094 132356
rect 422930 132300 422940 132356
rect 422996 132300 444136 132356
rect 149912 128716 154252 128772
rect 154308 128716 154318 128772
rect 421250 128716 421260 128772
rect 421316 128716 444136 128772
rect 595560 126084 597000 126280
rect 591042 126028 591052 126084
rect 591108 126056 597000 126084
rect 591108 126028 595672 126056
rect 149912 125132 157276 125188
rect 157332 125132 157342 125188
rect 157490 125132 157500 125188
rect 157556 125132 170716 125188
rect 170772 125132 170782 125188
rect 434578 125132 434588 125188
rect 434644 125132 444136 125188
rect 154466 123452 154476 123508
rect 154532 123452 168924 123508
rect 168980 123452 168990 123508
rect -960 121492 480 121688
rect 149912 121548 167244 121604
rect 167300 121548 167310 121604
rect 436482 121548 436492 121604
rect 436548 121548 444136 121604
rect -960 121464 8204 121492
rect 392 121436 8204 121464
rect 8260 121436 8270 121492
rect 422706 120092 422716 120148
rect 422772 120092 440188 120148
rect 440244 120092 440254 120148
rect 149912 117964 154476 118020
rect 154532 117964 154542 118020
rect 440178 117964 440188 118020
rect 440244 117964 444136 118020
rect 149912 114380 160636 114436
rect 160692 114380 160702 114436
rect 441298 114380 441308 114436
rect 441364 114380 444136 114436
rect 595560 112868 597000 113064
rect 590482 112812 590492 112868
rect 590548 112840 597000 112868
rect 590548 112812 595672 112840
rect 151106 112588 151116 112644
rect 151172 112588 152908 112644
rect 152964 112588 152974 112644
rect 149912 110796 157164 110852
rect 157220 110796 157230 110852
rect 419346 110796 419356 110852
rect 419412 110796 444136 110852
rect -960 107380 480 107576
rect -960 107352 7644 107380
rect 392 107324 7644 107352
rect 7700 107324 7710 107380
rect 149912 107212 173068 107268
rect 173124 107212 173134 107268
rect 427634 107212 427644 107268
rect 427700 107212 444136 107268
rect 174066 105196 174076 105252
rect 174132 105196 174636 105252
rect 174692 105196 174702 105252
rect 422818 104972 422828 105028
rect 422884 104972 440188 105028
rect 440244 104972 440254 105028
rect 149912 103628 162428 103684
rect 162484 103628 162494 103684
rect 422594 103628 422604 103684
rect 422660 103628 444136 103684
rect 191090 101948 191100 102004
rect 191156 101948 281372 102004
rect 281428 101948 281438 102004
rect 183026 101836 183036 101892
rect 183092 101836 278460 101892
rect 278516 101836 278526 101892
rect 181010 101724 181020 101780
rect 181076 101724 277116 101780
rect 277172 101724 277182 101780
rect 178322 101612 178332 101668
rect 178388 101612 275324 101668
rect 275380 101612 275390 101668
rect 199826 101500 199836 101556
rect 199892 101500 289660 101556
rect 289716 101500 289726 101556
rect 218642 101388 218652 101444
rect 218708 101388 302204 101444
rect 302260 101388 302270 101444
rect 266242 100828 266252 100884
rect 266308 100828 439740 100884
rect 439796 100828 439806 100884
rect 246194 100604 246204 100660
rect 246260 100604 442876 100660
rect 442932 100604 442942 100660
rect 234322 100492 234332 100548
rect 234388 100492 275772 100548
rect 275828 100492 275838 100548
rect 203858 100380 203868 100436
rect 203924 100380 292348 100436
rect 292404 100380 292414 100436
rect 192434 100268 192444 100324
rect 192500 100268 285740 100324
rect 285796 100268 285806 100324
rect 174962 100156 174972 100212
rect 175028 100156 277228 100212
rect 277284 100156 277294 100212
rect 149912 100044 153804 100100
rect 153860 100044 153870 100100
rect 440178 100044 440188 100100
rect 440244 100044 444136 100100
rect 244850 99932 244860 99988
rect 244916 99932 443100 99988
rect 443156 99932 443166 99988
rect 595560 99652 597000 99848
rect 587458 99596 587468 99652
rect 587524 99624 597000 99652
rect 587524 99596 595672 99624
rect 174738 99484 174748 99540
rect 174804 99484 179676 99540
rect 179732 99484 179742 99540
rect 173842 99036 173852 99092
rect 173908 99036 177772 99092
rect 177828 99036 177838 99092
rect 205874 98812 205884 98868
rect 205940 98812 293692 98868
rect 293748 98812 293758 98868
rect 200498 98700 200508 98756
rect 200564 98700 290108 98756
rect 290164 98700 290174 98756
rect 188402 98588 188412 98644
rect 188468 98588 282044 98644
rect 282100 98588 282110 98644
rect 180562 98476 180572 98532
rect 180628 98476 274876 98532
rect 274932 98476 274942 98532
rect 185714 98364 185724 98420
rect 185780 98364 280252 98420
rect 280308 98364 280318 98420
rect 235442 98252 235452 98308
rect 235508 98252 439964 98308
rect 440020 98252 440030 98308
rect 266466 97692 266476 97748
rect 266532 97692 443212 97748
rect 443268 97692 443278 97748
rect 266242 97580 266252 97636
rect 266308 97580 444108 97636
rect 444164 97580 444174 97636
rect 248882 97468 248892 97524
rect 248948 97468 442876 97524
rect 442932 97468 442942 97524
rect 209906 97020 209916 97076
rect 209972 97020 296380 97076
rect 296436 97020 296446 97076
rect 195794 96908 195804 96964
rect 195860 96908 283052 96964
rect 283108 96908 283118 96964
rect 189074 96796 189084 96852
rect 189140 96796 278348 96852
rect 278404 96796 278414 96852
rect 177762 96684 177772 96740
rect 177828 96684 221340 96740
rect 221396 96684 221406 96740
rect 245522 96684 245532 96740
rect 245588 96684 442988 96740
rect 443044 96684 443054 96740
rect 153794 96572 153804 96628
rect 153860 96572 158732 96628
rect 158788 96572 158798 96628
rect 179666 96572 179676 96628
rect 179732 96572 223356 96628
rect 223412 96572 223422 96628
rect 242834 96572 242844 96628
rect 242900 96572 442764 96628
rect 442820 96572 442830 96628
rect 149912 96460 152908 96516
rect 152964 96460 152974 96516
rect 268146 96460 268156 96516
rect 268212 96460 273084 96516
rect 273140 96460 273150 96516
rect 421026 96460 421036 96516
rect 421092 96460 444136 96516
rect 269602 96012 269612 96068
rect 269668 96012 286412 96068
rect 286468 96012 286478 96068
rect 258290 95900 258300 95956
rect 258356 95900 431004 95956
rect 431060 95900 431070 95956
rect 248210 95788 248220 95844
rect 248276 95788 432684 95844
rect 432740 95788 432750 95844
rect 211250 95228 211260 95284
rect 211316 95228 297276 95284
rect 297332 95228 297342 95284
rect 183698 95116 183708 95172
rect 183764 95116 278908 95172
rect 278964 95116 278974 95172
rect 219986 95004 219996 95060
rect 220052 95004 319004 95060
rect 319060 95004 319070 95060
rect 177202 94892 177212 94948
rect 177268 94892 273532 94948
rect 273588 94892 273598 94948
rect 309138 94892 309148 94948
rect 309204 94892 419132 94948
rect 419188 94892 419198 94948
rect 256274 94556 256284 94612
rect 256340 94556 432796 94612
rect 432852 94556 432862 94612
rect 266354 94444 266364 94500
rect 266420 94444 443436 94500
rect 443492 94444 443502 94500
rect 260978 94332 260988 94388
rect 261044 94332 442764 94388
rect 442820 94332 442830 94388
rect 257618 94220 257628 94276
rect 257684 94220 439404 94276
rect 439460 94220 439470 94276
rect 247538 94108 247548 94164
rect 247604 94108 432572 94164
rect 432628 94108 432638 94164
rect 273970 93996 273980 94052
rect 274036 93996 442652 94052
rect 442708 93996 442718 94052
rect 209234 93660 209244 93716
rect 209300 93660 285292 93716
rect 285348 93660 285358 93716
rect 207890 93548 207900 93604
rect 207956 93548 295036 93604
rect 295092 93548 295102 93604
rect -960 93268 480 93464
rect 181682 93436 181692 93492
rect 181748 93436 272972 93492
rect 273028 93436 273038 93492
rect 273746 93436 273756 93492
rect 273812 93436 309148 93492
rect 309204 93436 309214 93492
rect 173618 93324 173628 93380
rect 173684 93324 273868 93380
rect 273924 93324 273934 93380
rect 311602 93324 311612 93380
rect 311668 93324 426860 93380
rect 426916 93324 426926 93380
rect -960 93240 8988 93268
rect 392 93212 8988 93240
rect 9044 93212 9054 93268
rect 243506 93212 243516 93268
rect 243572 93212 435932 93268
rect 435988 93212 435998 93268
rect 149912 92876 157052 92932
rect 157108 92876 157118 92932
rect 419234 92876 419244 92932
rect 419300 92876 444136 92932
rect 270610 92764 270620 92820
rect 270676 92764 428764 92820
rect 428820 92764 428830 92820
rect 260306 92652 260316 92708
rect 260372 92652 431116 92708
rect 431172 92652 431182 92708
rect 250226 92540 250236 92596
rect 250292 92540 432908 92596
rect 432964 92540 432974 92596
rect 252242 92428 252252 92484
rect 252308 92428 437724 92484
rect 437780 92428 437790 92484
rect 201170 92092 201180 92148
rect 201236 92092 290556 92148
rect 290612 92092 290622 92148
rect 195682 91980 195692 92036
rect 195748 91980 285180 92036
rect 285236 91980 285246 92036
rect 187282 91868 187292 91924
rect 187348 91868 279804 91924
rect 279860 91868 279870 91924
rect 184370 91756 184380 91812
rect 184436 91756 279356 91812
rect 279412 91756 279422 91812
rect 182354 91644 182364 91700
rect 182420 91644 278012 91700
rect 278068 91644 278078 91700
rect 318434 91644 318444 91700
rect 318500 91644 420700 91700
rect 420756 91644 420766 91700
rect 154466 91532 154476 91588
rect 154532 91532 172284 91588
rect 172340 91532 172350 91588
rect 179666 91532 179676 91588
rect 179732 91532 276220 91588
rect 276276 91532 276286 91588
rect 315074 91532 315084 91588
rect 315140 91532 426972 91588
rect 427028 91532 427038 91588
rect 271282 91084 271292 91140
rect 271348 91084 298956 91140
rect 299012 91084 299022 91140
rect 276322 90972 276332 91028
rect 276388 90972 429212 91028
rect 429268 90972 429278 91028
rect 266690 90860 266700 90916
rect 266756 90860 439292 90916
rect 439348 90860 439358 90916
rect 255602 90748 255612 90804
rect 255668 90748 435932 90804
rect 435988 90748 435998 90804
rect 238578 90636 238588 90692
rect 238644 90636 289212 90692
rect 289268 90636 289278 90692
rect 207218 90524 207228 90580
rect 207284 90524 294588 90580
rect 294644 90524 294654 90580
rect 205202 90412 205212 90468
rect 205268 90412 293244 90468
rect 293300 90412 293310 90468
rect 203186 90300 203196 90356
rect 203252 90300 291900 90356
rect 291956 90300 291966 90356
rect 318658 90300 318668 90356
rect 318724 90300 422044 90356
rect 422100 90300 422110 90356
rect 198146 90188 198156 90244
rect 198212 90188 287420 90244
rect 287476 90188 287486 90244
rect 318322 90188 318332 90244
rect 318388 90188 425068 90244
rect 425124 90188 425134 90244
rect 198482 90076 198492 90132
rect 198548 90076 288764 90132
rect 288820 90076 288830 90132
rect 315074 90076 315084 90132
rect 315140 90076 443548 90132
rect 443604 90076 443614 90132
rect 192658 89964 192668 90020
rect 192724 89964 283388 90020
rect 283444 89964 283454 90020
rect 311826 89964 311836 90020
rect 311892 89964 442988 90020
rect 443044 89964 443054 90020
rect 155474 89852 155484 89908
rect 155540 89852 170492 89908
rect 170548 89852 170558 89908
rect 186386 89852 186396 89908
rect 186452 89852 280700 89908
rect 280756 89852 280766 89908
rect 286402 89852 286412 89908
rect 286468 89852 421596 89908
rect 421652 89852 421662 89908
rect 149912 89292 154476 89348
rect 154532 89292 154542 89348
rect 425954 89292 425964 89348
rect 426020 89292 444136 89348
rect 269602 89068 269612 89124
rect 269668 89068 429660 89124
rect 429716 89068 429726 89124
rect 273298 88508 273308 88564
rect 273364 88508 442652 88564
rect 442708 88508 442718 88564
rect 216738 88396 216748 88452
rect 216804 88396 295484 88452
rect 295540 88396 295550 88452
rect 210578 88284 210588 88340
rect 210644 88284 296828 88340
rect 296884 88284 296894 88340
rect 195122 88172 195132 88228
rect 195188 88172 284956 88228
rect 285012 88172 285022 88228
rect 295586 88060 295596 88116
rect 295652 88060 351036 88116
rect 351092 88060 351102 88116
rect 269714 87948 269724 88004
rect 269780 87948 315644 88004
rect 315700 87948 315710 88004
rect 317426 87948 317436 88004
rect 317492 87948 429660 88004
rect 429716 87948 429726 88004
rect 272962 87836 272972 87892
rect 273028 87836 429436 87892
rect 429492 87836 429502 87892
rect 265234 87724 265244 87780
rect 265300 87724 421932 87780
rect 421988 87724 421998 87780
rect 270274 87612 270284 87668
rect 270340 87612 432684 87668
rect 432740 87612 432750 87668
rect 270610 87500 270620 87556
rect 270676 87500 436044 87556
rect 436100 87500 436110 87556
rect 287298 87388 287308 87444
rect 287364 87388 299068 87444
rect 299124 87388 299134 87444
rect 421586 87276 421596 87332
rect 421652 87276 430332 87332
rect 430388 87276 430398 87332
rect 224690 87052 224700 87108
rect 224756 87052 273756 87108
rect 273812 87052 273822 87108
rect 315186 87052 315196 87108
rect 315252 87052 421484 87108
rect 421540 87052 421550 87108
rect 237682 86940 237692 86996
rect 237748 86940 287868 86996
rect 287924 86940 287934 86996
rect 318546 86940 318556 86996
rect 318612 86940 421036 86996
rect 421092 86940 421102 86996
rect 212594 86828 212604 86884
rect 212660 86828 298172 86884
rect 298228 86828 298238 86884
rect 318882 86828 318892 86884
rect 318948 86828 421708 86884
rect 421764 86828 421774 86884
rect 193778 86716 193788 86772
rect 193844 86716 284732 86772
rect 284788 86716 284798 86772
rect 318322 86716 318332 86772
rect 318388 86716 421820 86772
rect 421876 86716 421886 86772
rect 191762 86604 191772 86660
rect 191828 86604 284284 86660
rect 284340 86604 284350 86660
rect 187730 86492 187740 86548
rect 187796 86492 281596 86548
rect 281652 86492 281662 86548
rect 314962 86492 314972 86548
rect 315028 86492 422268 86548
rect 422324 86492 422334 86548
rect 426066 86492 426076 86548
rect 426132 86492 441644 86548
rect 441700 86492 441710 86548
rect 595560 86436 597000 86632
rect 591266 86380 591276 86436
rect 591332 86408 597000 86436
rect 591332 86380 595672 86408
rect 273522 86268 273532 86324
rect 273588 86268 443100 86324
rect 443156 86268 443166 86324
rect 292226 86156 292236 86212
rect 292292 86156 319116 86212
rect 319172 86156 319182 86212
rect 269714 86044 269724 86100
rect 269780 86044 340956 86100
rect 341012 86044 341022 86100
rect 414978 86044 414988 86100
rect 415044 86044 431228 86100
rect 431284 86044 431294 86100
rect 273074 85932 273084 85988
rect 273140 85932 436716 85988
rect 436772 85932 436782 85988
rect 268370 85820 268380 85876
rect 268436 85820 436268 85876
rect 436324 85820 436334 85876
rect 149912 85708 153692 85764
rect 153748 85708 153758 85764
rect 268790 85708 268828 85764
rect 268884 85708 268894 85764
rect 283826 85708 283836 85764
rect 283892 85708 299180 85764
rect 299236 85708 299246 85764
rect 441074 85708 441084 85764
rect 441140 85708 444136 85764
rect 266914 85260 266924 85316
rect 266980 85260 276332 85316
rect 276388 85260 276398 85316
rect 299058 85260 299068 85316
rect 299124 85260 315756 85316
rect 315812 85260 315822 85316
rect 174178 85148 174188 85204
rect 174244 85148 222684 85204
rect 222740 85148 222750 85204
rect 225138 85148 225148 85204
rect 225204 85148 301308 85204
rect 301364 85148 301374 85204
rect 215954 85036 215964 85092
rect 216020 85036 300412 85092
rect 300468 85036 300478 85092
rect 420802 85036 420812 85092
rect 420868 85036 441532 85092
rect 441588 85036 441598 85092
rect 215282 84924 215292 84980
rect 215348 84924 299964 84980
rect 300020 84924 300030 84980
rect 315634 84924 315644 84980
rect 315700 84924 429884 84980
rect 429940 84924 429950 84980
rect 154242 84812 154252 84868
rect 154308 84812 172172 84868
rect 172228 84812 172238 84868
rect 211922 84812 211932 84868
rect 211988 84812 297724 84868
rect 297780 84812 297790 84868
rect 298946 84812 298956 84868
rect 299012 84812 425180 84868
rect 425236 84812 425246 84868
rect 317314 84588 317324 84644
rect 317380 84588 429324 84644
rect 429380 84588 429390 84644
rect 270610 84476 270620 84532
rect 270676 84476 314972 84532
rect 315028 84476 315038 84532
rect 317426 84476 317436 84532
rect 317492 84476 436156 84532
rect 436212 84476 436222 84532
rect 282146 84364 282156 84420
rect 282212 84364 428988 84420
rect 429044 84364 429054 84420
rect 269826 84252 269836 84308
rect 269892 84252 422828 84308
rect 422884 84252 422894 84308
rect 270274 84140 270284 84196
rect 270340 84140 425740 84196
rect 425796 84140 425806 84196
rect 270834 84028 270844 84084
rect 270900 84028 443324 84084
rect 443380 84028 443390 84084
rect 271058 83916 271068 83972
rect 271124 83916 287308 83972
rect 287364 83916 287374 83972
rect 319106 83916 319116 83972
rect 319172 83916 414988 83972
rect 415044 83916 415054 83972
rect 230178 83804 230188 83860
rect 230244 83804 268156 83860
rect 268212 83804 268222 83860
rect 274642 83804 274652 83860
rect 274708 83804 317324 83860
rect 317380 83804 317390 83860
rect 173954 83692 173964 83748
rect 174020 83692 218428 83748
rect 218484 83692 218494 83748
rect 228610 83692 228620 83748
rect 228676 83692 267932 83748
rect 267988 83692 267998 83748
rect 273186 83692 273196 83748
rect 273252 83692 317436 83748
rect 317492 83692 317502 83748
rect 216626 83580 216636 83636
rect 216692 83580 298284 83636
rect 298340 83580 298350 83636
rect 351026 83580 351036 83636
rect 351092 83580 434028 83636
rect 434084 83580 434094 83636
rect 217970 83468 217980 83524
rect 218036 83468 301756 83524
rect 301812 83468 301822 83524
rect 340946 83468 340956 83524
rect 341012 83468 431452 83524
rect 431508 83468 431518 83524
rect 201842 83356 201852 83412
rect 201908 83356 291004 83412
rect 291060 83356 291070 83412
rect 321682 83356 321692 83412
rect 321748 83356 422156 83412
rect 422212 83356 422222 83412
rect 180338 83244 180348 83300
rect 180404 83244 267932 83300
rect 267988 83244 267998 83300
rect 271170 83244 271180 83300
rect 271236 83244 282156 83300
rect 282212 83244 282222 83300
rect 315746 83244 315756 83300
rect 315812 83244 419132 83300
rect 419188 83244 419198 83300
rect 420914 83244 420924 83300
rect 420980 83244 441308 83300
rect 441364 83244 441374 83300
rect 176978 83132 176988 83188
rect 177044 83132 274428 83188
rect 274484 83132 274494 83188
rect 276658 83132 276668 83188
rect 276724 83132 276734 83188
rect 299170 83132 299180 83188
rect 299236 83132 425068 83188
rect 425124 83132 425134 83188
rect 276668 83076 276724 83132
rect 267922 83020 267932 83076
rect 267988 83020 276724 83076
rect 266578 82684 266588 82740
rect 266644 82684 428204 82740
rect 428260 82684 428270 82740
rect 416658 82572 416668 82628
rect 416724 82572 429548 82628
rect 429604 82572 429614 82628
rect 282146 82460 282156 82516
rect 282212 82460 429100 82516
rect 429156 82460 429166 82516
rect 268902 82348 268940 82404
rect 268996 82348 269006 82404
rect 422818 82236 422828 82292
rect 422884 82236 425628 82292
rect 425684 82236 425694 82292
rect 149912 82124 160412 82180
rect 160468 82124 160478 82180
rect 421138 82124 421148 82180
rect 421204 82124 444136 82180
rect 270162 81788 270172 81844
rect 270228 81788 295596 81844
rect 295652 81788 295662 81844
rect 213266 81676 213276 81732
rect 213332 81676 298620 81732
rect 298676 81676 298686 81732
rect 197810 81564 197820 81620
rect 197876 81564 288316 81620
rect 288372 81564 288382 81620
rect 187058 81452 187068 81508
rect 187124 81452 278124 81508
rect 278180 81452 278190 81508
rect 287186 81452 287196 81508
rect 287252 81452 416668 81508
rect 416724 81452 416734 81508
rect 419122 81452 419132 81508
rect 419188 81452 440412 81508
rect 440468 81452 440478 81508
rect 295586 81228 295596 81284
rect 295652 81228 428316 81284
rect 428372 81228 428382 81284
rect 273634 81116 273644 81172
rect 273700 81116 420812 81172
rect 420868 81116 420878 81172
rect 266578 81004 266588 81060
rect 266644 81004 423836 81060
rect 423892 81004 423902 81060
rect 271282 80892 271292 80948
rect 271348 80892 439516 80948
rect 439572 80892 439582 80948
rect 268258 80780 268268 80836
rect 268324 80780 442428 80836
rect 442484 80780 442494 80836
rect 220658 80668 220668 80724
rect 220724 80668 433020 80724
rect 433076 80668 433086 80724
rect 175634 80556 175644 80612
rect 175700 80556 177212 80612
rect 177268 80556 177278 80612
rect 177650 80556 177660 80612
rect 177716 80556 180572 80612
rect 180628 80556 180638 80612
rect 185042 80556 185052 80612
rect 185108 80556 187292 80612
rect 187348 80556 187358 80612
rect 189494 80556 189532 80612
rect 189588 80556 189598 80612
rect 190418 80556 190428 80612
rect 190484 80556 192668 80612
rect 192724 80556 192734 80612
rect 193106 80556 193116 80612
rect 193172 80556 195692 80612
rect 195748 80556 195758 80612
rect 202486 80556 202524 80612
rect 202580 80556 202590 80612
rect 204838 80556 204876 80612
rect 204932 80556 204942 80612
rect 206518 80556 206556 80612
rect 206612 80556 206622 80612
rect 213910 80556 213948 80612
rect 214004 80556 214014 80612
rect 214806 80556 214844 80612
rect 214900 80556 214910 80612
rect 226566 80556 226604 80612
rect 226660 80556 226670 80612
rect 228358 80556 228396 80612
rect 228452 80556 228462 80612
rect 229926 80556 229964 80612
rect 230020 80556 230030 80612
rect 232054 80556 232092 80612
rect 232148 80556 232158 80612
rect 233398 80556 233436 80612
rect 233492 80556 233502 80612
rect 234098 80556 234108 80612
rect 234164 80556 235116 80612
rect 235172 80556 235182 80612
rect 236114 80556 236124 80612
rect 236180 80556 236796 80612
rect 236852 80556 236862 80612
rect 238438 80556 238476 80612
rect 238532 80556 238542 80612
rect 241798 80556 241836 80612
rect 241892 80556 241902 80612
rect 242162 80556 242172 80612
rect 242228 80556 243516 80612
rect 243572 80556 243582 80612
rect 244178 80556 244188 80612
rect 244244 80556 245196 80612
rect 245252 80556 245262 80612
rect 246838 80556 246876 80612
rect 246932 80556 246942 80612
rect 249526 80556 249564 80612
rect 249620 80556 249630 80612
rect 251878 80556 251916 80612
rect 251972 80556 251982 80612
rect 253446 80556 253484 80612
rect 253540 80556 253550 80612
rect 254258 80556 254268 80612
rect 254324 80556 254716 80612
rect 254772 80556 254782 80612
rect 259606 80556 259644 80612
rect 259700 80556 259710 80612
rect 425058 80556 425068 80612
rect 425124 80556 429436 80612
rect 429492 80556 429502 80612
rect 208562 80444 208572 80500
rect 208628 80444 216748 80500
rect 216804 80444 216814 80500
rect 226034 80444 226044 80500
rect 226100 80444 226716 80500
rect 226772 80444 226782 80500
rect 228722 80444 228732 80500
rect 228788 80444 230076 80500
rect 230132 80444 230142 80500
rect 254454 80444 254492 80500
rect 254548 80444 254558 80500
rect 274082 80444 274092 80500
rect 274148 80444 292236 80500
rect 292292 80444 292302 80500
rect 425170 80444 425180 80500
rect 425236 80444 429996 80500
rect 430052 80444 430062 80500
rect 199154 80332 199164 80388
rect 199220 80332 238588 80388
rect 238644 80332 238654 80388
rect 240818 80332 240828 80388
rect 240884 80332 425852 80388
rect 425908 80332 425918 80388
rect 176306 80220 176316 80276
rect 176372 80220 181468 80276
rect 181524 80220 181534 80276
rect 220052 80220 225148 80276
rect 225204 80220 225214 80276
rect 225362 80220 225372 80276
rect 225428 80220 228620 80276
rect 228676 80220 228686 80276
rect 237458 80220 237468 80276
rect 237524 80220 424396 80276
rect 424452 80220 424462 80276
rect 220052 80164 220108 80220
rect 217298 80108 217308 80164
rect 217364 80108 220108 80164
rect 224018 80108 224028 80164
rect 224084 80108 230188 80164
rect 230244 80108 230254 80164
rect 236786 80108 236796 80164
rect 236852 80108 424172 80164
rect 424228 80108 424238 80164
rect 197138 79996 197148 80052
rect 197204 79996 237692 80052
rect 237748 79996 237758 80052
rect 239474 79996 239484 80052
rect 239540 79996 429212 80052
rect 429268 79996 429278 80052
rect 172162 79884 172172 79940
rect 172228 79884 219324 79940
rect 219380 79884 219390 79940
rect 240146 79884 240156 79940
rect 240212 79884 430892 79940
rect 430948 79884 430958 79940
rect 178994 79772 179004 79828
rect 179060 79772 234332 79828
rect 234388 79772 234398 79828
rect 234742 79772 234780 79828
rect 234836 79772 234846 79828
rect 238802 79772 238812 79828
rect 238868 79772 434252 79828
rect 434308 79772 434318 79828
rect 229954 79660 229964 79716
rect 230020 79660 230076 79716
rect 230132 79660 230142 79716
rect 252886 79660 252924 79716
rect 252980 79660 252990 79716
rect 256918 79660 256956 79716
rect 257012 79660 257022 79716
rect 231382 79548 231420 79604
rect 231476 79548 231486 79604
rect 270498 79548 270508 79604
rect 270564 79548 282156 79604
rect 282212 79548 282222 79604
rect 232726 79436 232764 79492
rect 232820 79436 232830 79492
rect -960 79156 480 79352
rect 230710 79324 230748 79380
rect 230804 79324 230814 79380
rect 408212 79212 434476 79268
rect 434532 79212 434542 79268
rect -960 79128 9660 79156
rect 392 79100 9660 79128
rect 9716 79100 9726 79156
rect 258962 79100 258972 79156
rect 259028 79100 262108 79156
rect 262052 79044 262108 79100
rect 408212 79044 408268 79212
rect 153682 78988 153692 79044
rect 153748 78988 170940 79044
rect 170996 78988 171006 79044
rect 172946 78988 172956 79044
rect 173012 78988 173852 79044
rect 173908 78988 173918 79044
rect 196466 78988 196476 79044
rect 196532 78988 198156 79044
rect 198212 78988 198222 79044
rect 218418 78988 218428 79044
rect 218484 78988 222012 79044
rect 222068 78988 222078 79044
rect 227350 78988 227388 79044
rect 227444 78988 227454 79044
rect 262052 78988 408268 79044
rect 268146 78876 268156 78932
rect 268212 78876 271292 78932
rect 271348 78876 271358 78932
rect 149912 78540 153804 78596
rect 153860 78540 153870 78596
rect 268594 78540 268604 78596
rect 268660 78540 271180 78596
rect 271236 78540 271246 78596
rect 441410 78540 441420 78596
rect 441476 78540 444136 78596
rect 266690 78428 266700 78484
rect 266756 78428 274652 78484
rect 274708 78428 274718 78484
rect 419122 78428 419132 78484
rect 419188 78428 430892 78484
rect 430948 78428 430958 78484
rect 267026 78316 267036 78372
rect 267092 78316 287196 78372
rect 287252 78316 287262 78372
rect 422482 78316 422492 78372
rect 422548 78316 440188 78372
rect 440244 78316 440254 78372
rect 194450 78204 194460 78260
rect 194516 78204 271516 78260
rect 271572 78204 271582 78260
rect 273410 78204 273420 78260
rect 273476 78204 295596 78260
rect 295652 78204 295662 78260
rect 314962 78204 314972 78260
rect 315028 78204 423948 78260
rect 424004 78204 424014 78260
rect 267922 78092 267932 78148
rect 267988 78092 428204 78148
rect 428260 78092 428270 78148
rect 250870 77308 250908 77364
rect 250964 77308 250974 77364
rect 268034 77196 268044 77252
rect 268100 77196 270620 77252
rect 270676 77196 270686 77252
rect 269826 77084 269836 77140
rect 269892 77084 270620 77140
rect 270676 77084 270686 77140
rect 262052 76860 270620 76916
rect 270676 76860 270686 76916
rect 262052 76468 262108 76860
rect 267810 76748 267820 76804
rect 267876 76748 270508 76804
rect 270564 76748 270574 76804
rect 169586 76412 169596 76468
rect 169652 76412 262108 76468
rect 266802 76300 266812 76356
rect 266868 76300 270620 76356
rect 270676 76300 270686 76356
rect 268818 75404 268828 75460
rect 268884 75404 270088 75460
rect 428642 75404 428652 75460
rect 428708 75404 441084 75460
rect 441140 75404 441150 75460
rect 153682 75292 153692 75348
rect 153748 75292 168812 75348
rect 168868 75292 168878 75348
rect 149912 74956 155596 75012
rect 155652 74956 155662 75012
rect 440402 74956 440412 75012
rect 440468 74956 444136 75012
rect 154018 74732 154028 74788
rect 154084 74732 167132 74788
rect 167188 74732 167198 74788
rect 164546 73948 164556 74004
rect 164612 73948 169708 74004
rect 169764 73948 169774 74004
rect 268930 73836 268940 73892
rect 268996 73836 270088 73892
rect 595560 73220 597000 73416
rect 591154 73164 591164 73220
rect 591220 73192 597000 73220
rect 591220 73164 595672 73192
rect 265906 72604 265916 72660
rect 265972 72604 270116 72660
rect 270060 72296 270116 72604
rect 265944 72044 268828 72100
rect 268884 72044 268894 72100
rect 149912 71372 154252 71428
rect 154308 71372 154318 71428
rect 438050 71372 438060 71428
rect 438116 71372 444136 71428
rect 265944 70700 268940 70756
rect 268996 70700 269006 70756
rect 270050 70700 270060 70756
rect 270116 70700 270126 70756
rect 162194 69580 162204 69636
rect 162260 69580 166040 69636
rect 265906 69356 265916 69412
rect 265972 69356 265982 69412
rect 268818 69132 268828 69188
rect 268884 69132 270088 69188
rect 162642 68684 162652 68740
rect 162708 68684 166040 68740
rect 265916 68460 270060 68516
rect 270116 68460 270126 68516
rect 265916 68040 265972 68460
rect 149884 67900 165452 67956
rect 165508 67900 165518 67956
rect 149884 67816 149940 67900
rect 162418 67788 162428 67844
rect 162484 67788 166040 67844
rect 440178 67788 440188 67844
rect 440244 67788 444136 67844
rect 270050 67564 270060 67620
rect 270116 67564 270126 67620
rect 162306 66892 162316 66948
rect 162372 66892 166040 66948
rect 265944 66668 268828 66724
rect 268884 66668 268894 66724
rect 162082 65996 162092 66052
rect 162148 65996 166040 66052
rect 265906 65996 265916 66052
rect 265972 65996 270088 66052
rect 265944 65324 270060 65380
rect 270116 65324 270126 65380
rect -960 65044 480 65240
rect 164210 65100 164220 65156
rect 164276 65100 166040 65156
rect -960 65016 4732 65044
rect 392 64988 4732 65016
rect 4788 64988 4798 65044
rect 149912 64204 153916 64260
rect 153972 64204 153982 64260
rect 164546 64204 164556 64260
rect 164612 64204 166040 64260
rect 265906 63980 265916 64036
rect 265972 63980 265982 64036
rect 270060 63364 270116 64456
rect 441186 64204 441196 64260
rect 441252 64204 444136 64260
rect 164098 63308 164108 63364
rect 164164 63308 166040 63364
rect 265916 63308 270116 63364
rect 265916 62664 265972 63308
rect 164322 62412 164332 62468
rect 164388 62412 166040 62468
rect 270060 62132 270116 62888
rect 265916 62076 270116 62132
rect 163986 61516 163996 61572
rect 164052 61516 166040 61572
rect 265916 61320 265972 62076
rect 270060 60676 270116 61320
rect 436370 61292 436380 61348
rect 436436 61292 441196 61348
rect 441252 61292 441262 61348
rect 149912 60620 160524 60676
rect 160580 60620 160590 60676
rect 163762 60620 163772 60676
rect 163828 60620 166040 60676
rect 265916 60620 270116 60676
rect 440962 60620 440972 60676
rect 441028 60620 444136 60676
rect 166338 60284 166348 60340
rect 166404 60284 166414 60340
rect 166348 59752 166404 60284
rect 265916 59976 265972 60620
rect 595560 60004 597000 60200
rect 590258 59948 590268 60004
rect 590324 59976 597000 60004
rect 590324 59948 595672 59976
rect 270060 59332 270116 59752
rect 265916 59276 270116 59332
rect 152226 58828 152236 58884
rect 152292 58828 166040 58884
rect 265916 58632 265972 59276
rect 163986 57932 163996 57988
rect 164052 57932 166040 57988
rect 270060 57764 270116 58184
rect 265916 57708 270116 57764
rect 166002 57260 166012 57316
rect 166068 57260 166078 57316
rect 265916 57288 265972 57708
rect 149912 57036 154140 57092
rect 154196 57036 154206 57092
rect 166012 57064 166068 57260
rect 441634 57036 441644 57092
rect 441700 57036 444136 57092
rect 265916 56588 270088 56644
rect 162306 56140 162316 56196
rect 162372 56140 166040 56196
rect 265916 55944 265972 56588
rect 163874 55244 163884 55300
rect 163940 55244 166040 55300
rect 265916 55020 270088 55076
rect 265916 54600 265972 55020
rect 166002 54348 166012 54404
rect 166068 54348 166078 54404
rect 152002 53564 152012 53620
rect 152068 53564 161308 53620
rect 161252 53508 161308 53564
rect 149912 53452 154028 53508
rect 154084 53452 154094 53508
rect 161252 53452 166040 53508
rect 265916 53452 270088 53508
rect 441522 53452 441532 53508
rect 441588 53452 444136 53508
rect 265916 53256 265972 53452
rect 165778 52556 165788 52612
rect 165844 52556 166040 52612
rect 265944 51884 270088 51940
rect 152114 51660 152124 51716
rect 152180 51660 166040 51716
rect -960 50932 480 51128
rect -960 50904 4844 50932
rect 392 50876 4844 50904
rect 4900 50876 4910 50932
rect 162194 50764 162204 50820
rect 162260 50764 166040 50820
rect 265916 50372 265972 50568
rect 265916 50316 270088 50372
rect 149912 49868 155372 49924
rect 155428 49868 155438 49924
rect 163762 49868 163772 49924
rect 163828 49868 166040 49924
rect 441186 49868 441196 49924
rect 441252 49868 444136 49924
rect 430882 49532 430892 49588
rect 430948 49532 440972 49588
rect 441028 49532 441038 49588
rect 162082 48972 162092 49028
rect 162148 48972 166040 49028
rect 265916 48804 265972 49224
rect 265916 48748 270088 48804
rect 166226 48076 166236 48132
rect 166292 48076 166302 48132
rect 152226 47852 152236 47908
rect 152292 47852 163660 47908
rect 163716 47852 163726 47908
rect 265916 47572 265972 47880
rect 265916 47516 270116 47572
rect 150770 47180 150780 47236
rect 150836 47180 166040 47236
rect 270060 47208 270116 47516
rect 595560 46788 597000 46984
rect 590034 46732 590044 46788
rect 590100 46760 597000 46788
rect 590100 46732 595672 46760
rect 149912 46284 157500 46340
rect 157556 46284 157566 46340
rect 164546 46284 164556 46340
rect 164612 46284 166040 46340
rect 265916 46116 265972 46536
rect 441298 46284 441308 46340
rect 441364 46284 444136 46340
rect 265916 46060 270116 46116
rect 270060 45640 270116 46060
rect 163650 45388 163660 45444
rect 163716 45388 166040 45444
rect 432786 45276 432796 45332
rect 432852 45276 440188 45332
rect 440244 45276 440254 45332
rect 265916 44660 265972 45192
rect 265916 44604 270116 44660
rect 150546 44492 150556 44548
rect 150612 44492 166040 44548
rect 270060 44072 270116 44604
rect 150322 43596 150332 43652
rect 150388 43596 166040 43652
rect 265916 43204 265972 43848
rect 265916 43148 270116 43204
rect 149912 42700 156044 42756
rect 156100 42700 156110 42756
rect 163762 42700 163772 42756
rect 163828 42700 166040 42756
rect 270060 42504 270116 43148
rect 440962 42700 440972 42756
rect 441028 42700 444136 42756
rect 152002 41804 152012 41860
rect 152068 41804 166040 41860
rect 265916 41748 265972 42504
rect 265916 41692 270116 41748
rect 163986 40908 163996 40964
rect 164052 40908 166040 40964
rect 265916 40516 265972 41160
rect 270060 40936 270116 41692
rect 265916 40460 270116 40516
rect 150322 40012 150332 40068
rect 150388 40012 166040 40068
rect 265944 39788 268828 39844
rect 268884 39788 268894 39844
rect 270060 39368 270116 40460
rect 149912 39116 155484 39172
rect 155540 39116 155550 39172
rect 164546 39116 164556 39172
rect 164612 39116 166040 39172
rect 440178 39116 440188 39172
rect 440244 39116 444136 39172
rect 265944 38444 270060 38500
rect 270116 38444 270126 38500
rect 155362 38220 155372 38276
rect 155428 38220 166040 38276
rect 268818 37772 268828 37828
rect 268884 37772 270088 37828
rect 164434 37324 164444 37380
rect 164500 37324 166040 37380
rect 265906 37100 265916 37156
rect 265972 37100 265982 37156
rect -960 36820 480 37016
rect 3378 36876 3388 36932
rect 3444 36876 4172 36932
rect 4228 36876 4238 36932
rect -960 36792 4956 36820
rect 392 36764 4956 36792
rect 5012 36764 5022 36820
rect 150322 36428 150332 36484
rect 150388 36428 166040 36484
rect 270050 36204 270060 36260
rect 270116 36204 270126 36260
rect 265916 35588 265972 35784
rect 149912 35532 153692 35588
rect 153748 35532 153758 35588
rect 164210 35532 164220 35588
rect 164276 35532 166040 35588
rect 265916 35532 270060 35588
rect 270116 35532 270126 35588
rect 441074 35532 441084 35588
rect 441140 35532 444136 35588
rect 265906 35084 265916 35140
rect 265972 35084 270116 35140
rect 163538 34636 163548 34692
rect 163604 34636 166040 34692
rect 270060 34664 270116 35084
rect 265944 34412 266140 34468
rect 266196 34412 266206 34468
rect 428978 34412 428988 34468
rect 429044 34412 441644 34468
rect 441700 34412 441710 34468
rect 163762 33740 163772 33796
rect 163828 33740 166040 33796
rect 595560 33684 597000 33768
rect 589810 33628 589820 33684
rect 589876 33628 597000 33684
rect 595560 33544 597000 33628
rect 265944 33068 268828 33124
rect 268884 33068 268894 33124
rect 270050 33068 270060 33124
rect 270116 33068 270126 33124
rect 152226 32844 152236 32900
rect 152292 32844 166040 32900
rect 149912 31948 153692 32004
rect 153748 31948 153758 32004
rect 163874 31948 163884 32004
rect 163940 31948 166040 32004
rect 433010 31948 433020 32004
rect 433076 31948 444136 32004
rect 265906 31724 265916 31780
rect 265972 31724 265982 31780
rect 266130 31500 266140 31556
rect 266196 31500 270088 31556
rect 152114 31052 152124 31108
rect 152180 31052 166040 31108
rect 265944 30380 268940 30436
rect 268996 30380 269006 30436
rect 153682 30156 153692 30212
rect 153748 30156 166040 30212
rect 268818 29932 268828 29988
rect 268884 29932 270088 29988
rect 429426 29372 429436 29428
rect 429492 29372 437836 29428
rect 437892 29372 437902 29428
rect 164098 29260 164108 29316
rect 164164 29260 166040 29316
rect 265944 29036 268828 29092
rect 268884 29036 268894 29092
rect 163986 28364 163996 28420
rect 164052 28364 166040 28420
rect 265906 28364 265916 28420
rect 265972 28364 270088 28420
rect 265944 27692 270060 27748
rect 270116 27692 270126 27748
rect 164210 27468 164220 27524
rect 164276 27468 166040 27524
rect 268930 26796 268940 26852
rect 268996 26796 270088 26852
rect 4162 26572 4172 26628
rect 4228 26572 4508 26628
rect 4564 26572 4574 26628
rect 164322 26572 164332 26628
rect 164388 26572 166040 26628
rect 4498 26348 4508 26404
rect 4564 26348 4732 26404
rect 4788 26348 4798 26404
rect 265906 26348 265916 26404
rect 265972 26348 265982 26404
rect 150434 25676 150444 25732
rect 150500 25676 166040 25732
rect 268818 25228 268828 25284
rect 268884 25228 270088 25284
rect 265944 25004 267036 25060
rect 267092 25004 267102 25060
rect 153906 24780 153916 24836
rect 153972 24780 166040 24836
rect 152338 23884 152348 23940
rect 152404 23884 166040 23940
rect 265944 23660 268940 23716
rect 268996 23660 269006 23716
rect 270050 23660 270060 23716
rect 270116 23660 270126 23716
rect 3462 23436 3500 23492
rect 3556 23436 3566 23492
rect 265458 23100 265468 23156
rect 265524 23100 270284 23156
rect 270340 23100 270350 23156
rect 159730 22988 159740 23044
rect 159796 22988 166040 23044
rect -960 22708 480 22904
rect 429986 22764 429996 22820
rect 430052 22764 439964 22820
rect 440020 22764 440030 22820
rect -960 22680 4956 22708
rect 392 22652 4956 22680
rect 5012 22652 5022 22708
rect 429650 22652 429660 22708
rect 429716 22652 440076 22708
rect 440132 22652 440142 22708
rect 265944 22316 268828 22372
rect 268884 22316 268894 22372
rect 149762 22092 149772 22148
rect 149828 22092 166040 22148
rect 265906 22092 265916 22148
rect 265972 22092 270088 22148
rect 4050 20972 4060 21028
rect 4116 20972 155372 21028
rect 155428 20972 155438 21028
rect 265944 20972 270060 21028
rect 270116 20972 270126 21028
rect 439058 20972 439068 21028
rect 439124 20972 591052 21028
rect 591108 20972 591118 21028
rect 438834 20860 438844 20916
rect 438900 20860 590828 20916
rect 590884 20860 590894 20916
rect 438610 20748 438620 20804
rect 438676 20748 590604 20804
rect 590660 20748 590670 20804
rect 443202 20636 443212 20692
rect 443268 20636 591276 20692
rect 591332 20636 591342 20692
rect 267026 20524 267036 20580
rect 267092 20524 270088 20580
rect 595560 20356 597000 20552
rect 591266 20300 591276 20356
rect 591332 20328 597000 20356
rect 591332 20300 595672 20328
rect 7746 20076 7756 20132
rect 7812 20076 164220 20132
rect 164276 20076 164286 20132
rect 430994 20076 431004 20132
rect 431060 20076 590268 20132
rect 590324 20076 590334 20132
rect 7522 19964 7532 20020
rect 7588 19964 163772 20020
rect 163828 19964 163838 20020
rect 431218 19964 431228 20020
rect 431284 19964 589820 20020
rect 589876 19964 589886 20020
rect 8194 19852 8204 19908
rect 8260 19852 164108 19908
rect 164164 19852 164174 19908
rect 432450 19852 432460 19908
rect 432516 19852 590940 19908
rect 590996 19852 591006 19908
rect 7970 19740 7980 19796
rect 8036 19740 163548 19796
rect 163604 19740 163614 19796
rect 433010 19740 433020 19796
rect 433076 19740 590716 19796
rect 590772 19740 590782 19796
rect 9202 19628 9212 19684
rect 9268 19628 163996 19684
rect 164052 19628 164062 19684
rect 265906 19628 265916 19684
rect 265972 19628 265982 19684
rect 434466 19628 434476 19684
rect 434532 19628 590044 19684
rect 590100 19628 590110 19684
rect 9650 19516 9660 19572
rect 9716 19516 164332 19572
rect 164388 19516 164398 19572
rect 432786 19516 432796 19572
rect 432852 19516 587468 19572
rect 587524 19516 587534 19572
rect 9426 19404 9436 19460
rect 9492 19404 163884 19460
rect 163940 19404 163950 19460
rect 437714 19404 437724 19460
rect 437780 19404 587244 19460
rect 587300 19404 587310 19460
rect 4834 19292 4844 19348
rect 4900 19292 152348 19348
rect 152404 19292 152414 19348
rect 442866 19292 442876 19348
rect 442932 19292 590492 19348
rect 590548 19292 590558 19348
rect 4274 19180 4284 19236
rect 4340 19180 150332 19236
rect 150388 19180 150398 19236
rect 440066 19180 440076 19236
rect 440132 19180 464492 19236
rect 464548 19180 464558 19236
rect 268930 18956 268940 19012
rect 268996 18956 270088 19012
rect 164518 18508 164556 18564
rect 164612 18508 164622 18564
rect 265234 18508 265244 18564
rect 265300 18508 269836 18564
rect 269892 18508 269902 18564
rect 6178 18396 6188 18452
rect 6244 18396 163772 18452
rect 163828 18396 163838 18452
rect 256946 18396 256956 18452
rect 257012 18396 268828 18452
rect 268884 18396 268894 18452
rect 431106 18396 431116 18452
rect 431172 18396 591276 18452
rect 591332 18396 591342 18452
rect 4946 18284 4956 18340
rect 5012 18284 159740 18340
rect 159796 18284 159806 18340
rect 164434 18284 164444 18340
rect 164500 18284 164510 18340
rect 268902 18284 268940 18340
rect 268996 18284 269006 18340
rect 433346 18284 433356 18340
rect 433412 18284 590828 18340
rect 590884 18284 590894 18340
rect 8978 18172 8988 18228
rect 9044 18172 164220 18228
rect 164276 18172 164286 18228
rect 164444 18116 164500 18284
rect 432562 18172 432572 18228
rect 432628 18172 587356 18228
rect 587412 18172 587422 18228
rect 9874 18060 9884 18116
rect 9940 18060 164500 18116
rect 433122 18060 433132 18116
rect 433188 18060 587804 18116
rect 587860 18060 587870 18116
rect 4610 17948 4620 18004
rect 4676 17948 153692 18004
rect 153748 17948 153758 18004
rect 252802 17948 252812 18004
rect 252868 17948 265020 18004
rect 265076 17948 265086 18004
rect 432898 17948 432908 18004
rect 432964 17948 587580 18004
rect 587636 17948 587646 18004
rect 4722 17836 4732 17892
rect 4788 17836 153916 17892
rect 153972 17836 153982 17892
rect 241714 17836 241724 17892
rect 241780 17836 266924 17892
rect 266980 17836 266990 17892
rect 435922 17836 435932 17892
rect 435988 17836 590492 17892
rect 590548 17836 590558 17892
rect 4386 17724 4396 17780
rect 4452 17724 152236 17780
rect 152292 17724 152302 17780
rect 222450 17724 222460 17780
rect 222516 17724 252028 17780
rect 252084 17724 252094 17780
rect 439394 17724 439404 17780
rect 439460 17724 591164 17780
rect 591220 17724 591230 17780
rect 3490 17612 3500 17668
rect 3556 17612 150332 17668
rect 150388 17612 150398 17668
rect 222898 17612 222908 17668
rect 222964 17612 256844 17668
rect 256900 17612 256910 17668
rect 429202 17612 429212 17668
rect 429268 17612 438508 17668
rect 438564 17612 438574 17668
rect 440066 17612 440076 17668
rect 440132 17612 587132 17668
rect 587188 17612 587198 17668
rect 228834 17500 228844 17556
rect 228900 17500 269052 17556
rect 269108 17500 269118 17556
rect 437826 17500 437836 17556
rect 437892 17500 460684 17556
rect 460740 17500 460750 17556
rect 223122 17388 223132 17444
rect 223188 17388 265468 17444
rect 265524 17388 265534 17444
rect 268818 17388 268828 17444
rect 268884 17388 270088 17444
rect 223346 17276 223356 17332
rect 223412 17276 269500 17332
rect 269556 17276 269566 17332
rect 219538 17164 219548 17220
rect 219604 17164 269388 17220
rect 269444 17164 269454 17220
rect 216860 17052 268380 17108
rect 268436 17052 268446 17108
rect 216860 16772 216916 17052
rect 217532 16940 243628 16996
rect 217532 16772 217588 16940
rect 243572 16884 243628 16940
rect 262052 16940 270452 16996
rect 262052 16884 262108 16940
rect 219324 16828 219548 16884
rect 219604 16828 219614 16884
rect 221116 16828 222460 16884
rect 222516 16828 222526 16884
rect 222684 16828 222908 16884
rect 222964 16828 222974 16884
rect 223132 16828 223356 16884
rect 223412 16828 223422 16884
rect 225820 16828 228844 16884
rect 228900 16828 228910 16884
rect 240156 16828 241724 16884
rect 241780 16828 241790 16884
rect 243572 16828 262108 16884
rect 265468 16828 268604 16884
rect 268660 16828 268670 16884
rect 219324 16772 219380 16828
rect 221116 16772 221172 16828
rect 222684 16772 222740 16828
rect 223132 16772 223188 16828
rect 225820 16772 225876 16828
rect 240156 16772 240212 16828
rect 4134 16716 4172 16772
rect 4228 16716 4238 16772
rect 216850 16716 216860 16772
rect 216916 16716 216926 16772
rect 217522 16716 217532 16772
rect 217588 16716 217598 16772
rect 219090 16716 219100 16772
rect 219156 16716 219380 16772
rect 221106 16716 221116 16772
rect 221172 16716 221182 16772
rect 222450 16716 222460 16772
rect 222516 16716 222740 16772
rect 222898 16716 222908 16772
rect 222964 16716 223188 16772
rect 225810 16716 225820 16772
rect 225876 16716 225886 16772
rect 226230 16716 226268 16772
rect 226324 16716 226334 16772
rect 230710 16716 230748 16772
rect 230804 16716 230814 16772
rect 231158 16716 231196 16772
rect 231252 16716 231262 16772
rect 236534 16716 236572 16772
rect 236628 16716 236638 16772
rect 239222 16716 239260 16772
rect 239316 16716 239326 16772
rect 239922 16716 239932 16772
rect 239988 16716 240212 16772
rect 240342 16716 240380 16772
rect 240436 16716 240446 16772
rect 240594 16716 240604 16772
rect 240660 16716 240698 16772
rect 243702 16716 243740 16772
rect 243796 16716 243806 16772
rect 245046 16716 245084 16772
rect 245140 16716 245150 16772
rect 7634 16604 7644 16660
rect 7700 16604 163996 16660
rect 164052 16604 164062 16660
rect 223094 16604 223132 16660
rect 223188 16604 223198 16660
rect 238578 16604 238588 16660
rect 238644 16604 241948 16660
rect 242004 16604 242014 16660
rect 4386 16492 4396 16548
rect 4452 16492 152124 16548
rect 152180 16492 152190 16548
rect 4498 16380 4508 16436
rect 4564 16380 150444 16436
rect 150500 16380 150510 16436
rect 265468 16324 265524 16828
rect 270396 16772 270452 16940
rect 270386 16716 270396 16772
rect 270452 16716 270462 16772
rect 442642 16716 442652 16772
rect 442708 16716 487340 16772
rect 487396 16716 487406 16772
rect 439506 16604 439516 16660
rect 439572 16604 491148 16660
rect 491204 16604 491214 16660
rect 436706 16492 436716 16548
rect 436772 16492 514108 16548
rect 514164 16492 514174 16548
rect 436034 16380 436044 16436
rect 436100 16380 525420 16436
rect 525476 16380 525486 16436
rect 2482 16268 2492 16324
rect 2548 16268 164556 16324
rect 164612 16268 164622 16324
rect 245270 16268 245308 16324
rect 245364 16268 245374 16324
rect 249554 16268 249564 16324
rect 249620 16268 265524 16324
rect 436258 16268 436268 16324
rect 436324 16268 538748 16324
rect 538804 16268 538814 16324
rect 216626 16156 216636 16212
rect 216692 16156 231868 16212
rect 248546 16156 248556 16212
rect 248612 16156 269724 16212
rect 269780 16156 269790 16212
rect 443090 16156 443100 16212
rect 443156 16156 565404 16212
rect 565460 16156 565470 16212
rect 231812 16100 231868 16156
rect 114258 16044 114268 16100
rect 114324 16044 197820 16100
rect 197876 16044 197886 16100
rect 200498 16044 200508 16100
rect 200564 16044 200574 16100
rect 217270 16044 217308 16100
rect 217364 16044 217374 16100
rect 219762 16044 219772 16100
rect 219828 16044 220108 16100
rect 226006 16044 226044 16100
rect 226100 16044 226110 16100
rect 231812 16044 266476 16100
rect 266532 16044 266542 16100
rect 436482 16044 436492 16100
rect 436548 16044 567308 16100
rect 567364 16044 567374 16100
rect 200508 15988 200564 16044
rect 136994 15932 137004 15988
rect 137060 15932 200564 15988
rect 220052 15988 220108 16044
rect 220052 15932 269276 15988
rect 269332 15932 269342 15988
rect 439954 15932 439964 15988
rect 440020 15932 578732 15988
rect 578788 15932 578798 15988
rect 148418 15820 148428 15876
rect 148484 15820 201852 15876
rect 201908 15820 201918 15876
rect 215954 15820 215964 15876
rect 216020 15820 260764 15876
rect 260820 15820 260830 15876
rect 270050 15820 270060 15876
rect 270116 15820 270126 15876
rect 439954 15820 439964 15876
rect 440020 15820 447356 15876
rect 447412 15820 447422 15876
rect 226482 15708 226492 15764
rect 226548 15708 269948 15764
rect 270004 15708 270014 15764
rect 215282 15596 215292 15652
rect 215348 15596 255052 15652
rect 255108 15596 255118 15652
rect 214610 15484 214620 15540
rect 214676 15484 249228 15540
rect 249284 15484 249294 15540
rect 226818 15372 226828 15428
rect 226884 15372 247772 15428
rect 247828 15372 247838 15428
rect 253698 15372 253708 15428
rect 253764 15372 269164 15428
rect 269220 15372 269230 15428
rect 142818 15260 142828 15316
rect 142884 15260 201180 15316
rect 201236 15260 201246 15316
rect 230402 15260 230412 15316
rect 230468 15260 265468 15316
rect 265524 15260 265534 15316
rect 117954 15148 117964 15204
rect 118020 15148 198156 15204
rect 198212 15148 198222 15204
rect 227154 15148 227164 15204
rect 227220 15148 270508 15204
rect 270564 15148 270574 15204
rect 220052 15036 253708 15092
rect 253764 15036 253774 15092
rect 256834 15036 256844 15092
rect 256900 15036 265692 15092
rect 265748 15036 265758 15092
rect 438498 15036 438508 15092
rect 438564 15036 441868 15092
rect 441924 15036 441934 15092
rect 219986 14924 219996 14980
rect 220052 14924 220108 15036
rect 221302 14924 221340 14980
rect 221396 14924 221406 14980
rect 222198 14924 222236 14980
rect 222292 14924 222302 14980
rect 243030 14924 243068 14980
rect 243124 14924 243134 14980
rect 244850 14924 244860 14980
rect 244916 14924 266924 14980
rect 266980 14924 266990 14980
rect 144610 14812 144620 14868
rect 144676 14812 201404 14868
rect 201460 14812 201470 14868
rect 432674 14812 432684 14868
rect 432740 14812 508284 14868
rect 508340 14812 508350 14868
rect 133186 14700 133196 14756
rect 133252 14700 200060 14756
rect 200116 14700 200126 14756
rect 429874 14700 429884 14756
rect 429940 14700 519708 14756
rect 519764 14700 519774 14756
rect 106530 14588 106540 14644
rect 106596 14588 196924 14644
rect 196980 14588 196990 14644
rect 233874 14588 233884 14644
rect 233940 14588 244524 14644
rect 244580 14588 244590 14644
rect 252018 14588 252028 14644
rect 252084 14588 268716 14644
rect 268772 14588 268782 14644
rect 429090 14588 429100 14644
rect 429156 14588 529228 14644
rect 529284 14588 529294 14644
rect 69682 14476 69692 14532
rect 69748 14476 192444 14532
rect 192500 14476 192510 14532
rect 218866 14476 218876 14532
rect 218932 14476 270620 14532
rect 270676 14476 270686 14532
rect 437826 14476 437836 14532
rect 437892 14476 546812 14532
rect 546868 14476 546878 14532
rect 4162 14364 4172 14420
rect 4228 14364 149772 14420
rect 149828 14364 149838 14420
rect 167458 14364 167468 14420
rect 167524 14364 204092 14420
rect 204148 14364 204158 14420
rect 228498 14364 228508 14420
rect 228564 14364 269724 14420
rect 269780 14364 269790 14420
rect 432898 14364 432908 14420
rect 432964 14364 569212 14420
rect 569268 14364 569278 14420
rect 42802 14252 42812 14308
rect 42868 14252 189308 14308
rect 189364 14252 189374 14308
rect 215730 14252 215740 14308
rect 215796 14252 258860 14308
rect 258916 14252 258926 14308
rect 265906 14252 265916 14308
rect 265972 14252 270088 14308
rect 429650 14252 429660 14308
rect 429716 14252 576828 14308
rect 576884 14252 576894 14308
rect 268146 14140 268156 14196
rect 268212 14140 268604 14196
rect 268660 14140 268670 14196
rect 233426 13804 233436 13860
rect 233492 13804 253148 13860
rect 253204 13804 253214 13860
rect 104626 13692 104636 13748
rect 104692 13692 196700 13748
rect 196756 13692 196766 13748
rect 240258 13692 240268 13748
rect 240324 13692 269724 13748
rect 269780 13692 269790 13748
rect 87490 13580 87500 13636
rect 87556 13580 191604 13636
rect 230178 13580 230188 13636
rect 230244 13580 270284 13636
rect 270340 13580 270350 13636
rect 53218 13468 53228 13524
rect 53284 13468 188244 13524
rect 188188 13412 188244 13468
rect 191548 13412 191604 13580
rect 218204 13468 264572 13524
rect 264628 13468 264638 13524
rect 218204 13412 218260 13468
rect 186806 13356 186844 13412
rect 186900 13356 186910 13412
rect 187030 13356 187068 13412
rect 187124 13356 187134 13412
rect 188188 13356 190652 13412
rect 190708 13356 190718 13412
rect 191548 13356 194684 13412
rect 194740 13356 194750 13412
rect 207554 13356 207564 13412
rect 207620 13356 208796 13412
rect 208852 13356 208862 13412
rect 209430 13356 209468 13412
rect 209524 13356 209534 13412
rect 209654 13356 209692 13412
rect 209748 13356 209758 13412
rect 209906 13356 209916 13412
rect 209972 13356 210010 13412
rect 210102 13356 210140 13412
rect 210196 13356 210206 13412
rect 216402 13356 216412 13412
rect 216468 13356 218260 13412
rect 218614 13356 218652 13412
rect 218708 13356 218718 13412
rect 224466 13356 224476 13412
rect 224532 13356 230412 13412
rect 230468 13356 230478 13412
rect 236086 13356 236124 13412
rect 236180 13356 236190 13412
rect 241462 13356 241500 13412
rect 241556 13356 241566 13412
rect 243282 13356 243292 13412
rect 243348 13356 243516 13412
rect 243572 13356 243582 13412
rect 245942 13356 245980 13412
rect 246036 13356 246046 13412
rect 265458 13356 265468 13412
rect 265524 13356 267820 13412
rect 267876 13356 267886 13412
rect 268482 13356 268492 13412
rect 268548 13356 269612 13412
rect 269668 13356 269678 13412
rect 270610 13356 270620 13412
rect 270676 13356 270686 13412
rect 442418 13356 442428 13412
rect 442484 13356 458780 13412
rect 458836 13356 458846 13412
rect 270620 13300 270676 13356
rect 154130 13244 154140 13300
rect 154196 13244 202524 13300
rect 202580 13244 202590 13300
rect 205538 13244 205548 13300
rect 205604 13244 208572 13300
rect 208628 13244 208638 13300
rect 217074 13244 217084 13300
rect 217140 13244 230188 13300
rect 230244 13244 230254 13300
rect 235218 13244 235228 13300
rect 235284 13244 243628 13300
rect 249442 13244 249452 13300
rect 249508 13244 268268 13300
rect 268324 13244 268334 13300
rect 268706 13244 268716 13300
rect 268772 13244 270676 13300
rect 434354 13244 434364 13300
rect 434420 13244 472108 13300
rect 472164 13244 472174 13300
rect 243572 13188 243628 13244
rect 116722 13132 116732 13188
rect 116788 13132 188412 13188
rect 188468 13132 188478 13188
rect 190194 13132 190204 13188
rect 190260 13132 190428 13188
rect 190484 13132 190494 13188
rect 193106 13132 193116 13188
rect 193172 13132 193182 13188
rect 220434 13132 220444 13188
rect 220500 13132 226828 13188
rect 226884 13132 226894 13188
rect 234770 13132 234780 13188
rect 234836 13132 239148 13188
rect 239204 13132 239214 13188
rect 243572 13132 266252 13188
rect 266308 13132 266318 13188
rect 268594 13132 268604 13188
rect 268660 13132 270620 13188
rect 270676 13132 270686 13188
rect 436146 13132 436156 13188
rect 436212 13132 481628 13188
rect 481684 13132 481694 13188
rect 193116 13076 193172 13132
rect 92306 13020 92316 13076
rect 92372 13020 185724 13076
rect 185780 13020 185790 13076
rect 186060 13020 193172 13076
rect 194450 13020 194460 13076
rect 194516 13020 194526 13076
rect 243572 13020 268716 13076
rect 268772 13020 268782 13076
rect 270498 13020 270508 13076
rect 270564 13020 270574 13076
rect 442642 13020 442652 13076
rect 442708 13020 493052 13076
rect 493108 13020 493118 13076
rect 81442 12908 81452 12964
rect 81508 12908 185836 12964
rect 185892 12908 185902 12964
rect 186060 12852 186116 13020
rect 194460 12964 194516 13020
rect 243572 12964 243628 13020
rect 270508 12964 270564 13020
rect 186498 12908 186508 12964
rect 186564 12908 191772 12964
rect 191828 12908 191838 12964
rect 191996 12908 194516 12964
rect 221974 12908 222012 12964
rect 222068 12908 222078 12964
rect 236786 12908 236796 12964
rect 236852 12908 240492 12964
rect 240548 12908 240558 12964
rect 240818 12908 240828 12964
rect 240884 12908 243628 12964
rect 243964 12908 266812 12964
rect 266868 12908 266878 12964
rect 268706 12908 268716 12964
rect 268772 12908 270564 12964
rect 443090 12908 443100 12964
rect 443156 12908 498764 12964
rect 498820 12908 498830 12964
rect 191996 12852 192052 12908
rect 74162 12796 74172 12852
rect 74228 12796 186116 12852
rect 186386 12796 186396 12852
rect 186452 12796 192052 12852
rect 194114 12796 194124 12852
rect 194180 12796 207228 12852
rect 207284 12796 207294 12852
rect 211922 12796 211932 12852
rect 211988 12796 226492 12852
rect 226548 12796 226558 12852
rect 227378 12796 227388 12852
rect 227444 12796 241052 12852
rect 241108 12796 241118 12852
rect 242358 12796 242396 12852
rect 242452 12796 242462 12852
rect 243964 12740 244020 12908
rect 244178 12796 244188 12852
rect 244244 12796 270620 12852
rect 270676 12796 270686 12852
rect 443314 12796 443324 12852
rect 443380 12796 504476 12852
rect 504532 12796 504542 12852
rect 54562 12684 54572 12740
rect 54628 12684 190428 12740
rect 190484 12684 190494 12740
rect 190642 12684 190652 12740
rect 190708 12684 204540 12740
rect 204596 12684 204606 12740
rect 212146 12684 212156 12740
rect 212212 12684 228508 12740
rect 228564 12684 228574 12740
rect 231382 12684 231420 12740
rect 231476 12684 231486 12740
rect 232082 12684 232092 12740
rect 232148 12684 234892 12740
rect 234948 12684 234958 12740
rect 239026 12684 239036 12740
rect 239092 12684 244020 12740
rect 249442 12684 249452 12740
rect 249508 12684 270396 12740
rect 270452 12684 270462 12740
rect 436706 12684 436716 12740
rect 436772 12684 510188 12740
rect 510244 12684 510254 12740
rect 37762 12572 37772 12628
rect 37828 12572 188636 12628
rect 188692 12572 188702 12628
rect 192546 12572 192556 12628
rect 192612 12572 207004 12628
rect 207060 12572 207070 12628
rect 220658 12572 220668 12628
rect 220724 12572 269836 12628
rect 269892 12572 269902 12628
rect 428306 12572 428316 12628
rect 428372 12572 435932 12628
rect 435988 12572 435998 12628
rect 442866 12572 442876 12628
rect 442932 12572 584444 12628
rect 584500 12572 584510 12628
rect 185042 12460 185052 12516
rect 185108 12460 186396 12516
rect 186452 12460 186462 12516
rect 192322 12460 192332 12516
rect 192388 12460 194236 12516
rect 194292 12460 194302 12516
rect 220882 12460 220892 12516
rect 220948 12460 240268 12516
rect 240324 12460 240334 12516
rect 240482 12460 240492 12516
rect 240548 12460 249452 12516
rect 249508 12460 249518 12516
rect 179106 12348 179116 12404
rect 179172 12348 199836 12404
rect 199892 12348 199902 12404
rect 224018 12348 224028 12404
rect 224084 12348 225036 12404
rect 225092 12348 225102 12404
rect 225362 12348 225372 12404
rect 225428 12348 226604 12404
rect 226660 12348 226670 12404
rect 232530 12348 232540 12404
rect 232596 12348 235116 12404
rect 235172 12348 235182 12404
rect 237906 12348 237916 12404
rect 237972 12348 238476 12404
rect 238532 12348 238542 12404
rect 239138 12348 239148 12404
rect 239204 12348 242004 12404
rect 242162 12348 242172 12404
rect 242228 12348 243292 12404
rect 243348 12348 243358 12404
rect 244402 12348 244412 12404
rect 244468 12348 245196 12404
rect 245252 12348 245262 12404
rect 241948 12292 242004 12348
rect 184930 12236 184940 12292
rect 184996 12236 185948 12292
rect 186004 12236 186014 12292
rect 186162 12236 186172 12292
rect 186228 12236 186266 12292
rect 186498 12236 186508 12292
rect 186564 12236 187516 12292
rect 187572 12236 187582 12292
rect 188178 12236 188188 12292
rect 188244 12236 189084 12292
rect 189140 12236 189150 12292
rect 190418 12236 190428 12292
rect 190484 12236 190876 12292
rect 190932 12236 190942 12292
rect 191426 12236 191436 12292
rect 191492 12236 192668 12292
rect 192724 12236 192734 12292
rect 193442 12236 193452 12292
rect 193508 12236 195580 12292
rect 195636 12236 195646 12292
rect 197474 12236 197484 12292
rect 197540 12236 199164 12292
rect 199220 12236 199230 12292
rect 204082 12236 204092 12292
rect 204148 12236 205436 12292
rect 205492 12236 205502 12292
rect 223318 12236 223356 12292
rect 223412 12236 223422 12292
rect 224690 12236 224700 12292
rect 224756 12236 224924 12292
rect 224980 12236 224990 12292
rect 226678 12236 226716 12292
rect 226772 12236 226782 12292
rect 228050 12236 228060 12292
rect 228116 12236 228396 12292
rect 228452 12236 228462 12292
rect 229394 12236 229404 12292
rect 229460 12236 230076 12292
rect 230132 12236 230142 12292
rect 231606 12236 231644 12292
rect 231700 12236 231710 12292
rect 232978 12236 232988 12292
rect 233044 12236 237804 12292
rect 237860 12236 237870 12292
rect 238326 12236 238364 12292
rect 238420 12236 238430 12292
rect 240118 12236 240156 12292
rect 240212 12236 240222 12292
rect 241266 12236 241276 12292
rect 241332 12236 241724 12292
rect 241780 12236 241790 12292
rect 241948 12236 270172 12292
rect 270228 12236 270238 12292
rect 189298 12124 189308 12180
rect 189364 12124 191100 12180
rect 191156 12124 191166 12180
rect 192434 12124 192444 12180
rect 192500 12124 193788 12180
rect 193844 12124 193854 12180
rect 228274 12124 228284 12180
rect 228340 12124 238588 12180
rect 238644 12124 238654 12180
rect 243282 12124 243292 12180
rect 243348 12124 244412 12180
rect 244468 12124 244478 12180
rect 244626 12124 244636 12180
rect 244692 12124 245084 12180
rect 245140 12124 245150 12180
rect 245522 12124 245532 12180
rect 245588 12124 246876 12180
rect 246932 12124 246942 12180
rect 249442 12124 249452 12180
rect 249508 12124 249518 12180
rect 249452 12068 249508 12124
rect 165554 12012 165564 12068
rect 165620 12012 203868 12068
rect 203924 12012 203934 12068
rect 215058 12012 215068 12068
rect 215124 12012 233436 12068
rect 233492 12012 233502 12068
rect 238130 12012 238140 12068
rect 238196 12012 249508 12068
rect 199490 11900 199500 11956
rect 199556 11900 202300 11956
rect 202356 11900 202366 11956
rect 244402 11900 244412 11956
rect 244468 11900 248556 11956
rect 248612 11900 248622 11956
rect 237234 11788 237244 11844
rect 237300 11788 238364 11844
rect 238420 11788 238430 11844
rect 238802 11788 238812 11844
rect 238868 11788 240156 11844
rect 240212 11788 240222 11844
rect 242610 11788 242620 11844
rect 242676 11788 243404 11844
rect 243460 11788 243470 11844
rect 175298 11676 175308 11732
rect 175364 11676 200788 11732
rect 201282 11676 201292 11732
rect 201348 11676 202748 11732
rect 202804 11676 202814 11732
rect 213490 11676 213500 11732
rect 213556 11676 216748 11732
rect 216804 11676 216814 11732
rect 229170 11676 229180 11732
rect 229236 11676 231868 11732
rect 233314 11676 233324 11732
rect 233380 11676 268716 11732
rect 268772 11676 268782 11732
rect 158162 11564 158172 11620
rect 158228 11564 200564 11620
rect 135314 11452 135324 11508
rect 135380 11452 200284 11508
rect 200340 11452 200350 11508
rect 200508 11396 200564 11564
rect 200732 11508 200788 11676
rect 211026 11564 211036 11620
rect 211092 11564 218876 11620
rect 218932 11564 218942 11620
rect 231812 11508 231868 11676
rect 237010 11564 237020 11620
rect 237076 11564 267036 11620
rect 267092 11564 267102 11620
rect 200732 11452 204988 11508
rect 205044 11452 205054 11508
rect 212370 11452 212380 11508
rect 212436 11452 230188 11508
rect 230244 11452 230254 11508
rect 231812 11452 249340 11508
rect 249396 11452 249406 11508
rect 129602 11340 129612 11396
rect 129668 11340 199612 11396
rect 199668 11340 199678 11396
rect 200508 11340 202972 11396
rect 203028 11340 203038 11396
rect 217746 11340 217756 11396
rect 217812 11340 251916 11396
rect 251972 11340 251982 11396
rect 49634 11228 49644 11284
rect 49700 11228 134428 11284
rect 134484 11228 134494 11284
rect 141026 11228 141036 11284
rect 141092 11228 200956 11284
rect 201012 11228 201022 11284
rect 228946 11228 228956 11284
rect 229012 11228 270284 11284
rect 270340 11228 270350 11284
rect 430882 11228 430892 11284
rect 430948 11228 468300 11284
rect 468356 11228 468366 11284
rect 78194 11116 78204 11172
rect 78260 11116 193564 11172
rect 193620 11116 193630 11172
rect 223794 11116 223804 11172
rect 223860 11116 265468 11172
rect 265524 11116 265534 11172
rect 265682 11116 265692 11172
rect 265748 11116 270508 11172
rect 270564 11116 270574 11172
rect 431442 11116 431452 11172
rect 431508 11116 544460 11172
rect 544516 11116 544526 11172
rect 47730 11004 47740 11060
rect 47796 11004 189980 11060
rect 190036 11004 190046 11060
rect 196130 11004 196140 11060
rect 196196 11004 207452 11060
rect 207508 11004 207518 11060
rect 227826 11004 227836 11060
rect 227892 11004 269164 11060
rect 269220 11004 269230 11060
rect 441858 11004 441868 11060
rect 441924 11004 561596 11060
rect 561652 11004 561662 11060
rect 32498 10892 32508 10948
rect 32564 10892 188188 10948
rect 188244 10892 188254 10948
rect 190530 10892 190540 10948
rect 190596 10892 206780 10948
rect 206836 10892 206846 10948
rect 221554 10892 221564 10948
rect 221620 10892 268940 10948
rect 268996 10892 269006 10948
rect 431218 10892 431228 10948
rect 431284 10892 563500 10948
rect 563556 10892 563566 10948
rect 171490 10780 171500 10836
rect 171556 10780 190652 10836
rect 190708 10780 190718 10836
rect 218418 10780 218428 10836
rect 218484 10780 236796 10836
rect 236852 10780 236862 10836
rect 220210 10444 220220 10500
rect 220276 10444 275324 10500
rect 275380 10444 275390 10500
rect 312386 10444 312396 10500
rect 312452 10444 420476 10500
rect 420532 10444 420542 10500
rect 420690 10444 420700 10500
rect 420756 10444 425740 10500
rect 425796 10444 425806 10500
rect 269938 10332 269948 10388
rect 270004 10332 287084 10388
rect 287140 10332 287150 10388
rect 413074 10332 413084 10388
rect 413140 10332 423948 10388
rect 424004 10332 424014 10388
rect 218194 10108 218204 10164
rect 218260 10108 220108 10164
rect 249442 10108 249452 10164
rect 249508 10108 264460 10164
rect 264516 10108 264526 10164
rect 265458 10108 265468 10164
rect 265524 10108 269500 10164
rect 269556 10108 269566 10164
rect 273858 10108 273868 10164
rect 273924 10108 310716 10164
rect 310772 10108 310782 10164
rect 169586 9996 169596 10052
rect 169652 9996 200396 10052
rect 200452 9996 200462 10052
rect 201954 9996 201964 10052
rect 202020 9996 208124 10052
rect 208180 9996 208190 10052
rect 160066 9884 160076 9940
rect 160132 9884 199892 9940
rect 200050 9884 200060 9940
rect 200116 9884 207900 9940
rect 207956 9884 207966 9940
rect 199836 9828 199892 9884
rect 220052 9828 220108 10108
rect 230066 9996 230076 10052
rect 230132 9996 268156 10052
rect 268212 9996 268222 10052
rect 270274 9996 270284 10052
rect 270340 9996 275212 10052
rect 275268 9996 275278 10052
rect 239698 9884 239708 9940
rect 239764 9884 266364 9940
rect 266420 9884 266430 9940
rect 269378 9884 269388 9940
rect 269444 9884 269836 9940
rect 269892 9884 269902 9940
rect 272962 9884 272972 9940
rect 273028 9884 314188 9940
rect 314244 9884 314254 9940
rect 152450 9772 152460 9828
rect 152516 9772 199500 9828
rect 199556 9772 199566 9828
rect 199836 9772 203196 9828
rect 203252 9772 203262 9828
rect 204306 9772 204316 9828
rect 204372 9772 204382 9828
rect 220052 9772 277228 9828
rect 277284 9772 277294 9828
rect 204316 9716 204372 9772
rect 112466 9660 112476 9716
rect 112532 9660 197596 9716
rect 197652 9660 197662 9716
rect 200386 9660 200396 9716
rect 200452 9660 204372 9716
rect 216178 9660 216188 9716
rect 216244 9660 238476 9716
rect 238532 9660 238542 9716
rect 241714 9660 241724 9716
rect 241780 9660 267148 9716
rect 267204 9660 267214 9716
rect 272066 9660 272076 9716
rect 272132 9660 365484 9716
rect 365540 9660 365550 9716
rect 398178 9660 398188 9716
rect 398244 9660 428204 9716
rect 428260 9660 428270 9716
rect 97234 9548 97244 9604
rect 97300 9548 195804 9604
rect 195860 9548 195870 9604
rect 224242 9548 224252 9604
rect 224308 9548 331212 9604
rect 331268 9548 331278 9604
rect 370402 9548 370412 9604
rect 370468 9548 421036 9604
rect 421092 9548 421102 9604
rect 89618 9436 89628 9492
rect 89684 9436 194908 9492
rect 194964 9436 194974 9492
rect 224914 9436 224924 9492
rect 224980 9436 336924 9492
rect 336980 9436 336990 9492
rect 358082 9436 358092 9492
rect 358148 9436 426972 9492
rect 427028 9436 427038 9492
rect 61058 9324 61068 9380
rect 61124 9324 191548 9380
rect 191604 9324 191614 9380
rect 211250 9324 211260 9380
rect 211316 9324 220780 9380
rect 220836 9324 220846 9380
rect 225586 9324 225596 9380
rect 225652 9324 342748 9380
rect 342804 9324 342814 9380
rect 346658 9324 346668 9380
rect 346724 9324 420700 9380
rect 420756 9324 420766 9380
rect 24882 9212 24892 9268
rect 24948 9212 187292 9268
rect 187348 9212 187358 9268
rect 188626 9212 188636 9268
rect 188692 9212 206556 9268
rect 206612 9212 206622 9268
rect 212594 9212 212604 9268
rect 212660 9212 232204 9268
rect 232260 9212 232270 9268
rect 234882 9212 234892 9268
rect 234948 9212 399868 9268
rect 399924 9212 399934 9268
rect 408258 9212 408268 9268
rect 408324 9212 426748 9268
rect 426804 9212 426814 9268
rect 177202 9100 177212 9156
rect 177268 9100 205212 9156
rect 205268 9100 205278 9156
rect 235106 9100 235116 9156
rect 235172 9100 249452 9156
rect 249508 9100 249518 9156
rect 269154 9100 269164 9156
rect 269220 9100 277564 9156
rect 277620 9100 277630 9156
rect 249330 8876 249340 8932
rect 249396 8876 257068 8932
rect 257124 8876 257134 8932
rect 392 8792 4172 8820
rect -960 8764 4172 8792
rect 4228 8764 4238 8820
rect 277442 8764 277452 8820
rect 277508 8764 290668 8820
rect 290724 8764 290734 8820
rect 290892 8764 297164 8820
rect 297220 8764 297230 8820
rect -960 8568 480 8764
rect 290892 8708 290948 8764
rect 277330 8652 277340 8708
rect 277396 8652 288988 8708
rect 289044 8652 289054 8708
rect 290612 8652 290948 8708
rect 296268 8652 304108 8708
rect 304164 8652 304174 8708
rect 290612 8596 290668 8652
rect 269714 8540 269724 8596
rect 269780 8540 279132 8596
rect 279188 8540 279198 8596
rect 289090 8540 289100 8596
rect 289156 8540 290668 8596
rect 296268 8484 296324 8652
rect 85810 8428 85820 8484
rect 85876 8428 92316 8484
rect 92372 8428 92382 8484
rect 203858 8428 203868 8484
rect 203924 8428 208348 8484
rect 208404 8428 208414 8484
rect 278898 8428 278908 8484
rect 278964 8428 296324 8484
rect 297276 8540 357196 8596
rect 357252 8540 357262 8596
rect 297276 8372 297332 8540
rect 304098 8428 304108 8484
rect 304164 8428 514220 8484
rect 514276 8428 514286 8484
rect 173394 8316 173404 8372
rect 173460 8316 204764 8372
rect 204820 8316 204830 8372
rect 222674 8316 222684 8372
rect 222740 8316 266700 8372
rect 266756 8316 266766 8372
rect 269266 8316 269276 8372
rect 269332 8316 277340 8372
rect 277396 8316 277406 8372
rect 288978 8316 288988 8372
rect 289044 8316 297332 8372
rect 131506 8204 131516 8260
rect 131572 8204 179116 8260
rect 179172 8204 179182 8260
rect 184706 8204 184716 8260
rect 184772 8204 206108 8260
rect 206164 8204 206174 8260
rect 213938 8204 213948 8260
rect 214004 8204 236796 8260
rect 236852 8204 236862 8260
rect 241042 8204 241052 8260
rect 241108 8204 264572 8260
rect 264628 8204 264638 8260
rect 265458 8204 265468 8260
rect 265524 8204 270172 8260
rect 270228 8204 270238 8260
rect 274082 8204 274092 8260
rect 274148 8204 283612 8260
rect 283668 8204 283678 8260
rect 357186 8204 357196 8260
rect 357252 8204 361676 8260
rect 361732 8204 361742 8260
rect 413186 8204 413196 8260
rect 413252 8204 423724 8260
rect 423780 8204 423790 8260
rect 146738 8092 146748 8148
rect 146804 8092 201628 8148
rect 201684 8092 201694 8148
rect 213266 8092 213276 8148
rect 213332 8092 237916 8148
rect 237972 8092 237982 8148
rect 245746 8092 245756 8148
rect 245812 8092 266476 8148
rect 266532 8092 266542 8148
rect 269266 8092 269276 8148
rect 269332 8092 293132 8148
rect 293188 8092 293198 8148
rect 403778 8092 403788 8148
rect 403844 8092 423612 8148
rect 423668 8092 423678 8148
rect 442978 8092 442988 8148
rect 443044 8092 449260 8148
rect 449316 8092 449326 8148
rect 108658 7980 108668 8036
rect 108724 7980 197148 8036
rect 197204 7980 197214 8036
rect 226930 7980 226940 8036
rect 226996 7980 265804 8036
rect 265860 7980 265870 8036
rect 269490 7980 269500 8036
rect 269556 7980 319788 8036
rect 319844 7980 319854 8036
rect 398066 7980 398076 8036
rect 398132 7980 422044 8036
rect 422100 7980 422110 8036
rect 429426 7980 429436 8036
rect 429492 7980 456988 8036
rect 457044 7980 457054 8036
rect 91522 7868 91532 7924
rect 91588 7868 195132 7924
rect 195188 7868 195198 7924
rect 229618 7868 229628 7924
rect 229684 7868 376908 7924
rect 376964 7868 376974 7924
rect 380930 7868 380940 7924
rect 380996 7868 421484 7924
rect 421540 7868 421550 7924
rect 439282 7868 439292 7924
rect 439348 7868 500668 7924
rect 500724 7868 500734 7924
rect 83906 7756 83916 7812
rect 83972 7756 192332 7812
rect 192388 7756 192398 7812
rect 214162 7756 214172 7812
rect 214228 7756 228620 7812
rect 228676 7756 228686 7812
rect 230402 7756 230412 7812
rect 230468 7756 382620 7812
rect 382676 7756 382686 7812
rect 386642 7756 386652 7812
rect 386708 7756 422268 7812
rect 422324 7756 422334 7812
rect 444098 7756 444108 7812
rect 444164 7756 552076 7812
rect 552132 7756 552142 7812
rect 62962 7644 62972 7700
rect 63028 7644 81452 7700
rect 81508 7644 81518 7700
rect 82002 7644 82012 7700
rect 82068 7644 194012 7700
rect 194068 7644 194078 7700
rect 215506 7644 215516 7700
rect 215572 7644 233436 7700
rect 233492 7644 233502 7700
rect 234322 7644 234332 7700
rect 234388 7644 428428 7700
rect 428484 7644 428494 7700
rect 436258 7644 436268 7700
rect 436324 7644 580636 7700
rect 580692 7644 580702 7700
rect 21074 7532 21084 7588
rect 21140 7532 44492 7588
rect 44548 7532 44558 7588
rect 72482 7532 72492 7588
rect 72548 7532 192892 7588
rect 192948 7532 192958 7588
rect 213714 7532 213724 7588
rect 213780 7532 235116 7588
rect 235172 7532 235182 7588
rect 235666 7532 235676 7588
rect 235732 7532 445452 7588
rect 445508 7532 445518 7588
rect 179106 7420 179116 7476
rect 179172 7420 204092 7476
rect 204148 7420 204158 7476
rect 595560 7140 597000 7336
rect 290612 7084 302652 7140
rect 302708 7084 302718 7140
rect 442754 7084 442764 7140
rect 442820 7112 597000 7140
rect 442820 7084 595672 7112
rect 270498 6972 270508 7028
rect 270564 6972 275436 7028
rect 275492 6972 275502 7028
rect 280802 6972 280812 7028
rect 280868 6972 285852 7028
rect 285908 6972 285918 7028
rect 290612 6916 290668 7084
rect 295810 6972 295820 7028
rect 295876 6972 354060 7028
rect 354116 6972 354126 7028
rect 363794 6972 363804 7028
rect 363860 6972 370412 7028
rect 370468 6972 370478 7028
rect 273298 6860 273308 6916
rect 273364 6860 281708 6916
rect 281764 6860 281774 6916
rect 285618 6860 285628 6916
rect 285684 6860 290668 6916
rect 303986 6860 303996 6916
rect 304052 6860 373100 6916
rect 373156 6860 373166 6916
rect 390450 6860 390460 6916
rect 390516 6860 398188 6916
rect 398244 6860 398254 6916
rect 51538 6748 51548 6804
rect 51604 6748 54572 6804
rect 54628 6748 54638 6804
rect 210578 6748 210588 6804
rect 210644 6748 215068 6804
rect 215124 6748 215134 6804
rect 267092 6748 411180 6804
rect 411236 6748 411246 6804
rect 425058 6748 425068 6804
rect 425124 6748 428764 6804
rect 428820 6748 428830 6804
rect 514210 6748 514220 6804
rect 514276 6748 521612 6804
rect 521668 6748 521678 6804
rect 571218 6748 571228 6804
rect 571284 6748 574924 6804
rect 574980 6748 574990 6804
rect 163874 6636 163884 6692
rect 163940 6636 203644 6692
rect 203700 6636 203710 6692
rect 228722 6636 228732 6692
rect 228788 6636 266252 6692
rect 266308 6636 266318 6692
rect 267092 6580 267148 6748
rect 272962 6636 272972 6692
rect 273028 6636 289100 6692
rect 289156 6636 289166 6692
rect 290658 6636 290668 6692
rect 290724 6636 295820 6692
rect 295876 6636 295886 6692
rect 127586 6524 127596 6580
rect 127652 6524 199388 6580
rect 199444 6524 199454 6580
rect 237794 6524 237804 6580
rect 237860 6524 267148 6580
rect 268930 6524 268940 6580
rect 268996 6524 308364 6580
rect 308420 6524 308430 6580
rect 121986 6412 121996 6468
rect 122052 6412 198716 6468
rect 198772 6412 198782 6468
rect 211474 6412 211484 6468
rect 211540 6412 222684 6468
rect 222740 6412 222750 6468
rect 237458 6412 237468 6468
rect 237524 6412 266812 6468
rect 266868 6412 266878 6468
rect 269714 6412 269724 6468
rect 269780 6412 285628 6468
rect 285684 6412 285694 6468
rect 297154 6412 297164 6468
rect 297220 6412 348348 6468
rect 348404 6412 348414 6468
rect 394818 6412 394828 6468
rect 394884 6412 408268 6468
rect 408324 6412 408334 6468
rect 116274 6300 116284 6356
rect 116340 6300 198044 6356
rect 198100 6300 198110 6356
rect 214386 6300 214396 6356
rect 214452 6300 230188 6356
rect 230244 6300 230254 6356
rect 244514 6300 244524 6356
rect 244580 6300 265244 6356
rect 265300 6300 265310 6356
rect 271618 6300 271628 6356
rect 271684 6300 280812 6356
rect 280868 6300 280878 6356
rect 287074 6300 287084 6356
rect 287140 6300 350252 6356
rect 350308 6300 350318 6356
rect 401874 6300 401884 6356
rect 401940 6300 425628 6356
rect 425684 6300 425694 6356
rect 34402 6188 34412 6244
rect 34468 6188 116732 6244
rect 116788 6188 116798 6244
rect 120082 6188 120092 6244
rect 120148 6188 198492 6244
rect 198548 6188 198558 6244
rect 217970 6188 217980 6244
rect 218036 6188 277900 6244
rect 277956 6188 277966 6244
rect 288978 6188 288988 6244
rect 289044 6188 295372 6244
rect 295428 6188 295438 6244
rect 340946 6188 340956 6244
rect 341012 6188 426860 6244
rect 426916 6188 426926 6244
rect 70466 6076 70476 6132
rect 70532 6076 191436 6132
rect 191492 6076 191502 6132
rect 211698 6076 211708 6132
rect 211764 6076 224588 6132
rect 224644 6076 224654 6132
rect 227602 6076 227612 6132
rect 227668 6076 359772 6132
rect 359828 6076 359838 6132
rect 362786 6076 362796 6132
rect 362852 6076 425068 6132
rect 425124 6076 425134 6132
rect 66770 5964 66780 6020
rect 66836 5964 192220 6020
rect 192276 5964 192286 6020
rect 219538 5964 219548 6020
rect 219604 5964 291228 6020
rect 291284 5964 291294 6020
rect 310706 5964 310716 6020
rect 310772 5964 451164 6020
rect 451220 5964 451230 6020
rect 30594 5852 30604 5908
rect 30660 5852 187964 5908
rect 188020 5852 188030 5908
rect 214834 5852 214844 5908
rect 214900 5852 226828 5908
rect 226884 5852 226894 5908
rect 230962 5852 230972 5908
rect 231028 5852 388332 5908
rect 388388 5852 388398 5908
rect 392354 5852 392364 5908
rect 392420 5852 423500 5908
rect 423556 5852 423566 5908
rect 429538 5852 429548 5908
rect 429604 5852 462588 5908
rect 462644 5852 462654 5908
rect 181010 5740 181020 5796
rect 181076 5740 205660 5796
rect 205716 5740 205726 5796
rect 269938 5740 269948 5796
rect 270004 5740 300748 5796
rect 300804 5740 300814 5796
rect 275202 5292 275212 5348
rect 275268 5292 275660 5348
rect 275716 5292 275726 5348
rect 275426 5180 275436 5236
rect 275492 5180 285740 5236
rect 285796 5180 285806 5236
rect 295474 5180 295484 5236
rect 295540 5180 324268 5236
rect 324324 5180 324334 5236
rect 265458 5068 265468 5124
rect 265524 5068 268044 5124
rect 268100 5068 268110 5124
rect 275538 5068 275548 5124
rect 275604 5068 295764 5124
rect 296482 5068 296492 5124
rect 296548 5068 303996 5124
rect 304052 5068 304062 5124
rect 307346 5068 307356 5124
rect 307412 5068 337708 5124
rect 295708 5012 295764 5068
rect 186722 4956 186732 5012
rect 186788 4956 206332 5012
rect 206388 4956 206398 5012
rect 239474 4956 239484 5012
rect 239540 4956 268492 5012
rect 268548 4956 268558 5012
rect 295708 4956 298900 5012
rect 298844 4900 298900 4956
rect 182914 4844 182924 4900
rect 182980 4844 205884 4900
rect 205940 4844 205950 4900
rect 235106 4844 235116 4900
rect 235172 4844 241724 4900
rect 241780 4844 241790 4900
rect 241938 4844 241948 4900
rect 242004 4844 268044 4900
rect 268100 4844 268110 4900
rect 277218 4844 277228 4900
rect 277284 4844 279804 4900
rect 279860 4844 279870 4900
rect 287298 4844 287308 4900
rect 287364 4844 296492 4900
rect 296548 4844 296558 4900
rect 298834 4844 298844 4900
rect 298900 4844 298910 4900
rect 337652 4788 337708 5068
rect 546802 4956 546812 5012
rect 546868 4956 550172 5012
rect 550228 4956 550238 5012
rect 419010 4844 419020 4900
rect 419076 4844 424172 4900
rect 424228 4844 424238 4900
rect 442754 4844 442764 4900
rect 442820 4844 454972 4900
rect 455028 4844 455038 4900
rect 156146 4732 156156 4788
rect 156212 4732 201292 4788
rect 201348 4732 201358 4788
rect 238466 4732 238476 4788
rect 238532 4732 243628 4788
rect 243954 4732 243964 4788
rect 244020 4732 265468 4788
rect 265524 4732 265534 4788
rect 271506 4732 271516 4788
rect 271572 4732 320908 4788
rect 320964 4732 320974 4788
rect 337652 4732 367388 4788
rect 367444 4732 367454 4788
rect 417106 4732 417116 4788
rect 417172 4732 425068 4788
rect 425124 4732 425134 4788
rect 442978 4732 442988 4788
rect 443044 4732 466396 4788
rect 466452 4732 466462 4788
rect 243572 4676 243628 4732
rect 93426 4620 93436 4676
rect 93492 4620 195356 4676
rect 195412 4620 195422 4676
rect 216738 4620 216748 4676
rect 216804 4620 239820 4676
rect 239876 4620 239886 4676
rect 243572 4620 256228 4676
rect 257058 4620 257068 4676
rect 257124 4620 265692 4676
rect 265748 4620 265758 4676
rect 273186 4620 273196 4676
rect 273252 4620 344540 4676
rect 344596 4620 344606 4676
rect 444210 4620 444220 4676
rect 444276 4620 483532 4676
rect 483588 4620 483598 4676
rect 256172 4564 256228 4620
rect 80098 4508 80108 4564
rect 80164 4508 192444 4564
rect 192500 4508 192510 4564
rect 226818 4508 226828 4564
rect 226884 4508 251244 4564
rect 251300 4508 251310 4564
rect 256172 4508 262108 4564
rect 267810 4508 267820 4564
rect 267876 4508 333116 4564
rect 333172 4508 333182 4564
rect 335234 4508 335244 4564
rect 335300 4508 413196 4564
rect 413252 4508 413262 4564
rect 415202 4508 415212 4564
rect 415268 4508 428428 4564
rect 428484 4508 428494 4564
rect 437602 4508 437612 4564
rect 437668 4508 477820 4564
rect 477876 4508 477886 4564
rect 43922 4396 43932 4452
rect 43988 4396 189532 4452
rect 189588 4396 189598 4452
rect 209234 4396 209244 4452
rect 209300 4396 211260 4452
rect 211316 4396 211326 4452
rect 212818 4396 212828 4452
rect 212884 4396 220108 4452
rect 233426 4396 233436 4452
rect 233492 4396 257068 4452
rect 257124 4396 257134 4452
rect 220052 4340 220108 4396
rect 262052 4340 262108 4508
rect 270162 4396 270172 4452
rect 270228 4396 274372 4452
rect 275314 4396 275324 4452
rect 275380 4396 296940 4452
rect 296996 4396 297006 4452
rect 318098 4396 318108 4452
rect 318164 4396 394828 4452
rect 394884 4396 394894 4452
rect 407586 4396 407596 4452
rect 407652 4396 420700 4452
rect 420756 4396 420766 4452
rect 443426 4396 443436 4452
rect 443492 4396 496860 4452
rect 496916 4396 496926 4452
rect 502292 4396 537628 4452
rect 274316 4340 274372 4396
rect 502292 4340 502348 4396
rect 537572 4340 537628 4396
rect 22978 4284 22988 4340
rect 23044 4284 23436 4340
rect 23492 4284 23502 4340
rect 28690 4284 28700 4340
rect 28756 4284 187740 4340
rect 187796 4284 187806 4340
rect 210802 4284 210812 4340
rect 210868 4284 216972 4340
rect 217028 4284 217038 4340
rect 220052 4284 234108 4340
rect 234164 4284 234174 4340
rect 242834 4284 242844 4340
rect 242900 4284 249508 4340
rect 262052 4284 262668 4340
rect 262724 4284 262734 4340
rect 270386 4284 270396 4340
rect 270452 4284 274092 4340
rect 274148 4284 274158 4340
rect 274316 4284 327404 4340
rect 327460 4284 327470 4340
rect 329522 4284 329532 4340
rect 329588 4284 420588 4340
rect 420644 4284 420654 4340
rect 421708 4284 428820 4340
rect 429314 4284 429324 4340
rect 429380 4284 502348 4340
rect 523478 4284 523516 4340
rect 523572 4284 523582 4340
rect 531094 4284 531132 4340
rect 531188 4284 531198 4340
rect 537572 4284 548268 4340
rect 548324 4284 548334 4340
rect 249452 4228 249508 4284
rect 421708 4228 421764 4284
rect 428764 4228 428820 4284
rect 17238 4172 17276 4228
rect 17332 4172 17342 4228
rect 19170 4172 19180 4228
rect 19236 4172 186620 4228
rect 186676 4172 186686 4228
rect 198146 4172 198156 4228
rect 198212 4172 207676 4228
rect 207732 4172 207742 4228
rect 210354 4172 210364 4228
rect 210420 4172 213164 4228
rect 213220 4172 213230 4228
rect 220052 4172 236012 4228
rect 236068 4172 236078 4228
rect 236786 4172 236796 4228
rect 236852 4172 243628 4228
rect 243684 4172 243694 4228
rect 249452 4172 272020 4228
rect 272150 4172 272188 4228
rect 272244 4172 272254 4228
rect 278852 4172 352716 4228
rect 352772 4172 352782 4228
rect 409490 4172 409500 4228
rect 409556 4172 421764 4228
rect 421922 4172 421932 4228
rect 421988 4172 422604 4228
rect 422660 4172 422670 4228
rect 423826 4172 423836 4228
rect 423892 4172 424508 4228
rect 424564 4172 424574 4228
rect 426626 4172 426636 4228
rect 426692 4172 428540 4228
rect 428596 4172 428606 4228
rect 428764 4172 430220 4228
rect 430276 4172 430286 4228
rect 431778 4172 431788 4228
rect 431844 4172 432124 4228
rect 432180 4172 432190 4228
rect 436818 4172 436828 4228
rect 436884 4172 437836 4228
rect 437892 4172 437902 4228
rect 443202 4172 443212 4228
rect 443268 4172 573020 4228
rect 573076 4172 573086 4228
rect 581298 4172 581308 4228
rect 581364 4172 582540 4228
rect 582596 4172 582606 4228
rect 220052 4116 220108 4172
rect 271964 4116 272020 4172
rect 278852 4116 278908 4172
rect 36306 4060 36316 4116
rect 36372 4060 37772 4116
rect 37828 4060 37838 4116
rect 42018 4060 42028 4116
rect 42084 4060 42812 4116
rect 42868 4060 42878 4116
rect 68674 4060 68684 4116
rect 68740 4060 69692 4116
rect 69748 4060 69758 4116
rect 213042 4060 213052 4116
rect 213108 4060 220108 4116
rect 230178 4060 230188 4116
rect 230244 4060 247436 4116
rect 247492 4060 247502 4116
rect 251906 4060 251916 4116
rect 251972 4060 267148 4116
rect 271964 4060 278908 4116
rect 352370 4060 352380 4116
rect 352436 4060 362796 4116
rect 362852 4060 362862 4116
rect 420914 4060 420924 4116
rect 420980 4060 430108 4116
rect 430164 4060 430174 4116
rect 479686 4060 479724 4116
rect 479780 4060 479790 4116
rect 267092 4004 267148 4060
rect 228610 3948 228620 4004
rect 228676 3948 245532 4004
rect 245588 3948 245598 4004
rect 267092 3948 275996 4004
rect 276052 3948 276062 4004
rect 540614 3948 540652 4004
rect 540708 3948 540718 4004
rect 55318 3836 55356 3892
rect 55412 3836 55422 3892
rect 546326 3836 546364 3892
rect 546420 3836 546430 3892
rect 40114 3724 40124 3780
rect 40180 3724 41804 3780
rect 41860 3724 41870 3780
rect 267092 3724 282156 3780
rect 282212 3724 282222 3780
rect 285618 3724 285628 3780
rect 285684 3724 290668 3780
rect 297378 3724 297388 3780
rect 297444 3724 310268 3780
rect 310324 3724 310334 3780
rect 323810 3724 323820 3780
rect 323876 3724 416668 3780
rect 416724 3724 416734 3780
rect 557750 3724 557788 3780
rect 557844 3724 557854 3780
rect 267092 3668 267148 3724
rect 248546 3612 248556 3668
rect 248612 3612 267148 3668
rect 280466 3612 280476 3668
rect 280532 3612 287420 3668
rect 287476 3612 287486 3668
rect 290612 3556 290668 3724
rect 375218 3612 375228 3668
rect 375284 3612 398076 3668
rect 398132 3612 398142 3668
rect 275762 3500 275772 3556
rect 275828 3500 287364 3556
rect 290612 3500 297612 3556
rect 297668 3500 297678 3556
rect 309138 3500 309148 3556
rect 309204 3500 321692 3556
rect 321748 3500 321758 3556
rect 361172 3500 378812 3556
rect 378868 3500 378878 3556
rect 11526 3388 11564 3444
rect 11620 3388 11630 3444
rect 13318 3388 13356 3444
rect 13412 3388 13422 3444
rect 26758 3388 26796 3444
rect 26852 3388 26862 3444
rect 265570 3388 265580 3444
rect 265636 3388 275604 3444
rect 275548 3332 275604 3388
rect 287308 3332 287364 3500
rect 296492 3388 315980 3444
rect 316036 3388 316046 3444
rect 296492 3332 296548 3388
rect 361172 3332 361228 3500
rect 369506 3388 369516 3444
rect 369572 3388 372988 3444
rect 394006 3388 394044 3444
rect 394100 3388 394110 3444
rect 397730 3388 397740 3444
rect 397796 3388 406588 3444
rect 406644 3388 406654 3444
rect 506342 3388 506380 3444
rect 506436 3388 506446 3444
rect 512054 3388 512092 3444
rect 512148 3388 512158 3444
rect 517766 3388 517804 3444
rect 517860 3388 517870 3444
rect 534902 3388 534940 3444
rect 534996 3388 535006 3444
rect 552626 3388 552636 3444
rect 552692 3388 555884 3444
rect 555940 3388 555950 3444
rect 559654 3388 559692 3444
rect 559748 3388 559758 3444
rect 571190 3388 571228 3444
rect 571284 3388 571294 3444
rect 150546 3276 150556 3332
rect 150612 3276 202076 3332
rect 202132 3276 202142 3332
rect 221778 3276 221788 3332
rect 221844 3276 230188 3332
rect 230244 3276 230254 3332
rect 234994 3276 235004 3332
rect 235060 3276 264684 3332
rect 264740 3276 264750 3332
rect 275548 3276 278908 3332
rect 278964 3276 278974 3332
rect 287308 3276 296548 3332
rect 304098 3276 304108 3332
rect 304164 3276 361228 3332
rect 372932 3332 372988 3388
rect 372932 3276 421820 3332
rect 421876 3276 421886 3332
rect 139122 3164 139132 3220
rect 139188 3164 200732 3220
rect 200788 3164 200798 3220
rect 225138 3164 225148 3220
rect 225204 3164 248556 3220
rect 248612 3164 248622 3220
rect 270498 3164 270508 3220
rect 270564 3164 275772 3220
rect 275828 3164 275838 3220
rect 294018 3164 294028 3220
rect 294084 3164 307356 3220
rect 307412 3164 307422 3220
rect 324258 3164 324268 3220
rect 324324 3164 371308 3220
rect 371364 3164 371374 3220
rect 123890 3052 123900 3108
rect 123956 3052 198940 3108
rect 198996 3052 199006 3108
rect 232306 3052 232316 3108
rect 232372 3052 265244 3108
rect 265300 3052 265310 3108
rect 265794 3052 265804 3108
rect 265860 3052 277452 3108
rect 277508 3052 277518 3108
rect 285730 3052 285740 3108
rect 285796 3052 355964 3108
rect 356020 3052 356030 3108
rect 416658 3052 416668 3108
rect 416724 3052 422156 3108
rect 422212 3052 422222 3108
rect 110562 2940 110572 2996
rect 110628 2940 197372 2996
rect 197428 2940 197438 2996
rect 264450 2940 264460 2996
rect 264516 2940 405468 2996
rect 405524 2940 405534 2996
rect 99026 2828 99036 2884
rect 99092 2828 196028 2884
rect 196084 2828 196094 2884
rect 234210 2828 234220 2884
rect 234276 2828 266588 2884
rect 266644 2828 266654 2884
rect 285572 2828 297388 2884
rect 297444 2828 297454 2884
rect 320898 2828 320908 2884
rect 320964 2828 489244 2884
rect 489300 2828 489310 2884
rect 285572 2772 285628 2828
rect 95330 2716 95340 2772
rect 95396 2716 193452 2772
rect 193508 2716 193518 2772
rect 235890 2716 235900 2772
rect 235956 2716 268156 2772
rect 268212 2716 268222 2772
rect 280354 2716 280364 2772
rect 280420 2716 285628 2772
rect 285740 2716 289324 2772
rect 289380 2716 289390 2772
rect 297602 2716 297612 2772
rect 297668 2716 325500 2772
rect 325556 2716 325566 2772
rect 352706 2716 352716 2772
rect 352772 2716 536844 2772
rect 536900 2716 536910 2772
rect 285740 2660 285796 2716
rect 57250 2604 57260 2660
rect 57316 2604 189308 2660
rect 189364 2604 189374 2660
rect 219314 2604 219324 2660
rect 219380 2604 285796 2660
rect 286066 2604 286076 2660
rect 286132 2604 304556 2660
rect 304612 2604 304622 2660
rect 308242 2604 308252 2660
rect 308308 2604 494956 2660
rect 495012 2604 495022 2660
rect 15362 2492 15372 2548
rect 15428 2492 185724 2548
rect 185780 2492 185790 2548
rect 265458 2492 265468 2548
rect 265524 2492 275548 2548
rect 275604 2492 275614 2548
rect 277218 2492 277228 2548
rect 277284 2492 502572 2548
rect 502628 2492 502638 2548
rect 161970 2380 161980 2436
rect 162036 2380 203420 2436
rect 203476 2380 203486 2436
rect 229842 2380 229852 2436
rect 229908 2380 265580 2436
rect 265636 2380 265646 2436
rect 277554 2380 277564 2436
rect 277620 2380 295036 2436
rect 295092 2380 295102 2436
rect 295362 2380 295372 2436
rect 295428 2380 308252 2436
rect 308308 2380 308318 2436
rect 223570 2268 223580 2324
rect 223636 2268 285628 2324
rect 285684 2268 285694 2324
rect 265682 2156 265692 2212
rect 265748 2156 287308 2212
rect 287364 2156 287374 2212
rect 233202 2044 233212 2100
rect 233268 2044 269836 2100
rect 269892 2044 269902 2100
rect 275650 2044 275660 2100
rect 275716 2044 295484 2100
rect 295540 2044 295550 2100
rect 305666 1932 305676 1988
rect 305732 1932 309148 1988
rect 309204 1932 309214 1988
rect 248668 1708 252812 1764
rect 252868 1708 252878 1764
rect 307356 1708 338828 1764
rect 338884 1708 338894 1764
rect 475878 1708 475916 1764
rect 475972 1708 475982 1764
rect 515862 1708 515900 1764
rect 515956 1708 515966 1764
rect 542630 1708 542668 1764
rect 542724 1708 542734 1764
rect 248668 1652 248724 1708
rect 307356 1652 307412 1708
rect 232754 1596 232764 1652
rect 232820 1596 248724 1652
rect 269826 1596 269836 1652
rect 269892 1596 280476 1652
rect 280532 1596 280542 1652
rect 282146 1596 282156 1652
rect 282212 1596 307412 1652
rect 398066 1596 398076 1652
rect 398132 1596 421708 1652
rect 421764 1596 421774 1652
rect 233650 1484 233660 1540
rect 233716 1484 267932 1540
rect 267988 1484 267998 1540
rect 273074 1484 273084 1540
rect 273140 1484 305676 1540
rect 305732 1484 305742 1540
rect 406578 1484 406588 1540
rect 406644 1484 423388 1540
rect 423444 1484 423454 1540
rect 234546 1372 234556 1428
rect 234612 1372 268492 1428
rect 268548 1372 268558 1428
rect 279122 1372 279132 1428
rect 279188 1372 294028 1428
rect 294084 1372 294094 1428
rect 230514 1260 230524 1316
rect 230580 1260 248668 1316
rect 248724 1260 248734 1316
rect 185602 1148 185612 1204
rect 185668 1148 196364 1204
rect 196420 1148 196430 1204
rect 235442 1148 235452 1204
rect 235508 1148 249564 1204
rect 249620 1148 249630 1204
rect 173012 1036 176428 1092
rect 186050 1036 186060 1092
rect 186116 1036 196476 1092
rect 196532 1036 196542 1092
rect 230178 1036 230188 1092
rect 230244 1036 280364 1092
rect 280420 1036 280430 1092
rect 173012 868 173068 1036
rect 176372 980 176428 1036
rect 176372 924 188188 980
rect 247762 924 247772 980
rect 247828 924 265468 980
rect 265524 924 265534 980
rect 125794 812 125804 868
rect 125860 812 173068 868
rect 188132 868 188188 924
rect 188132 812 197484 868
rect 197540 812 197550 868
rect 102946 700 102956 756
rect 103012 700 186060 756
rect 186116 700 186126 756
rect 193330 700 193340 756
rect 193396 700 193406 756
rect 193340 644 193396 700
rect 101042 588 101052 644
rect 101108 588 185612 644
rect 185668 588 185678 644
rect 191492 588 193396 644
rect 232082 588 232092 644
rect 232148 588 236628 644
rect 237682 588 237692 644
rect 237748 588 470204 644
rect 470260 588 470270 644
rect 473974 588 474012 644
rect 474068 588 474078 644
rect 485510 588 485548 644
rect 485604 588 485614 644
rect 527286 588 527324 644
rect 527380 588 527390 644
rect 532998 588 533036 644
rect 533092 588 533102 644
rect 553942 588 553980 644
rect 554036 588 554046 644
rect 191492 532 191548 588
rect 236572 532 236628 588
rect 76402 476 76412 532
rect 76468 476 191548 532
rect 191986 476 191996 532
rect 192052 476 192062 532
rect 236338 476 236348 532
rect 236404 476 236414 532
rect 236572 476 243628 532
rect 270610 476 270620 532
rect 270676 476 285404 532
rect 285460 476 285470 532
rect 306786 476 306796 532
rect 306852 476 397740 532
rect 397796 476 397806 532
rect 191996 420 192052 476
rect 65426 364 65436 420
rect 65492 364 192052 420
rect 59266 252 59276 308
rect 59332 252 191324 308
rect 191380 252 191390 308
rect 236348 196 236404 476
rect 243572 308 243628 476
rect 248658 364 248668 420
rect 248724 364 384412 420
rect 384468 364 384478 420
rect 243572 252 395836 308
rect 395892 252 395902 308
rect 45938 140 45948 196
rect 46004 140 189644 196
rect 189700 140 189710 196
rect 236348 140 452956 196
rect 453012 140 453022 196
rect 38322 28 38332 84
rect 38388 28 188860 84
rect 188916 28 188926 84
<< via3 >>
rect 549388 591052 549444 591108
rect 548044 590940 548100 590996
rect 29484 590828 29540 590884
rect 548156 590828 548212 590884
rect 28364 590716 28420 590772
rect 547708 590716 547764 590772
rect 26796 590604 26852 590660
rect 549612 590604 549668 590660
rect 28476 590492 28532 590548
rect 548268 590492 548324 590548
rect 590492 588588 590548 588644
rect 3388 587132 3444 587188
rect 29372 577276 29428 577332
rect 28028 576044 28084 576100
rect 29260 575932 29316 575988
rect 29148 575820 29204 575876
rect 28140 575708 28196 575764
rect 29036 575596 29092 575652
rect 547820 575596 547876 575652
rect 28252 575484 28308 575540
rect 549500 575484 549556 575540
rect 26460 575372 26516 575428
rect 547932 575372 547988 575428
rect 26572 575036 26628 575092
rect 26684 574476 26740 574532
rect 12572 573020 12628 573076
rect 590604 562156 590660 562212
rect 3500 558908 3556 558964
rect 590716 548940 590772 548996
rect 4172 544796 4228 544852
rect 14252 530684 14308 530740
rect 4284 516572 4340 516628
rect 590828 509292 590884 509348
rect 4396 502460 4452 502516
rect 4508 488348 4564 488404
rect 4732 474236 4788 474292
rect 4620 460124 4676 460180
rect 17612 446012 17668 446068
rect 4844 431900 4900 431956
rect 3948 417788 4004 417844
rect 3388 416668 3444 416724
rect 4956 403676 5012 403732
rect 3500 403228 3556 403284
rect 28028 394492 28084 394548
rect 4396 394268 4452 394324
rect 152012 394268 152068 394324
rect 442652 394268 442708 394324
rect 4844 394156 4900 394212
rect 162092 394156 162148 394212
rect 437612 394156 437668 394212
rect 4172 394044 4228 394100
rect 162316 394044 162372 394100
rect 427532 394044 427588 394100
rect 590604 394044 590660 394100
rect 3948 393932 4004 393988
rect 166012 393932 166068 393988
rect 28140 393148 28196 393204
rect 26460 393036 26516 393092
rect 443436 392924 443492 392980
rect 548268 392924 548324 392980
rect 442876 392812 442932 392868
rect 548156 392812 548212 392868
rect 443212 392700 443268 392756
rect 549612 392700 549668 392756
rect 4620 390684 4676 390740
rect 162204 390684 162260 390740
rect 436268 390684 436324 390740
rect 4284 390572 4340 390628
rect 165900 390572 165956 390628
rect 434252 390572 434308 390628
rect 590492 390572 590548 390628
rect 437724 390348 437780 390404
rect 26572 389788 26628 389844
rect 26684 389676 26740 389732
rect 29148 389676 29204 389732
rect 169708 389564 169764 389620
rect 29036 389452 29092 389508
rect 549388 389340 549444 389396
rect 440076 389004 440132 389060
rect 590716 389004 590772 389060
rect 432684 388892 432740 388948
rect 547708 386092 547764 386148
rect 432572 385532 432628 385588
rect 4732 383964 4788 384020
rect 152124 383964 152180 384020
rect 4508 383852 4564 383908
rect 165788 383852 165844 383908
rect 29260 382956 29316 383012
rect 434476 380604 434532 380660
rect 425852 378812 425908 378868
rect 28252 377356 28308 377412
rect 12572 377244 12628 377300
rect 163996 377244 164052 377300
rect 424172 377132 424228 377188
rect 29484 375564 29540 375620
rect 152236 375452 152292 375508
rect 165452 375452 165508 375508
rect 441196 375340 441252 375396
rect 153804 374780 153860 374836
rect 420924 374780 420980 374836
rect 29372 374556 29428 374612
rect 547932 374556 547988 374612
rect 160748 374108 160804 374164
rect 422604 374108 422660 374164
rect 28364 373996 28420 374052
rect 26796 373884 26852 373940
rect 549500 373884 549556 373940
rect 14252 373772 14308 373828
rect 163884 373772 163940 373828
rect 160524 373436 160580 373492
rect 417564 373436 417620 373492
rect 437948 373100 438004 373156
rect 153692 372764 153748 372820
rect 432908 372764 432964 372820
rect 28476 372316 28532 372372
rect 4956 372204 5012 372260
rect 150780 372204 150836 372260
rect 547820 372204 547876 372260
rect 17612 372092 17668 372148
rect 163772 372092 163828 372148
rect 168812 372092 168868 372148
rect 417676 372092 417732 372148
rect 4284 371420 4340 371476
rect 150332 371420 150388 371476
rect 157164 371420 157220 371476
rect 417900 371420 417956 371476
rect 4172 371308 4228 371364
rect 150556 371308 150612 371364
rect 160412 370748 160468 370804
rect 421036 370748 421092 370804
rect 169820 370076 169876 370132
rect 425964 370076 426020 370132
rect 155036 369404 155092 369460
rect 427980 369404 428036 369460
rect 155596 368732 155652 368788
rect 418348 368732 418404 368788
rect 155372 368060 155428 368116
rect 440972 368060 441028 368116
rect 156828 367388 156884 367444
rect 429436 367388 429492 367444
rect 157052 367052 157108 367108
rect 169820 367052 169876 367108
rect 155148 366716 155204 366772
rect 432796 366716 432852 366772
rect 157836 366044 157892 366100
rect 419020 366044 419076 366100
rect 418348 365484 418404 365540
rect 441084 365484 441140 365540
rect 170828 365372 170884 365428
rect 419916 365372 419972 365428
rect 153916 364700 153972 364756
rect 416108 364700 416164 364756
rect 169820 364028 169876 364084
rect 420812 364028 420868 364084
rect 170492 363356 170548 363412
rect 437388 363356 437444 363412
rect 154364 362796 154420 362852
rect 160748 362796 160804 362852
rect 172620 362684 172676 362740
rect 438396 362684 438452 362740
rect 160300 362124 160356 362180
rect 169820 362124 169876 362180
rect 167468 362012 167524 362068
rect 422492 362012 422548 362068
rect 165452 361676 165508 361732
rect 441196 361676 441252 361732
rect 4172 361564 4228 361620
rect 161196 361340 161252 361396
rect 420700 361340 420756 361396
rect 170268 360668 170324 360724
rect 419804 360668 419860 360724
rect 156940 360332 156996 360388
rect 170828 360332 170884 360388
rect 421036 360332 421092 360388
rect 441196 360332 441252 360388
rect 169260 359996 169316 360052
rect 434924 359996 434980 360052
rect 166124 359324 166180 359380
rect 417452 359324 417508 359380
rect 157724 358652 157780 358708
rect 442540 358652 442596 358708
rect 153804 358092 153860 358148
rect 420924 358092 420980 358148
rect 154476 357868 154532 357924
rect 160524 357868 160580 357924
rect 419692 357980 419748 358036
rect 173180 357532 173236 357588
rect 171052 357308 171108 357364
rect 431228 357308 431284 357364
rect 422604 356972 422660 357028
rect 440188 356972 440244 357028
rect 169372 356636 169428 356692
rect 417788 356636 417844 356692
rect 158508 355964 158564 356020
rect 421596 355964 421652 356020
rect 169820 355292 169876 355348
rect 436604 355292 436660 355348
rect 167580 355068 167636 355124
rect 170268 355068 170324 355124
rect 172508 354620 172564 354676
rect 433244 354620 433300 354676
rect 154364 354508 154420 354564
rect 440188 354508 440244 354564
rect 156156 353948 156212 354004
rect 415772 353948 415828 354004
rect 150892 353612 150948 353668
rect 169820 353612 169876 353668
rect 417676 353612 417732 353668
rect 441308 353612 441364 353668
rect 158620 353276 158676 353332
rect 418012 353276 418068 353332
rect 171276 352604 171332 352660
rect 429212 352604 429268 352660
rect 170828 351932 170884 351988
rect 427868 351932 427924 351988
rect 420924 351260 420980 351316
rect 162540 351036 162596 351092
rect 154476 350924 154532 350980
rect 417564 350924 417620 350980
rect 170940 350588 170996 350644
rect 418236 350588 418292 350644
rect 169148 349916 169204 349972
rect 438956 349916 439012 349972
rect 169036 349244 169092 349300
rect 426412 349244 426468 349300
rect 417900 348684 417956 348740
rect 440188 348684 440244 348740
rect 154364 348572 154420 348628
rect 417564 348572 417620 348628
rect 418236 348572 418292 348628
rect 443324 348572 443380 348628
rect 165676 347900 165732 347956
rect 416668 347900 416724 347956
rect 4172 347452 4228 347508
rect 153692 347340 153748 347396
rect 432908 347340 432964 347396
rect 173740 347228 173796 347284
rect 416780 347228 416836 347284
rect 416668 346892 416724 346948
rect 433132 346892 433188 346948
rect 174076 346556 174132 346612
rect 426300 346556 426356 346612
rect 170604 345884 170660 345940
rect 417676 345884 417732 345940
rect 418012 345324 418068 345380
rect 429324 345324 429380 345380
rect 161084 345212 161140 345268
rect 418236 345212 418292 345268
rect 172396 344540 172452 344596
rect 424396 344540 424452 344596
rect 156044 343868 156100 343924
rect 427756 343868 427812 343924
rect 168812 343756 168868 343812
rect 441308 343756 441364 343812
rect 416780 343532 416836 343588
rect 438172 343532 438228 343588
rect 154252 343196 154308 343252
rect 423276 343196 423332 343252
rect 170716 342524 170772 342580
rect 434812 342524 434868 342580
rect 151004 341852 151060 341908
rect 416668 341852 416724 341908
rect 425964 341852 426020 341908
rect 441644 341852 441700 341908
rect 155932 341180 155988 341236
rect 424284 341180 424340 341236
rect 165564 340508 165620 340564
rect 423164 340508 423220 340564
rect 152348 340284 152404 340340
rect 170940 340284 170996 340340
rect 427980 340284 428036 340340
rect 440300 340284 440356 340340
rect 157164 340172 157220 340228
rect 416668 340172 416724 340228
rect 439068 340172 439124 340228
rect 440188 340172 440244 340228
rect 160860 339836 160916 339892
rect 415996 339836 416052 339892
rect 157612 339164 157668 339220
rect 426188 339164 426244 339220
rect 155820 338492 155876 338548
rect 433020 338492 433076 338548
rect 154140 337820 154196 337876
rect 423052 337820 423108 337876
rect 414092 337708 414148 337764
rect 174076 337148 174132 337204
rect 421484 337148 421540 337204
rect 420924 336812 420980 336868
rect 441532 336812 441588 336868
rect 160412 336588 160468 336644
rect 441196 336588 441252 336644
rect 157500 336476 157556 336532
rect 432908 336476 432964 336532
rect 169820 335804 169876 335860
rect 431004 335804 431060 335860
rect 167356 335132 167412 335188
rect 438284 335132 438340 335188
rect 160748 334460 160804 334516
rect 421372 334460 421428 334516
rect 164220 334348 164276 334404
rect 170492 334348 170548 334404
rect 432796 334348 432852 334404
rect 441308 334348 441364 334404
rect 157388 333788 157444 333844
rect 419468 333788 419524 333844
rect 7532 333116 7588 333172
rect 170492 333116 170548 333172
rect 434700 333116 434756 333172
rect 157052 333004 157108 333060
rect 441644 333004 441700 333060
rect 154028 332444 154084 332500
rect 422940 332444 422996 332500
rect 420812 331884 420868 331940
rect 440748 331884 440804 331940
rect 158844 331772 158900 331828
rect 421260 331772 421316 331828
rect 157276 331100 157332 331156
rect 434588 331100 434644 331156
rect 167244 330428 167300 330484
rect 436492 330428 436548 330484
rect 155708 330092 155764 330148
rect 169820 330092 169876 330148
rect 422492 330092 422548 330148
rect 440860 330092 440916 330148
rect 168924 329756 168980 329812
rect 422716 329756 422772 329812
rect 155036 329420 155092 329476
rect 440188 329420 440244 329476
rect 164108 329196 164164 329252
rect 170716 329196 170772 329252
rect 160636 329084 160692 329140
rect 424508 329084 424564 329140
rect 169820 328412 169876 328468
rect 419356 328412 419412 328468
rect 427644 327740 427700 327796
rect 173068 327292 173124 327348
rect 162428 327068 162484 327124
rect 422604 327068 422660 327124
rect 153804 326396 153860 326452
rect 422828 326396 422884 326452
rect 155596 325836 155652 325892
rect 441084 325836 441140 325892
rect 151116 325724 151172 325780
rect 421036 325724 421092 325780
rect 157164 325276 157220 325332
rect 169820 325276 169876 325332
rect 169820 325052 169876 325108
rect 419244 325052 419300 325108
rect 172284 324380 172340 324436
rect 425964 324380 426020 324436
rect 153692 323708 153748 323764
rect 416668 323708 416724 323764
rect 418236 323484 418292 323540
rect 431116 323484 431172 323540
rect 417788 323372 417844 323428
rect 441196 323372 441252 323428
rect 160412 323036 160468 323092
rect 418012 323036 418068 323092
rect 158732 322364 158788 322420
rect 419580 322364 419636 322420
rect 155372 322252 155428 322308
rect 440972 322252 441028 322308
rect 169932 321692 169988 321748
rect 419132 321692 419188 321748
rect 172172 321020 172228 321076
rect 417788 321020 417844 321076
rect 165452 320348 165508 320404
rect 422492 320348 422548 320404
rect 429436 320124 429492 320180
rect 440188 320124 440244 320180
rect 155484 320012 155540 320068
rect 170492 320012 170548 320068
rect 416668 320012 416724 320068
rect 441084 320012 441140 320068
rect 161980 319676 162036 319732
rect 438844 319676 438900 319732
rect 3388 319004 3444 319060
rect 171164 319004 171220 319060
rect 429436 319004 429492 319060
rect 156828 318668 156884 318724
rect 440188 318668 440244 318724
rect 157052 318444 157108 318500
rect 169820 318444 169876 318500
rect 160972 318332 161028 318388
rect 426076 318332 426132 318388
rect 167132 317660 167188 317716
rect 420812 317660 420868 317716
rect 168812 316988 168868 317044
rect 427980 316988 428036 317044
rect 169820 316316 169876 316372
rect 436380 316316 436436 316372
rect 170716 315644 170772 315700
rect 420924 315644 420980 315700
rect 155148 315084 155204 315140
rect 155596 315084 155652 315140
rect 169932 315084 169988 315140
rect 441308 315084 441364 315140
rect 155372 314972 155428 315028
rect 169820 314972 169876 315028
rect 170940 314972 170996 315028
rect 430892 314972 430948 315028
rect 170492 314300 170548 314356
rect 432796 314300 432852 314356
rect 417564 313292 417620 313348
rect 441644 313292 441700 313348
rect 157836 311500 157892 311556
rect 419020 311500 419076 311556
rect 156940 307916 156996 307972
rect 419916 307916 419972 307972
rect 272188 305676 272244 305732
rect 320684 305676 320740 305732
rect 324156 305676 324212 305732
rect 324604 305676 324660 305732
rect 327292 305676 327348 305732
rect 330428 305676 330484 305732
rect 336476 305676 336532 305732
rect 342524 305676 342580 305732
rect 342972 305676 343028 305732
rect 352380 305676 352436 305732
rect 357756 305676 357812 305732
rect 360892 305676 360948 305732
rect 369404 305676 369460 305732
rect 379596 305676 379652 305732
rect 381052 305676 381108 305732
rect 331548 305564 331604 305620
rect 362684 305564 362740 305620
rect 320012 305452 320068 305508
rect 330876 305452 330932 305508
rect 349580 305452 349636 305508
rect 378812 305452 378868 305508
rect 296492 305340 296548 305396
rect 273980 305228 274036 305284
rect 282604 305228 282660 305284
rect 286300 305228 286356 305284
rect 290668 305228 290724 305284
rect 292348 305228 292404 305284
rect 294140 305228 294196 305284
rect 299068 305228 299124 305284
rect 310828 305228 310884 305284
rect 352828 305340 352884 305396
rect 334236 305116 334292 305172
rect 322588 305004 322644 305060
rect 371084 305228 371140 305284
rect 394492 305228 394548 305284
rect 378812 305116 378868 305172
rect 361900 305004 361956 305060
rect 9212 304892 9268 304948
rect 154476 304892 154532 304948
rect 169372 304892 169428 304948
rect 364588 304892 364644 304948
rect 330988 304780 331044 304836
rect 352828 304780 352884 304836
rect 320796 304668 320852 304724
rect 383068 304668 383124 304724
rect 388444 304668 388500 304724
rect 341404 304556 341460 304612
rect 366268 304556 366324 304612
rect 372988 304556 373044 304612
rect 191772 304444 191828 304500
rect 320012 304444 320068 304500
rect 354396 304444 354452 304500
rect 153916 304332 153972 304388
rect 329196 304332 329252 304388
rect 361900 304332 361956 304388
rect 416108 304332 416164 304388
rect 398076 304220 398132 304276
rect 327740 304108 327796 304164
rect 344652 304108 344708 304164
rect 355852 304108 355908 304164
rect 376460 304108 376516 304164
rect 388444 304108 388500 304164
rect 401548 304108 401604 304164
rect 405244 304108 405300 304164
rect 309148 303996 309204 304052
rect 366268 303996 366324 304052
rect 377580 303996 377636 304052
rect 336028 303884 336084 303940
rect 330988 303660 331044 303716
rect 319004 303324 319060 303380
rect 160524 303212 160580 303268
rect 171164 303212 171220 303268
rect 429436 303212 429492 303268
rect 440972 303212 441028 303268
rect 191772 303100 191828 303156
rect 381388 303100 381444 303156
rect 389900 303100 389956 303156
rect 398412 303100 398468 303156
rect 329196 302876 329252 302932
rect 351036 302876 351092 302932
rect 369516 302876 369572 302932
rect 398076 302876 398132 302932
rect 324492 302764 324548 302820
rect 322588 302540 322644 302596
rect 347788 302540 347844 302596
rect 354396 302540 354452 302596
rect 363468 302428 363524 302484
rect 383068 302428 383124 302484
rect 367612 302316 367668 302372
rect 377580 302316 377636 302372
rect 393148 302204 393204 302260
rect 374332 302092 374388 302148
rect 344316 301980 344372 302036
rect 417452 301868 417508 301924
rect 424620 301868 424676 301924
rect 417676 301756 417732 301812
rect 436716 301756 436772 301812
rect 415996 301644 416052 301700
rect 441420 301644 441476 301700
rect 415772 301532 415828 301588
rect 441756 301532 441812 301588
rect 321692 301420 321748 301476
rect 371084 301420 371140 301476
rect 334236 301308 334292 301364
rect 357756 301308 357812 301364
rect 369516 301308 369572 301364
rect 310828 301084 310884 301140
rect 341404 301084 341460 301140
rect 344428 300972 344484 301028
rect 332556 300860 332612 300916
rect 349580 300860 349636 300916
rect 374556 300860 374612 300916
rect 160300 300748 160356 300804
rect 218428 300748 218484 300804
rect 228732 300748 228788 300804
rect 229180 300748 229236 300804
rect 242172 300748 242228 300804
rect 260540 300748 260596 300804
rect 329420 300748 329476 300804
rect 329868 300748 329924 300804
rect 331548 300748 331604 300804
rect 342636 300748 342692 300804
rect 351372 300748 351428 300804
rect 364812 300748 364868 300804
rect 372428 300748 372484 300804
rect 372988 300748 373044 300804
rect 379708 300748 379764 300804
rect 388108 300748 388164 300804
rect 394828 300748 394884 300804
rect 399756 300748 399812 300804
rect 414988 300748 415044 300804
rect 440748 300748 440804 300804
rect 223356 299516 223412 299572
rect 237692 299516 237748 299572
rect 217980 299404 218036 299460
rect 428540 299404 428596 299460
rect 428428 299180 428484 299236
rect 442988 298956 443044 299012
rect 423724 298844 423780 298900
rect 414092 298732 414148 298788
rect 418012 298732 418068 298788
rect 421148 298732 421204 298788
rect 426748 298620 426804 298676
rect 423612 298508 423668 298564
rect 255612 298284 255668 298340
rect 260092 298284 260148 298340
rect 332332 298284 332388 298340
rect 352716 298284 352772 298340
rect 337708 298172 337764 298228
rect 343532 298172 343588 298228
rect 356188 298172 356244 298228
rect 384972 298284 385028 298340
rect 423388 298284 423444 298340
rect 371084 298172 371140 298228
rect 384860 298172 384916 298228
rect 332332 297948 332388 298004
rect 352716 297948 352772 298004
rect 384972 297948 385028 298004
rect 414092 298060 414148 298116
rect 337708 297836 337764 297892
rect 343532 297836 343588 297892
rect 356188 297836 356244 297892
rect 371084 297836 371140 297892
rect 384860 297836 384916 297892
rect 164220 297164 164276 297220
rect 437388 297164 437444 297220
rect 255612 296940 255668 296996
rect 260092 296828 260148 296884
rect 405244 296716 405300 296772
rect 413980 296604 414036 296660
rect 417788 296604 417844 296660
rect 438060 296604 438116 296660
rect 314972 296492 315028 296548
rect 424508 294812 424564 294868
rect 441308 294812 441364 294868
rect 172620 293580 172676 293636
rect 438396 293580 438452 293636
rect 3500 290780 3556 290836
rect 167468 289996 167524 290052
rect 440860 289996 440916 290052
rect 167692 288988 167748 289044
rect 171052 288988 171108 289044
rect 161196 286412 161252 286468
rect 420700 286412 420756 286468
rect 420476 285628 420532 285684
rect 167580 282828 167636 282884
rect 419804 282828 419860 282884
rect 169260 279244 169316 279300
rect 434924 279244 434980 279300
rect 2492 276668 2548 276724
rect 166124 275660 166180 275716
rect 424620 275660 424676 275716
rect 157724 272076 157780 272132
rect 442540 272076 442596 272132
rect 173180 268492 173236 268548
rect 419692 268492 419748 268548
rect 153916 265468 153972 265524
rect 161980 265468 162036 265524
rect 167692 264908 167748 264964
rect 431228 264908 431284 264964
rect 4172 262556 4228 262612
rect 154476 261324 154532 261380
rect 441196 261324 441252 261380
rect 420588 258636 420644 258692
rect 587132 258188 587188 258244
rect 158508 257740 158564 257796
rect 421596 257740 421652 257796
rect 150892 254156 150948 254212
rect 436604 254156 436660 254212
rect 172508 250572 172564 250628
rect 433244 250572 433300 250628
rect 438844 248556 438900 248612
rect 441196 248556 441252 248612
rect 9884 248444 9940 248500
rect 156156 246988 156212 247044
rect 441756 246988 441812 247044
rect 590492 244972 590548 245028
rect 158620 243404 158676 243460
rect 429324 243404 429380 243460
rect 171388 239820 171444 239876
rect 429212 239820 429268 239876
rect 272972 236796 273028 236852
rect 170828 236236 170884 236292
rect 427868 236236 427924 236292
rect 4284 234332 4340 234388
rect 438284 233436 438340 233492
rect 441756 233436 441812 233492
rect 162540 232652 162596 232708
rect 441532 232652 441588 232708
rect 590716 231868 590772 231924
rect 152348 229068 152404 229124
rect 443324 229068 443380 229124
rect 169148 225484 169204 225540
rect 438956 225484 439012 225540
rect 169036 221900 169092 221956
rect 426412 221900 426468 221956
rect 7756 220220 7812 220276
rect 154364 218316 154420 218372
rect 441644 218316 441700 218372
rect 165676 214732 165732 214788
rect 433132 214732 433188 214788
rect 173740 211148 173796 211204
rect 438172 211148 438228 211204
rect 173964 207564 174020 207620
rect 426300 207564 426356 207620
rect 7980 206108 8036 206164
rect 590604 205324 590660 205380
rect 434812 204988 434868 205044
rect 441532 204988 441588 205044
rect 170604 203980 170660 204036
rect 436716 203980 436772 204036
rect 161084 200396 161140 200452
rect 431116 200396 431172 200452
rect 172396 196812 172452 196868
rect 424396 196812 424452 196868
rect 156044 193228 156100 193284
rect 427756 193228 427812 193284
rect 590828 192108 590884 192164
rect 6188 191996 6244 192052
rect 154252 189644 154308 189700
rect 423276 189644 423332 189700
rect 164108 186060 164164 186116
rect 441532 186060 441588 186116
rect 151004 182476 151060 182532
rect 439068 182476 439124 182532
rect 155932 178892 155988 178948
rect 424284 178892 424340 178948
rect 4396 177884 4452 177940
rect 165564 175308 165620 175364
rect 423164 175308 423220 175364
rect 421484 173852 421540 173908
rect 441532 173852 441588 173908
rect 160860 171724 160916 171780
rect 441420 171724 441476 171780
rect 419580 170492 419636 170548
rect 441420 170492 441476 170548
rect 157612 168140 157668 168196
rect 426188 168140 426244 168196
rect 155820 164556 155876 164612
rect 433020 164556 433076 164612
rect 9436 163772 9492 163828
rect 156044 163772 156100 163828
rect 170940 163772 170996 163828
rect 154140 160972 154196 161028
rect 423052 160972 423108 161028
rect 154364 160412 154420 160468
rect 167356 160412 167412 160468
rect 154140 157948 154196 158004
rect 160972 157948 161028 158004
rect 174076 157388 174132 157444
rect 441532 157388 441588 157444
rect 157500 153804 157556 153860
rect 432908 153804 432964 153860
rect 155708 150220 155764 150276
rect 431004 150220 431060 150276
rect 4508 149660 4564 149716
rect 154364 146636 154420 146692
rect 441756 146636 441812 146692
rect 160748 143052 160804 143108
rect 421372 143052 421428 143108
rect 157388 139468 157444 139524
rect 419468 139468 419524 139524
rect 155484 135884 155540 135940
rect 434700 135884 434756 135940
rect 4620 135548 4676 135604
rect 154252 132412 154308 132468
rect 158844 132412 158900 132468
rect 154028 132300 154084 132356
rect 422940 132300 422996 132356
rect 154252 128716 154308 128772
rect 421260 128716 421316 128772
rect 157276 125132 157332 125188
rect 157500 125132 157556 125188
rect 170716 125132 170772 125188
rect 434588 125132 434644 125188
rect 154476 123452 154532 123508
rect 168924 123452 168980 123508
rect 167244 121548 167300 121604
rect 436492 121548 436548 121604
rect 8204 121436 8260 121492
rect 422716 120092 422772 120148
rect 440188 120092 440244 120148
rect 154476 117964 154532 118020
rect 440188 117964 440244 118020
rect 160636 114380 160692 114436
rect 441308 114380 441364 114436
rect 151116 112588 151172 112644
rect 152908 112588 152964 112644
rect 157164 110796 157220 110852
rect 419356 110796 419412 110852
rect 7644 107324 7700 107380
rect 173068 107212 173124 107268
rect 427644 107212 427700 107268
rect 174636 105196 174692 105252
rect 422828 104972 422884 105028
rect 440188 104972 440244 105028
rect 162428 103628 162484 103684
rect 422604 103628 422660 103684
rect 153804 100044 153860 100100
rect 440188 100044 440244 100100
rect 174748 99484 174804 99540
rect 439964 98252 440020 98308
rect 266476 97692 266532 97748
rect 266252 97580 266308 97636
rect 153804 96572 153860 96628
rect 158732 96572 158788 96628
rect 152908 96460 152964 96516
rect 421036 96460 421092 96516
rect 432684 95788 432740 95844
rect 273980 93996 274036 94052
rect 311612 93324 311668 93380
rect 426860 93324 426916 93380
rect 8988 93212 9044 93268
rect 157052 92876 157108 92932
rect 419244 92876 419300 92932
rect 270620 92764 270676 92820
rect 420700 91644 420756 91700
rect 154476 91532 154532 91588
rect 172284 91532 172340 91588
rect 426972 91532 427028 91588
rect 429212 90972 429268 91028
rect 422044 90300 422100 90356
rect 318332 90188 318388 90244
rect 425068 90188 425124 90244
rect 315084 90076 315140 90132
rect 155484 89852 155540 89908
rect 170492 89852 170548 89908
rect 154476 89292 154532 89348
rect 425964 89292 426020 89348
rect 269612 89068 269668 89124
rect 273308 88508 273364 88564
rect 269724 87948 269780 88004
rect 317436 87948 317492 88004
rect 429660 87948 429716 88004
rect 272972 87836 273028 87892
rect 265244 87724 265300 87780
rect 421932 87724 421988 87780
rect 270284 87612 270340 87668
rect 270620 87500 270676 87556
rect 421484 87052 421540 87108
rect 421036 86940 421092 86996
rect 421708 86828 421764 86884
rect 421820 86716 421876 86772
rect 422268 86492 422324 86548
rect 426076 86492 426132 86548
rect 441644 86492 441700 86548
rect 273532 86268 273588 86324
rect 273084 85932 273140 85988
rect 268380 85820 268436 85876
rect 153692 85708 153748 85764
rect 268828 85708 268884 85764
rect 283836 85708 283892 85764
rect 441084 85708 441140 85764
rect 420812 85036 420868 85092
rect 441532 85036 441588 85092
rect 154252 84812 154308 84868
rect 172172 84812 172228 84868
rect 425740 84140 425796 84196
rect 270844 84028 270900 84084
rect 271068 83916 271124 83972
rect 267932 83692 267988 83748
rect 273196 83692 273252 83748
rect 321692 83356 321748 83412
rect 422156 83356 422212 83412
rect 420924 83244 420980 83300
rect 441308 83244 441364 83300
rect 266588 82684 266644 82740
rect 268940 82348 268996 82404
rect 425628 82236 425684 82292
rect 160412 82124 160468 82180
rect 421148 82124 421204 82180
rect 270172 81788 270228 81844
rect 419132 81452 419188 81508
rect 440412 81452 440468 81508
rect 428316 81228 428372 81284
rect 273644 81116 273700 81172
rect 420812 81116 420868 81172
rect 423836 81004 423892 81060
rect 271292 80892 271348 80948
rect 189532 80556 189588 80612
rect 202524 80556 202580 80612
rect 204876 80556 204932 80612
rect 206556 80556 206612 80612
rect 213948 80556 214004 80612
rect 214844 80556 214900 80612
rect 226604 80556 226660 80612
rect 228396 80556 228452 80612
rect 229964 80556 230020 80612
rect 232092 80556 232148 80612
rect 233436 80556 233492 80612
rect 235116 80556 235172 80612
rect 236796 80556 236852 80612
rect 238476 80556 238532 80612
rect 241836 80556 241892 80612
rect 243516 80556 243572 80612
rect 245196 80556 245252 80612
rect 246876 80556 246932 80612
rect 249564 80556 249620 80612
rect 251916 80556 251972 80612
rect 253484 80556 253540 80612
rect 254716 80556 254772 80612
rect 259644 80556 259700 80612
rect 429436 80556 429492 80612
rect 226716 80444 226772 80500
rect 230076 80444 230132 80500
rect 254492 80444 254548 80500
rect 274092 80444 274148 80500
rect 181468 80220 181524 80276
rect 234780 79772 234836 79828
rect 229964 79660 230020 79716
rect 252924 79660 252980 79716
rect 256956 79660 257012 79716
rect 231420 79548 231476 79604
rect 270508 79548 270564 79604
rect 232764 79436 232820 79492
rect 230748 79324 230804 79380
rect 9660 79100 9716 79156
rect 173852 78988 173908 79044
rect 227388 78988 227444 79044
rect 153804 78540 153860 78596
rect 441420 78540 441476 78596
rect 266700 78428 266756 78484
rect 422492 78316 422548 78372
rect 440188 78316 440244 78372
rect 271516 78204 271572 78260
rect 273420 78204 273476 78260
rect 423948 78204 424004 78260
rect 428204 78092 428260 78148
rect 250908 77308 250964 77364
rect 270620 77196 270676 77252
rect 269836 77084 269892 77140
rect 270620 76860 270676 76916
rect 267820 76748 267876 76804
rect 270508 76748 270564 76804
rect 169596 76412 169652 76468
rect 270620 76300 270676 76356
rect 268828 75404 268884 75460
rect 428652 75404 428708 75460
rect 441084 75404 441140 75460
rect 153692 75292 153748 75348
rect 168812 75292 168868 75348
rect 155596 74956 155652 75012
rect 440412 74956 440468 75012
rect 154028 74732 154084 74788
rect 167132 74732 167188 74788
rect 164556 73948 164612 74004
rect 169708 73948 169764 74004
rect 268940 73836 268996 73892
rect 265916 72604 265972 72660
rect 268828 72044 268884 72100
rect 154252 71372 154308 71428
rect 438060 71372 438116 71428
rect 268940 70700 268996 70756
rect 270060 70700 270116 70756
rect 265916 69356 265972 69412
rect 268828 69132 268884 69188
rect 270060 68460 270116 68516
rect 165452 67900 165508 67956
rect 440188 67788 440244 67844
rect 270060 67564 270116 67620
rect 268828 66668 268884 66724
rect 265916 65996 265972 66052
rect 270060 65324 270116 65380
rect 4732 64988 4788 65044
rect 153916 64204 153972 64260
rect 265916 63980 265972 64036
rect 441196 64204 441252 64260
rect 436380 61292 436436 61348
rect 441196 61292 441252 61348
rect 160524 60620 160580 60676
rect 440972 60620 441028 60676
rect 163996 57932 164052 57988
rect 154140 57036 154196 57092
rect 441644 57036 441700 57092
rect 162316 56140 162372 56196
rect 163884 55244 163940 55300
rect 166012 54348 166068 54404
rect 152012 53564 152068 53620
rect 154028 53452 154084 53508
rect 441532 53452 441588 53508
rect 165788 52556 165844 52612
rect 152124 51660 152180 51716
rect 4844 50876 4900 50932
rect 162204 50764 162260 50820
rect 155372 49868 155428 49924
rect 163772 49868 163828 49924
rect 441196 49868 441252 49924
rect 430892 49532 430948 49588
rect 440972 49532 441028 49588
rect 162092 48972 162148 49028
rect 166236 48076 166292 48132
rect 152236 47852 152292 47908
rect 163660 47852 163716 47908
rect 150780 47180 150836 47236
rect 157500 46284 157556 46340
rect 164556 46284 164612 46340
rect 441308 46284 441364 46340
rect 163660 45388 163716 45444
rect 432796 45276 432852 45332
rect 440188 45276 440244 45332
rect 150556 44492 150612 44548
rect 150332 43596 150388 43652
rect 156044 42700 156100 42756
rect 440972 42700 441028 42756
rect 152012 41804 152068 41860
rect 268828 39788 268884 39844
rect 155484 39116 155540 39172
rect 440188 39116 440244 39172
rect 270060 38444 270116 38500
rect 155372 38220 155428 38276
rect 268828 37772 268884 37828
rect 265916 37100 265972 37156
rect 3388 36876 3444 36932
rect 4956 36764 5012 36820
rect 150332 36428 150388 36484
rect 270060 36204 270116 36260
rect 153692 35532 153748 35588
rect 270060 35532 270116 35588
rect 441084 35532 441140 35588
rect 265916 35084 265972 35140
rect 163548 34636 163604 34692
rect 266140 34412 266196 34468
rect 163772 33740 163828 33796
rect 268828 33068 268884 33124
rect 270060 33068 270116 33124
rect 152236 32844 152292 32900
rect 163884 31948 163940 32004
rect 265916 31724 265972 31780
rect 266140 31500 266196 31556
rect 152124 31052 152180 31108
rect 268940 30380 268996 30436
rect 153692 30156 153748 30212
rect 268828 29932 268884 29988
rect 429436 29372 429492 29428
rect 164108 29260 164164 29316
rect 268828 29036 268884 29092
rect 163996 28364 164052 28420
rect 265916 28364 265972 28420
rect 270060 27692 270116 27748
rect 164220 27468 164276 27524
rect 268940 26796 268996 26852
rect 4172 26572 4228 26628
rect 4508 26572 4564 26628
rect 164332 26572 164388 26628
rect 4508 26348 4564 26404
rect 4732 26348 4788 26404
rect 265916 26348 265972 26404
rect 150444 25676 150500 25732
rect 268828 25228 268884 25284
rect 267036 25004 267092 25060
rect 153916 24780 153972 24836
rect 152348 23884 152404 23940
rect 268940 23660 268996 23716
rect 270060 23660 270116 23716
rect 3500 23436 3556 23492
rect 265468 23100 265524 23156
rect 159740 22988 159796 23044
rect 4956 22652 5012 22708
rect 268828 22316 268884 22372
rect 149772 22092 149828 22148
rect 265916 22092 265972 22148
rect 4060 20972 4116 21028
rect 155372 20972 155428 21028
rect 270060 20972 270116 21028
rect 439068 20972 439124 21028
rect 438844 20860 438900 20916
rect 438620 20748 438676 20804
rect 590604 20748 590660 20804
rect 443212 20636 443268 20692
rect 267036 20524 267092 20580
rect 7756 20076 7812 20132
rect 7532 19964 7588 20020
rect 431228 19964 431284 20020
rect 8204 19852 8260 19908
rect 164108 19852 164164 19908
rect 432460 19852 432516 19908
rect 7980 19740 8036 19796
rect 163548 19740 163604 19796
rect 433020 19740 433076 19796
rect 590716 19740 590772 19796
rect 9212 19628 9268 19684
rect 265916 19628 265972 19684
rect 9660 19516 9716 19572
rect 164332 19516 164388 19572
rect 9436 19404 9492 19460
rect 163884 19404 163940 19460
rect 4844 19292 4900 19348
rect 152348 19292 152404 19348
rect 590492 19292 590548 19348
rect 4284 19180 4340 19236
rect 150332 19180 150388 19236
rect 268940 18956 268996 19012
rect 164556 18508 164612 18564
rect 6188 18396 6244 18452
rect 163772 18396 163828 18452
rect 256956 18396 257012 18452
rect 4956 18284 5012 18340
rect 159740 18284 159796 18340
rect 268940 18284 268996 18340
rect 433356 18284 433412 18340
rect 590828 18284 590884 18340
rect 8988 18172 9044 18228
rect 164220 18172 164276 18228
rect 9884 18060 9940 18116
rect 433132 18060 433188 18116
rect 4620 17948 4676 18004
rect 153692 17948 153748 18004
rect 252812 17948 252868 18004
rect 265020 17948 265076 18004
rect 4732 17836 4788 17892
rect 153916 17836 153972 17892
rect 241724 17836 241780 17892
rect 266924 17836 266980 17892
rect 4396 17724 4452 17780
rect 152236 17724 152292 17780
rect 222460 17724 222516 17780
rect 252028 17724 252084 17780
rect 222908 17612 222964 17668
rect 256844 17612 256900 17668
rect 429212 17612 429268 17668
rect 440076 17612 440132 17668
rect 228844 17500 228900 17556
rect 269052 17500 269108 17556
rect 437836 17500 437892 17556
rect 223132 17388 223188 17444
rect 265468 17388 265524 17444
rect 268828 17388 268884 17444
rect 223356 17276 223412 17332
rect 219548 17164 219604 17220
rect 219548 16828 219604 16884
rect 222460 16828 222516 16884
rect 222908 16828 222964 16884
rect 223356 16828 223412 16884
rect 228844 16828 228900 16884
rect 241724 16828 241780 16884
rect 4172 16716 4228 16772
rect 226268 16716 226324 16772
rect 230748 16716 230804 16772
rect 231196 16716 231252 16772
rect 236572 16716 236628 16772
rect 239260 16716 239316 16772
rect 240380 16716 240436 16772
rect 240604 16716 240660 16772
rect 243740 16716 243796 16772
rect 245084 16716 245140 16772
rect 7644 16604 7700 16660
rect 163996 16604 164052 16660
rect 223132 16604 223188 16660
rect 241948 16604 242004 16660
rect 4396 16492 4452 16548
rect 152124 16492 152180 16548
rect 4508 16380 4564 16436
rect 150444 16380 150500 16436
rect 442652 16716 442708 16772
rect 2492 16268 2548 16324
rect 164556 16268 164612 16324
rect 245308 16268 245364 16324
rect 443100 16156 443156 16212
rect 217308 16044 217364 16100
rect 226044 16044 226100 16100
rect 436492 16044 436548 16100
rect 439964 15932 440020 15988
rect 270060 15820 270116 15876
rect 270508 15148 270564 15204
rect 256844 15036 256900 15092
rect 221340 14924 221396 14980
rect 222236 14924 222292 14980
rect 243068 14924 243124 14980
rect 252028 14588 252084 14644
rect 4172 14364 4228 14420
rect 149772 14364 149828 14420
rect 269724 14364 269780 14420
rect 432908 14364 432964 14420
rect 265916 14252 265972 14308
rect 429660 14252 429716 14308
rect 268156 14140 268212 14196
rect 268604 14140 268660 14196
rect 186844 13356 186900 13412
rect 187068 13356 187124 13412
rect 209468 13356 209524 13412
rect 209692 13356 209748 13412
rect 209916 13356 209972 13412
rect 210140 13356 210196 13412
rect 218652 13356 218708 13412
rect 236124 13356 236180 13412
rect 241500 13356 241556 13412
rect 243516 13356 243572 13412
rect 245980 13356 246036 13412
rect 270620 13356 270676 13412
rect 434364 13244 434420 13300
rect 190428 13132 190484 13188
rect 239148 13132 239204 13188
rect 268604 13132 268660 13188
rect 270620 13132 270676 13188
rect 185724 13020 185780 13076
rect 268716 13020 268772 13076
rect 270508 13020 270564 13076
rect 222012 12908 222068 12964
rect 266812 12908 266868 12964
rect 186396 12796 186452 12852
rect 241052 12796 241108 12852
rect 242396 12796 242452 12852
rect 270620 12796 270676 12852
rect 231420 12684 231476 12740
rect 249452 12684 249508 12740
rect 270396 12684 270452 12740
rect 436716 12684 436772 12740
rect 428316 12572 428372 12628
rect 442876 12572 442932 12628
rect 185052 12460 185108 12516
rect 225036 12348 225092 12404
rect 226604 12348 226660 12404
rect 238476 12348 238532 12404
rect 239148 12348 239204 12404
rect 243292 12348 243348 12404
rect 245196 12348 245252 12404
rect 184940 12236 184996 12292
rect 186172 12236 186228 12292
rect 186508 12236 186564 12292
rect 188188 12236 188244 12292
rect 190428 12236 190484 12292
rect 223356 12236 223412 12292
rect 224924 12236 224980 12292
rect 226716 12236 226772 12292
rect 228396 12236 228452 12292
rect 230076 12236 230132 12292
rect 231644 12236 231700 12292
rect 238364 12236 238420 12292
rect 240156 12236 240212 12292
rect 241724 12236 241780 12292
rect 270172 12236 270228 12292
rect 238588 12124 238644 12180
rect 245084 12124 245140 12180
rect 246876 12124 246932 12180
rect 249452 12124 249508 12180
rect 238364 11788 238420 11844
rect 240156 11788 240212 11844
rect 243404 11788 243460 11844
rect 134428 11228 134484 11284
rect 270284 11228 270340 11284
rect 269164 11004 269220 11060
rect 236796 10780 236852 10836
rect 420476 10444 420532 10500
rect 425740 10444 425796 10500
rect 423948 10332 424004 10388
rect 265468 10108 265524 10164
rect 269500 10108 269556 10164
rect 273868 10108 273924 10164
rect 268156 9996 268212 10052
rect 270284 9996 270340 10052
rect 272972 9884 273028 9940
rect 267148 9660 267204 9716
rect 272076 9660 272132 9716
rect 421036 9548 421092 9604
rect 426972 9436 427028 9492
rect 420700 9324 420756 9380
rect 426748 9212 426804 9268
rect 4172 8764 4228 8820
rect 269724 8540 269780 8596
rect 304108 8428 304164 8484
rect 269276 8316 269332 8372
rect 264572 8204 264628 8260
rect 274092 8204 274148 8260
rect 423724 8204 423780 8260
rect 266476 8092 266532 8148
rect 423612 8092 423668 8148
rect 422044 7980 422100 8036
rect 421484 7868 421540 7924
rect 422268 7756 422324 7812
rect 436268 7644 436324 7700
rect 44492 7532 44548 7588
rect 270508 6972 270564 7028
rect 273308 6860 273364 6916
rect 571228 6748 571284 6804
rect 266252 6636 266308 6692
rect 272972 6636 273028 6692
rect 265244 6300 265300 6356
rect 271628 6300 271684 6356
rect 425628 6300 425684 6356
rect 288988 6188 289044 6244
rect 426860 6188 426916 6244
rect 425068 6076 425124 6132
rect 423500 5852 423556 5908
rect 268044 5068 268100 5124
rect 268492 4956 268548 5012
rect 424172 4844 424228 4900
rect 442764 4844 442820 4900
rect 271516 4732 271572 4788
rect 442988 4732 443044 4788
rect 273196 4620 273252 4676
rect 428428 4508 428484 4564
rect 23436 4284 23492 4340
rect 420588 4284 420644 4340
rect 523516 4284 523572 4340
rect 531132 4284 531188 4340
rect 17276 4172 17332 4228
rect 272188 4172 272244 4228
rect 421932 4172 421988 4228
rect 423836 4172 423892 4228
rect 428540 4172 428596 4228
rect 431788 4172 431844 4228
rect 436828 4172 436884 4228
rect 581308 4172 581364 4228
rect 479724 4060 479780 4116
rect 540652 3948 540708 4004
rect 55356 3836 55412 3892
rect 546364 3836 546420 3892
rect 41804 3724 41860 3780
rect 557788 3724 557844 3780
rect 11564 3388 11620 3444
rect 13356 3388 13412 3444
rect 26796 3388 26852 3444
rect 394044 3388 394100 3444
rect 506380 3388 506436 3444
rect 512092 3388 512148 3444
rect 517804 3388 517860 3444
rect 534940 3388 534996 3444
rect 552636 3388 552692 3444
rect 559692 3388 559748 3444
rect 571228 3388 571284 3444
rect 264684 3276 264740 3332
rect 421820 3276 421876 3332
rect 422156 3052 422212 3108
rect 277228 2492 277284 2548
rect 269836 2044 269892 2100
rect 252812 1708 252868 1764
rect 475916 1708 475972 1764
rect 515900 1708 515956 1764
rect 542668 1708 542724 1764
rect 421708 1596 421764 1652
rect 273084 1484 273140 1540
rect 423388 1484 423444 1540
rect 185612 1148 185668 1204
rect 185612 588 185668 644
rect 474012 588 474068 644
rect 485548 588 485604 644
rect 527324 588 527380 644
rect 533036 588 533092 644
rect 553980 588 554036 644
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect 3388 587188 3444 587198
rect 3388 416724 3444 587132
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect 3388 416658 3444 416668
rect 3500 558964 3556 558974
rect 3500 403284 3556 558908
rect 4172 544852 4228 544862
rect 3500 403218 3556 403228
rect 3948 417844 4004 417854
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect 3948 393988 4004 417788
rect 4172 394100 4228 544796
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 4172 394034 4228 394044
rect 4284 516628 4340 516638
rect 3948 393922 4004 393932
rect 4284 390628 4340 516572
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 4396 502516 4452 502526
rect 4396 394324 4452 502460
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 4396 394258 4452 394268
rect 4508 488404 4564 488414
rect 4284 390562 4340 390572
rect 4508 383908 4564 488348
rect 4732 474292 4788 474302
rect 4620 460180 4676 460190
rect 4620 390740 4676 460124
rect 4620 390674 4676 390684
rect 4732 384020 4788 474236
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 4844 431956 4900 431966
rect 4844 394212 4900 431900
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 4844 394146 4900 394156
rect 4956 403732 5012 403742
rect 4732 383954 4788 383964
rect 4508 383842 4564 383852
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect 4956 372260 5012 403676
rect 4956 372194 5012 372204
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 4284 371476 4340 371486
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect 4172 371364 4228 371374
rect 4172 361620 4228 371308
rect 4172 361554 4228 361564
rect 4284 361228 4340 371420
rect 4172 361172 4340 361228
rect 5418 364350 6038 381922
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 29484 590884 29540 590894
rect 28364 590772 28420 590782
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 26796 590660 26852 590670
rect 26460 575428 26516 575438
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 9138 372094 9758 387922
rect 12572 573076 12628 573086
rect 12572 377300 12628 573020
rect 22448 562350 22768 562384
rect 22448 562294 22518 562350
rect 22574 562294 22642 562350
rect 22698 562294 22768 562350
rect 22448 562226 22768 562294
rect 22448 562170 22518 562226
rect 22574 562170 22642 562226
rect 22698 562170 22768 562226
rect 22448 562102 22768 562170
rect 22448 562046 22518 562102
rect 22574 562046 22642 562102
rect 22698 562046 22768 562102
rect 22448 561978 22768 562046
rect 22448 561922 22518 561978
rect 22574 561922 22642 561978
rect 22698 561922 22768 561978
rect 22448 561888 22768 561922
rect 22448 544350 22768 544384
rect 22448 544294 22518 544350
rect 22574 544294 22642 544350
rect 22698 544294 22768 544350
rect 22448 544226 22768 544294
rect 22448 544170 22518 544226
rect 22574 544170 22642 544226
rect 22698 544170 22768 544226
rect 22448 544102 22768 544170
rect 22448 544046 22518 544102
rect 22574 544046 22642 544102
rect 22698 544046 22768 544102
rect 22448 543978 22768 544046
rect 22448 543922 22518 543978
rect 22574 543922 22642 543978
rect 22698 543922 22768 543978
rect 22448 543888 22768 543922
rect 12572 377234 12628 377244
rect 14252 530740 14308 530750
rect 14252 373828 14308 530684
rect 22448 526350 22768 526384
rect 22448 526294 22518 526350
rect 22574 526294 22642 526350
rect 22698 526294 22768 526350
rect 22448 526226 22768 526294
rect 22448 526170 22518 526226
rect 22574 526170 22642 526226
rect 22698 526170 22768 526226
rect 22448 526102 22768 526170
rect 22448 526046 22518 526102
rect 22574 526046 22642 526102
rect 22698 526046 22768 526102
rect 22448 525978 22768 526046
rect 22448 525922 22518 525978
rect 22574 525922 22642 525978
rect 22698 525922 22768 525978
rect 22448 525888 22768 525922
rect 22448 508350 22768 508384
rect 22448 508294 22518 508350
rect 22574 508294 22642 508350
rect 22698 508294 22768 508350
rect 22448 508226 22768 508294
rect 22448 508170 22518 508226
rect 22574 508170 22642 508226
rect 22698 508170 22768 508226
rect 22448 508102 22768 508170
rect 22448 508046 22518 508102
rect 22574 508046 22642 508102
rect 22698 508046 22768 508102
rect 22448 507978 22768 508046
rect 22448 507922 22518 507978
rect 22574 507922 22642 507978
rect 22698 507922 22768 507978
rect 22448 507888 22768 507922
rect 22448 490350 22768 490384
rect 22448 490294 22518 490350
rect 22574 490294 22642 490350
rect 22698 490294 22768 490350
rect 22448 490226 22768 490294
rect 22448 490170 22518 490226
rect 22574 490170 22642 490226
rect 22698 490170 22768 490226
rect 22448 490102 22768 490170
rect 22448 490046 22518 490102
rect 22574 490046 22642 490102
rect 22698 490046 22768 490102
rect 22448 489978 22768 490046
rect 22448 489922 22518 489978
rect 22574 489922 22642 489978
rect 22698 489922 22768 489978
rect 22448 489888 22768 489922
rect 22448 472350 22768 472384
rect 22448 472294 22518 472350
rect 22574 472294 22642 472350
rect 22698 472294 22768 472350
rect 22448 472226 22768 472294
rect 22448 472170 22518 472226
rect 22574 472170 22642 472226
rect 22698 472170 22768 472226
rect 22448 472102 22768 472170
rect 22448 472046 22518 472102
rect 22574 472046 22642 472102
rect 22698 472046 22768 472102
rect 22448 471978 22768 472046
rect 22448 471922 22518 471978
rect 22574 471922 22642 471978
rect 22698 471922 22768 471978
rect 22448 471888 22768 471922
rect 22448 454350 22768 454384
rect 22448 454294 22518 454350
rect 22574 454294 22642 454350
rect 22698 454294 22768 454350
rect 22448 454226 22768 454294
rect 22448 454170 22518 454226
rect 22574 454170 22642 454226
rect 22698 454170 22768 454226
rect 22448 454102 22768 454170
rect 22448 454046 22518 454102
rect 22574 454046 22642 454102
rect 22698 454046 22768 454102
rect 22448 453978 22768 454046
rect 22448 453922 22518 453978
rect 22574 453922 22642 453978
rect 22698 453922 22768 453978
rect 22448 453888 22768 453922
rect 14252 373762 14308 373772
rect 17612 446068 17668 446078
rect 17612 372148 17668 446012
rect 22448 436350 22768 436384
rect 22448 436294 22518 436350
rect 22574 436294 22642 436350
rect 22698 436294 22768 436350
rect 22448 436226 22768 436294
rect 22448 436170 22518 436226
rect 22574 436170 22642 436226
rect 22698 436170 22768 436226
rect 22448 436102 22768 436170
rect 22448 436046 22518 436102
rect 22574 436046 22642 436102
rect 22698 436046 22768 436102
rect 22448 435978 22768 436046
rect 22448 435922 22518 435978
rect 22574 435922 22642 435978
rect 22698 435922 22768 435978
rect 22448 435888 22768 435922
rect 22448 418350 22768 418384
rect 22448 418294 22518 418350
rect 22574 418294 22642 418350
rect 22698 418294 22768 418350
rect 22448 418226 22768 418294
rect 22448 418170 22518 418226
rect 22574 418170 22642 418226
rect 22698 418170 22768 418226
rect 22448 418102 22768 418170
rect 22448 418046 22518 418102
rect 22574 418046 22642 418102
rect 22698 418046 22768 418102
rect 22448 417978 22768 418046
rect 22448 417922 22518 417978
rect 22574 417922 22642 417978
rect 22698 417922 22768 417978
rect 22448 417888 22768 417922
rect 22448 400350 22768 400384
rect 22448 400294 22518 400350
rect 22574 400294 22642 400350
rect 22698 400294 22768 400350
rect 22448 400226 22768 400294
rect 22448 400170 22518 400226
rect 22574 400170 22642 400226
rect 22698 400170 22768 400226
rect 22448 400102 22768 400170
rect 22448 400046 22518 400102
rect 22574 400046 22642 400102
rect 22698 400046 22768 400102
rect 22448 399978 22768 400046
rect 22448 399922 22518 399978
rect 22574 399922 22642 399978
rect 22698 399922 22768 399978
rect 22448 399888 22768 399922
rect 26460 393092 26516 575372
rect 26460 393026 26516 393036
rect 26572 575092 26628 575102
rect 26572 389844 26628 575036
rect 26572 389778 26628 389788
rect 26684 574532 26740 574542
rect 26684 389732 26740 574476
rect 26684 389666 26740 389676
rect 26796 373940 26852 590604
rect 28028 576100 28084 576110
rect 28028 394548 28084 576044
rect 28028 394482 28084 394492
rect 28140 575764 28196 575774
rect 28140 393204 28196 575708
rect 28140 393138 28196 393148
rect 28252 575540 28308 575550
rect 28252 377412 28308 575484
rect 28252 377346 28308 377356
rect 28364 374052 28420 590716
rect 28364 373986 28420 373996
rect 28476 590548 28532 590558
rect 26796 373874 26852 373884
rect 28476 372372 28532 590492
rect 29372 577332 29428 577342
rect 29260 575988 29316 575998
rect 29148 575876 29204 575886
rect 29036 575652 29092 575662
rect 29036 389508 29092 575596
rect 29148 389732 29204 575820
rect 29148 389666 29204 389676
rect 29036 389442 29092 389452
rect 29260 383012 29316 575932
rect 29260 382946 29316 382956
rect 29372 374612 29428 577276
rect 29484 375620 29540 590828
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 189738 575846 190358 579922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 575846 194078 585922
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 220458 575846 221078 579922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 575846 224798 585922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 251178 575846 251798 579922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 575846 255518 585922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 281898 575846 282518 579922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 575846 286238 585922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 312618 575846 313238 579922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 575846 316958 585922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 343338 575846 343958 579922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 575846 347678 585922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 374058 575846 374678 579922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 575846 378398 585922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 404778 575846 405398 579922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 575846 409118 585922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 435498 575846 436118 579922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 575846 439838 585922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 466218 575846 466838 579922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 575846 470558 585922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 496938 575846 497558 579922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 575846 501278 585922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 527658 575846 528278 579922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 549388 591108 549444 591118
rect 548044 590996 548100 591006
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 575846 531998 585922
rect 547708 590772 547764 590782
rect 37808 568350 38128 568384
rect 37808 568294 37878 568350
rect 37934 568294 38002 568350
rect 38058 568294 38128 568350
rect 37808 568226 38128 568294
rect 37808 568170 37878 568226
rect 37934 568170 38002 568226
rect 38058 568170 38128 568226
rect 37808 568102 38128 568170
rect 37808 568046 37878 568102
rect 37934 568046 38002 568102
rect 38058 568046 38128 568102
rect 37808 567978 38128 568046
rect 37808 567922 37878 567978
rect 37934 567922 38002 567978
rect 38058 567922 38128 567978
rect 37808 567888 38128 567922
rect 68528 568350 68848 568384
rect 68528 568294 68598 568350
rect 68654 568294 68722 568350
rect 68778 568294 68848 568350
rect 68528 568226 68848 568294
rect 68528 568170 68598 568226
rect 68654 568170 68722 568226
rect 68778 568170 68848 568226
rect 68528 568102 68848 568170
rect 68528 568046 68598 568102
rect 68654 568046 68722 568102
rect 68778 568046 68848 568102
rect 68528 567978 68848 568046
rect 68528 567922 68598 567978
rect 68654 567922 68722 567978
rect 68778 567922 68848 567978
rect 68528 567888 68848 567922
rect 99248 568350 99568 568384
rect 99248 568294 99318 568350
rect 99374 568294 99442 568350
rect 99498 568294 99568 568350
rect 99248 568226 99568 568294
rect 99248 568170 99318 568226
rect 99374 568170 99442 568226
rect 99498 568170 99568 568226
rect 99248 568102 99568 568170
rect 99248 568046 99318 568102
rect 99374 568046 99442 568102
rect 99498 568046 99568 568102
rect 99248 567978 99568 568046
rect 99248 567922 99318 567978
rect 99374 567922 99442 567978
rect 99498 567922 99568 567978
rect 99248 567888 99568 567922
rect 129968 568350 130288 568384
rect 129968 568294 130038 568350
rect 130094 568294 130162 568350
rect 130218 568294 130288 568350
rect 129968 568226 130288 568294
rect 129968 568170 130038 568226
rect 130094 568170 130162 568226
rect 130218 568170 130288 568226
rect 129968 568102 130288 568170
rect 129968 568046 130038 568102
rect 130094 568046 130162 568102
rect 130218 568046 130288 568102
rect 129968 567978 130288 568046
rect 129968 567922 130038 567978
rect 130094 567922 130162 567978
rect 130218 567922 130288 567978
rect 129968 567888 130288 567922
rect 160688 568350 161008 568384
rect 160688 568294 160758 568350
rect 160814 568294 160882 568350
rect 160938 568294 161008 568350
rect 160688 568226 161008 568294
rect 160688 568170 160758 568226
rect 160814 568170 160882 568226
rect 160938 568170 161008 568226
rect 160688 568102 161008 568170
rect 160688 568046 160758 568102
rect 160814 568046 160882 568102
rect 160938 568046 161008 568102
rect 160688 567978 161008 568046
rect 160688 567922 160758 567978
rect 160814 567922 160882 567978
rect 160938 567922 161008 567978
rect 160688 567888 161008 567922
rect 191408 568350 191728 568384
rect 191408 568294 191478 568350
rect 191534 568294 191602 568350
rect 191658 568294 191728 568350
rect 191408 568226 191728 568294
rect 191408 568170 191478 568226
rect 191534 568170 191602 568226
rect 191658 568170 191728 568226
rect 191408 568102 191728 568170
rect 191408 568046 191478 568102
rect 191534 568046 191602 568102
rect 191658 568046 191728 568102
rect 191408 567978 191728 568046
rect 191408 567922 191478 567978
rect 191534 567922 191602 567978
rect 191658 567922 191728 567978
rect 191408 567888 191728 567922
rect 222128 568350 222448 568384
rect 222128 568294 222198 568350
rect 222254 568294 222322 568350
rect 222378 568294 222448 568350
rect 222128 568226 222448 568294
rect 222128 568170 222198 568226
rect 222254 568170 222322 568226
rect 222378 568170 222448 568226
rect 222128 568102 222448 568170
rect 222128 568046 222198 568102
rect 222254 568046 222322 568102
rect 222378 568046 222448 568102
rect 222128 567978 222448 568046
rect 222128 567922 222198 567978
rect 222254 567922 222322 567978
rect 222378 567922 222448 567978
rect 222128 567888 222448 567922
rect 252848 568350 253168 568384
rect 252848 568294 252918 568350
rect 252974 568294 253042 568350
rect 253098 568294 253168 568350
rect 252848 568226 253168 568294
rect 252848 568170 252918 568226
rect 252974 568170 253042 568226
rect 253098 568170 253168 568226
rect 252848 568102 253168 568170
rect 252848 568046 252918 568102
rect 252974 568046 253042 568102
rect 253098 568046 253168 568102
rect 252848 567978 253168 568046
rect 252848 567922 252918 567978
rect 252974 567922 253042 567978
rect 253098 567922 253168 567978
rect 252848 567888 253168 567922
rect 283568 568350 283888 568384
rect 283568 568294 283638 568350
rect 283694 568294 283762 568350
rect 283818 568294 283888 568350
rect 283568 568226 283888 568294
rect 283568 568170 283638 568226
rect 283694 568170 283762 568226
rect 283818 568170 283888 568226
rect 283568 568102 283888 568170
rect 283568 568046 283638 568102
rect 283694 568046 283762 568102
rect 283818 568046 283888 568102
rect 283568 567978 283888 568046
rect 283568 567922 283638 567978
rect 283694 567922 283762 567978
rect 283818 567922 283888 567978
rect 283568 567888 283888 567922
rect 314288 568350 314608 568384
rect 314288 568294 314358 568350
rect 314414 568294 314482 568350
rect 314538 568294 314608 568350
rect 314288 568226 314608 568294
rect 314288 568170 314358 568226
rect 314414 568170 314482 568226
rect 314538 568170 314608 568226
rect 314288 568102 314608 568170
rect 314288 568046 314358 568102
rect 314414 568046 314482 568102
rect 314538 568046 314608 568102
rect 314288 567978 314608 568046
rect 314288 567922 314358 567978
rect 314414 567922 314482 567978
rect 314538 567922 314608 567978
rect 314288 567888 314608 567922
rect 345008 568350 345328 568384
rect 345008 568294 345078 568350
rect 345134 568294 345202 568350
rect 345258 568294 345328 568350
rect 345008 568226 345328 568294
rect 345008 568170 345078 568226
rect 345134 568170 345202 568226
rect 345258 568170 345328 568226
rect 345008 568102 345328 568170
rect 345008 568046 345078 568102
rect 345134 568046 345202 568102
rect 345258 568046 345328 568102
rect 345008 567978 345328 568046
rect 345008 567922 345078 567978
rect 345134 567922 345202 567978
rect 345258 567922 345328 567978
rect 345008 567888 345328 567922
rect 375728 568350 376048 568384
rect 375728 568294 375798 568350
rect 375854 568294 375922 568350
rect 375978 568294 376048 568350
rect 375728 568226 376048 568294
rect 375728 568170 375798 568226
rect 375854 568170 375922 568226
rect 375978 568170 376048 568226
rect 375728 568102 376048 568170
rect 375728 568046 375798 568102
rect 375854 568046 375922 568102
rect 375978 568046 376048 568102
rect 375728 567978 376048 568046
rect 375728 567922 375798 567978
rect 375854 567922 375922 567978
rect 375978 567922 376048 567978
rect 375728 567888 376048 567922
rect 406448 568350 406768 568384
rect 406448 568294 406518 568350
rect 406574 568294 406642 568350
rect 406698 568294 406768 568350
rect 406448 568226 406768 568294
rect 406448 568170 406518 568226
rect 406574 568170 406642 568226
rect 406698 568170 406768 568226
rect 406448 568102 406768 568170
rect 406448 568046 406518 568102
rect 406574 568046 406642 568102
rect 406698 568046 406768 568102
rect 406448 567978 406768 568046
rect 406448 567922 406518 567978
rect 406574 567922 406642 567978
rect 406698 567922 406768 567978
rect 406448 567888 406768 567922
rect 437168 568350 437488 568384
rect 437168 568294 437238 568350
rect 437294 568294 437362 568350
rect 437418 568294 437488 568350
rect 437168 568226 437488 568294
rect 437168 568170 437238 568226
rect 437294 568170 437362 568226
rect 437418 568170 437488 568226
rect 437168 568102 437488 568170
rect 437168 568046 437238 568102
rect 437294 568046 437362 568102
rect 437418 568046 437488 568102
rect 437168 567978 437488 568046
rect 437168 567922 437238 567978
rect 437294 567922 437362 567978
rect 437418 567922 437488 567978
rect 437168 567888 437488 567922
rect 467888 568350 468208 568384
rect 467888 568294 467958 568350
rect 468014 568294 468082 568350
rect 468138 568294 468208 568350
rect 467888 568226 468208 568294
rect 467888 568170 467958 568226
rect 468014 568170 468082 568226
rect 468138 568170 468208 568226
rect 467888 568102 468208 568170
rect 467888 568046 467958 568102
rect 468014 568046 468082 568102
rect 468138 568046 468208 568102
rect 467888 567978 468208 568046
rect 467888 567922 467958 567978
rect 468014 567922 468082 567978
rect 468138 567922 468208 567978
rect 467888 567888 468208 567922
rect 498608 568350 498928 568384
rect 498608 568294 498678 568350
rect 498734 568294 498802 568350
rect 498858 568294 498928 568350
rect 498608 568226 498928 568294
rect 498608 568170 498678 568226
rect 498734 568170 498802 568226
rect 498858 568170 498928 568226
rect 498608 568102 498928 568170
rect 498608 568046 498678 568102
rect 498734 568046 498802 568102
rect 498858 568046 498928 568102
rect 498608 567978 498928 568046
rect 498608 567922 498678 567978
rect 498734 567922 498802 567978
rect 498858 567922 498928 567978
rect 498608 567888 498928 567922
rect 529328 568350 529648 568384
rect 529328 568294 529398 568350
rect 529454 568294 529522 568350
rect 529578 568294 529648 568350
rect 529328 568226 529648 568294
rect 529328 568170 529398 568226
rect 529454 568170 529522 568226
rect 529578 568170 529648 568226
rect 529328 568102 529648 568170
rect 529328 568046 529398 568102
rect 529454 568046 529522 568102
rect 529578 568046 529648 568102
rect 529328 567978 529648 568046
rect 529328 567922 529398 567978
rect 529454 567922 529522 567978
rect 529578 567922 529648 567978
rect 529328 567888 529648 567922
rect 53168 562350 53488 562384
rect 53168 562294 53238 562350
rect 53294 562294 53362 562350
rect 53418 562294 53488 562350
rect 53168 562226 53488 562294
rect 53168 562170 53238 562226
rect 53294 562170 53362 562226
rect 53418 562170 53488 562226
rect 53168 562102 53488 562170
rect 53168 562046 53238 562102
rect 53294 562046 53362 562102
rect 53418 562046 53488 562102
rect 53168 561978 53488 562046
rect 53168 561922 53238 561978
rect 53294 561922 53362 561978
rect 53418 561922 53488 561978
rect 53168 561888 53488 561922
rect 83888 562350 84208 562384
rect 83888 562294 83958 562350
rect 84014 562294 84082 562350
rect 84138 562294 84208 562350
rect 83888 562226 84208 562294
rect 83888 562170 83958 562226
rect 84014 562170 84082 562226
rect 84138 562170 84208 562226
rect 83888 562102 84208 562170
rect 83888 562046 83958 562102
rect 84014 562046 84082 562102
rect 84138 562046 84208 562102
rect 83888 561978 84208 562046
rect 83888 561922 83958 561978
rect 84014 561922 84082 561978
rect 84138 561922 84208 561978
rect 83888 561888 84208 561922
rect 114608 562350 114928 562384
rect 114608 562294 114678 562350
rect 114734 562294 114802 562350
rect 114858 562294 114928 562350
rect 114608 562226 114928 562294
rect 114608 562170 114678 562226
rect 114734 562170 114802 562226
rect 114858 562170 114928 562226
rect 114608 562102 114928 562170
rect 114608 562046 114678 562102
rect 114734 562046 114802 562102
rect 114858 562046 114928 562102
rect 114608 561978 114928 562046
rect 114608 561922 114678 561978
rect 114734 561922 114802 561978
rect 114858 561922 114928 561978
rect 114608 561888 114928 561922
rect 145328 562350 145648 562384
rect 145328 562294 145398 562350
rect 145454 562294 145522 562350
rect 145578 562294 145648 562350
rect 145328 562226 145648 562294
rect 145328 562170 145398 562226
rect 145454 562170 145522 562226
rect 145578 562170 145648 562226
rect 145328 562102 145648 562170
rect 145328 562046 145398 562102
rect 145454 562046 145522 562102
rect 145578 562046 145648 562102
rect 145328 561978 145648 562046
rect 145328 561922 145398 561978
rect 145454 561922 145522 561978
rect 145578 561922 145648 561978
rect 145328 561888 145648 561922
rect 176048 562350 176368 562384
rect 176048 562294 176118 562350
rect 176174 562294 176242 562350
rect 176298 562294 176368 562350
rect 176048 562226 176368 562294
rect 176048 562170 176118 562226
rect 176174 562170 176242 562226
rect 176298 562170 176368 562226
rect 176048 562102 176368 562170
rect 176048 562046 176118 562102
rect 176174 562046 176242 562102
rect 176298 562046 176368 562102
rect 176048 561978 176368 562046
rect 176048 561922 176118 561978
rect 176174 561922 176242 561978
rect 176298 561922 176368 561978
rect 176048 561888 176368 561922
rect 206768 562350 207088 562384
rect 206768 562294 206838 562350
rect 206894 562294 206962 562350
rect 207018 562294 207088 562350
rect 206768 562226 207088 562294
rect 206768 562170 206838 562226
rect 206894 562170 206962 562226
rect 207018 562170 207088 562226
rect 206768 562102 207088 562170
rect 206768 562046 206838 562102
rect 206894 562046 206962 562102
rect 207018 562046 207088 562102
rect 206768 561978 207088 562046
rect 206768 561922 206838 561978
rect 206894 561922 206962 561978
rect 207018 561922 207088 561978
rect 206768 561888 207088 561922
rect 237488 562350 237808 562384
rect 237488 562294 237558 562350
rect 237614 562294 237682 562350
rect 237738 562294 237808 562350
rect 237488 562226 237808 562294
rect 237488 562170 237558 562226
rect 237614 562170 237682 562226
rect 237738 562170 237808 562226
rect 237488 562102 237808 562170
rect 237488 562046 237558 562102
rect 237614 562046 237682 562102
rect 237738 562046 237808 562102
rect 237488 561978 237808 562046
rect 237488 561922 237558 561978
rect 237614 561922 237682 561978
rect 237738 561922 237808 561978
rect 237488 561888 237808 561922
rect 268208 562350 268528 562384
rect 268208 562294 268278 562350
rect 268334 562294 268402 562350
rect 268458 562294 268528 562350
rect 268208 562226 268528 562294
rect 268208 562170 268278 562226
rect 268334 562170 268402 562226
rect 268458 562170 268528 562226
rect 268208 562102 268528 562170
rect 268208 562046 268278 562102
rect 268334 562046 268402 562102
rect 268458 562046 268528 562102
rect 268208 561978 268528 562046
rect 268208 561922 268278 561978
rect 268334 561922 268402 561978
rect 268458 561922 268528 561978
rect 268208 561888 268528 561922
rect 298928 562350 299248 562384
rect 298928 562294 298998 562350
rect 299054 562294 299122 562350
rect 299178 562294 299248 562350
rect 298928 562226 299248 562294
rect 298928 562170 298998 562226
rect 299054 562170 299122 562226
rect 299178 562170 299248 562226
rect 298928 562102 299248 562170
rect 298928 562046 298998 562102
rect 299054 562046 299122 562102
rect 299178 562046 299248 562102
rect 298928 561978 299248 562046
rect 298928 561922 298998 561978
rect 299054 561922 299122 561978
rect 299178 561922 299248 561978
rect 298928 561888 299248 561922
rect 329648 562350 329968 562384
rect 329648 562294 329718 562350
rect 329774 562294 329842 562350
rect 329898 562294 329968 562350
rect 329648 562226 329968 562294
rect 329648 562170 329718 562226
rect 329774 562170 329842 562226
rect 329898 562170 329968 562226
rect 329648 562102 329968 562170
rect 329648 562046 329718 562102
rect 329774 562046 329842 562102
rect 329898 562046 329968 562102
rect 329648 561978 329968 562046
rect 329648 561922 329718 561978
rect 329774 561922 329842 561978
rect 329898 561922 329968 561978
rect 329648 561888 329968 561922
rect 360368 562350 360688 562384
rect 360368 562294 360438 562350
rect 360494 562294 360562 562350
rect 360618 562294 360688 562350
rect 360368 562226 360688 562294
rect 360368 562170 360438 562226
rect 360494 562170 360562 562226
rect 360618 562170 360688 562226
rect 360368 562102 360688 562170
rect 360368 562046 360438 562102
rect 360494 562046 360562 562102
rect 360618 562046 360688 562102
rect 360368 561978 360688 562046
rect 360368 561922 360438 561978
rect 360494 561922 360562 561978
rect 360618 561922 360688 561978
rect 360368 561888 360688 561922
rect 391088 562350 391408 562384
rect 391088 562294 391158 562350
rect 391214 562294 391282 562350
rect 391338 562294 391408 562350
rect 391088 562226 391408 562294
rect 391088 562170 391158 562226
rect 391214 562170 391282 562226
rect 391338 562170 391408 562226
rect 391088 562102 391408 562170
rect 391088 562046 391158 562102
rect 391214 562046 391282 562102
rect 391338 562046 391408 562102
rect 391088 561978 391408 562046
rect 391088 561922 391158 561978
rect 391214 561922 391282 561978
rect 391338 561922 391408 561978
rect 391088 561888 391408 561922
rect 421808 562350 422128 562384
rect 421808 562294 421878 562350
rect 421934 562294 422002 562350
rect 422058 562294 422128 562350
rect 421808 562226 422128 562294
rect 421808 562170 421878 562226
rect 421934 562170 422002 562226
rect 422058 562170 422128 562226
rect 421808 562102 422128 562170
rect 421808 562046 421878 562102
rect 421934 562046 422002 562102
rect 422058 562046 422128 562102
rect 421808 561978 422128 562046
rect 421808 561922 421878 561978
rect 421934 561922 422002 561978
rect 422058 561922 422128 561978
rect 421808 561888 422128 561922
rect 452528 562350 452848 562384
rect 452528 562294 452598 562350
rect 452654 562294 452722 562350
rect 452778 562294 452848 562350
rect 452528 562226 452848 562294
rect 452528 562170 452598 562226
rect 452654 562170 452722 562226
rect 452778 562170 452848 562226
rect 452528 562102 452848 562170
rect 452528 562046 452598 562102
rect 452654 562046 452722 562102
rect 452778 562046 452848 562102
rect 452528 561978 452848 562046
rect 452528 561922 452598 561978
rect 452654 561922 452722 561978
rect 452778 561922 452848 561978
rect 452528 561888 452848 561922
rect 483248 562350 483568 562384
rect 483248 562294 483318 562350
rect 483374 562294 483442 562350
rect 483498 562294 483568 562350
rect 483248 562226 483568 562294
rect 483248 562170 483318 562226
rect 483374 562170 483442 562226
rect 483498 562170 483568 562226
rect 483248 562102 483568 562170
rect 483248 562046 483318 562102
rect 483374 562046 483442 562102
rect 483498 562046 483568 562102
rect 483248 561978 483568 562046
rect 483248 561922 483318 561978
rect 483374 561922 483442 561978
rect 483498 561922 483568 561978
rect 483248 561888 483568 561922
rect 513968 562350 514288 562384
rect 513968 562294 514038 562350
rect 514094 562294 514162 562350
rect 514218 562294 514288 562350
rect 513968 562226 514288 562294
rect 513968 562170 514038 562226
rect 514094 562170 514162 562226
rect 514218 562170 514288 562226
rect 513968 562102 514288 562170
rect 513968 562046 514038 562102
rect 514094 562046 514162 562102
rect 514218 562046 514288 562102
rect 513968 561978 514288 562046
rect 513968 561922 514038 561978
rect 514094 561922 514162 561978
rect 514218 561922 514288 561978
rect 513968 561888 514288 561922
rect 544688 562350 545008 562384
rect 544688 562294 544758 562350
rect 544814 562294 544882 562350
rect 544938 562294 545008 562350
rect 544688 562226 545008 562294
rect 544688 562170 544758 562226
rect 544814 562170 544882 562226
rect 544938 562170 545008 562226
rect 544688 562102 545008 562170
rect 544688 562046 544758 562102
rect 544814 562046 544882 562102
rect 544938 562046 545008 562102
rect 544688 561978 545008 562046
rect 544688 561922 544758 561978
rect 544814 561922 544882 561978
rect 544938 561922 545008 561978
rect 544688 561888 545008 561922
rect 37808 550350 38128 550384
rect 37808 550294 37878 550350
rect 37934 550294 38002 550350
rect 38058 550294 38128 550350
rect 37808 550226 38128 550294
rect 37808 550170 37878 550226
rect 37934 550170 38002 550226
rect 38058 550170 38128 550226
rect 37808 550102 38128 550170
rect 37808 550046 37878 550102
rect 37934 550046 38002 550102
rect 38058 550046 38128 550102
rect 37808 549978 38128 550046
rect 37808 549922 37878 549978
rect 37934 549922 38002 549978
rect 38058 549922 38128 549978
rect 37808 549888 38128 549922
rect 68528 550350 68848 550384
rect 68528 550294 68598 550350
rect 68654 550294 68722 550350
rect 68778 550294 68848 550350
rect 68528 550226 68848 550294
rect 68528 550170 68598 550226
rect 68654 550170 68722 550226
rect 68778 550170 68848 550226
rect 68528 550102 68848 550170
rect 68528 550046 68598 550102
rect 68654 550046 68722 550102
rect 68778 550046 68848 550102
rect 68528 549978 68848 550046
rect 68528 549922 68598 549978
rect 68654 549922 68722 549978
rect 68778 549922 68848 549978
rect 68528 549888 68848 549922
rect 99248 550350 99568 550384
rect 99248 550294 99318 550350
rect 99374 550294 99442 550350
rect 99498 550294 99568 550350
rect 99248 550226 99568 550294
rect 99248 550170 99318 550226
rect 99374 550170 99442 550226
rect 99498 550170 99568 550226
rect 99248 550102 99568 550170
rect 99248 550046 99318 550102
rect 99374 550046 99442 550102
rect 99498 550046 99568 550102
rect 99248 549978 99568 550046
rect 99248 549922 99318 549978
rect 99374 549922 99442 549978
rect 99498 549922 99568 549978
rect 99248 549888 99568 549922
rect 129968 550350 130288 550384
rect 129968 550294 130038 550350
rect 130094 550294 130162 550350
rect 130218 550294 130288 550350
rect 129968 550226 130288 550294
rect 129968 550170 130038 550226
rect 130094 550170 130162 550226
rect 130218 550170 130288 550226
rect 129968 550102 130288 550170
rect 129968 550046 130038 550102
rect 130094 550046 130162 550102
rect 130218 550046 130288 550102
rect 129968 549978 130288 550046
rect 129968 549922 130038 549978
rect 130094 549922 130162 549978
rect 130218 549922 130288 549978
rect 129968 549888 130288 549922
rect 160688 550350 161008 550384
rect 160688 550294 160758 550350
rect 160814 550294 160882 550350
rect 160938 550294 161008 550350
rect 160688 550226 161008 550294
rect 160688 550170 160758 550226
rect 160814 550170 160882 550226
rect 160938 550170 161008 550226
rect 160688 550102 161008 550170
rect 160688 550046 160758 550102
rect 160814 550046 160882 550102
rect 160938 550046 161008 550102
rect 160688 549978 161008 550046
rect 160688 549922 160758 549978
rect 160814 549922 160882 549978
rect 160938 549922 161008 549978
rect 160688 549888 161008 549922
rect 191408 550350 191728 550384
rect 191408 550294 191478 550350
rect 191534 550294 191602 550350
rect 191658 550294 191728 550350
rect 191408 550226 191728 550294
rect 191408 550170 191478 550226
rect 191534 550170 191602 550226
rect 191658 550170 191728 550226
rect 191408 550102 191728 550170
rect 191408 550046 191478 550102
rect 191534 550046 191602 550102
rect 191658 550046 191728 550102
rect 191408 549978 191728 550046
rect 191408 549922 191478 549978
rect 191534 549922 191602 549978
rect 191658 549922 191728 549978
rect 191408 549888 191728 549922
rect 222128 550350 222448 550384
rect 222128 550294 222198 550350
rect 222254 550294 222322 550350
rect 222378 550294 222448 550350
rect 222128 550226 222448 550294
rect 222128 550170 222198 550226
rect 222254 550170 222322 550226
rect 222378 550170 222448 550226
rect 222128 550102 222448 550170
rect 222128 550046 222198 550102
rect 222254 550046 222322 550102
rect 222378 550046 222448 550102
rect 222128 549978 222448 550046
rect 222128 549922 222198 549978
rect 222254 549922 222322 549978
rect 222378 549922 222448 549978
rect 222128 549888 222448 549922
rect 252848 550350 253168 550384
rect 252848 550294 252918 550350
rect 252974 550294 253042 550350
rect 253098 550294 253168 550350
rect 252848 550226 253168 550294
rect 252848 550170 252918 550226
rect 252974 550170 253042 550226
rect 253098 550170 253168 550226
rect 252848 550102 253168 550170
rect 252848 550046 252918 550102
rect 252974 550046 253042 550102
rect 253098 550046 253168 550102
rect 252848 549978 253168 550046
rect 252848 549922 252918 549978
rect 252974 549922 253042 549978
rect 253098 549922 253168 549978
rect 252848 549888 253168 549922
rect 283568 550350 283888 550384
rect 283568 550294 283638 550350
rect 283694 550294 283762 550350
rect 283818 550294 283888 550350
rect 283568 550226 283888 550294
rect 283568 550170 283638 550226
rect 283694 550170 283762 550226
rect 283818 550170 283888 550226
rect 283568 550102 283888 550170
rect 283568 550046 283638 550102
rect 283694 550046 283762 550102
rect 283818 550046 283888 550102
rect 283568 549978 283888 550046
rect 283568 549922 283638 549978
rect 283694 549922 283762 549978
rect 283818 549922 283888 549978
rect 283568 549888 283888 549922
rect 314288 550350 314608 550384
rect 314288 550294 314358 550350
rect 314414 550294 314482 550350
rect 314538 550294 314608 550350
rect 314288 550226 314608 550294
rect 314288 550170 314358 550226
rect 314414 550170 314482 550226
rect 314538 550170 314608 550226
rect 314288 550102 314608 550170
rect 314288 550046 314358 550102
rect 314414 550046 314482 550102
rect 314538 550046 314608 550102
rect 314288 549978 314608 550046
rect 314288 549922 314358 549978
rect 314414 549922 314482 549978
rect 314538 549922 314608 549978
rect 314288 549888 314608 549922
rect 345008 550350 345328 550384
rect 345008 550294 345078 550350
rect 345134 550294 345202 550350
rect 345258 550294 345328 550350
rect 345008 550226 345328 550294
rect 345008 550170 345078 550226
rect 345134 550170 345202 550226
rect 345258 550170 345328 550226
rect 345008 550102 345328 550170
rect 345008 550046 345078 550102
rect 345134 550046 345202 550102
rect 345258 550046 345328 550102
rect 345008 549978 345328 550046
rect 345008 549922 345078 549978
rect 345134 549922 345202 549978
rect 345258 549922 345328 549978
rect 345008 549888 345328 549922
rect 375728 550350 376048 550384
rect 375728 550294 375798 550350
rect 375854 550294 375922 550350
rect 375978 550294 376048 550350
rect 375728 550226 376048 550294
rect 375728 550170 375798 550226
rect 375854 550170 375922 550226
rect 375978 550170 376048 550226
rect 375728 550102 376048 550170
rect 375728 550046 375798 550102
rect 375854 550046 375922 550102
rect 375978 550046 376048 550102
rect 375728 549978 376048 550046
rect 375728 549922 375798 549978
rect 375854 549922 375922 549978
rect 375978 549922 376048 549978
rect 375728 549888 376048 549922
rect 406448 550350 406768 550384
rect 406448 550294 406518 550350
rect 406574 550294 406642 550350
rect 406698 550294 406768 550350
rect 406448 550226 406768 550294
rect 406448 550170 406518 550226
rect 406574 550170 406642 550226
rect 406698 550170 406768 550226
rect 406448 550102 406768 550170
rect 406448 550046 406518 550102
rect 406574 550046 406642 550102
rect 406698 550046 406768 550102
rect 406448 549978 406768 550046
rect 406448 549922 406518 549978
rect 406574 549922 406642 549978
rect 406698 549922 406768 549978
rect 406448 549888 406768 549922
rect 437168 550350 437488 550384
rect 437168 550294 437238 550350
rect 437294 550294 437362 550350
rect 437418 550294 437488 550350
rect 437168 550226 437488 550294
rect 437168 550170 437238 550226
rect 437294 550170 437362 550226
rect 437418 550170 437488 550226
rect 437168 550102 437488 550170
rect 437168 550046 437238 550102
rect 437294 550046 437362 550102
rect 437418 550046 437488 550102
rect 437168 549978 437488 550046
rect 437168 549922 437238 549978
rect 437294 549922 437362 549978
rect 437418 549922 437488 549978
rect 437168 549888 437488 549922
rect 467888 550350 468208 550384
rect 467888 550294 467958 550350
rect 468014 550294 468082 550350
rect 468138 550294 468208 550350
rect 467888 550226 468208 550294
rect 467888 550170 467958 550226
rect 468014 550170 468082 550226
rect 468138 550170 468208 550226
rect 467888 550102 468208 550170
rect 467888 550046 467958 550102
rect 468014 550046 468082 550102
rect 468138 550046 468208 550102
rect 467888 549978 468208 550046
rect 467888 549922 467958 549978
rect 468014 549922 468082 549978
rect 468138 549922 468208 549978
rect 467888 549888 468208 549922
rect 498608 550350 498928 550384
rect 498608 550294 498678 550350
rect 498734 550294 498802 550350
rect 498858 550294 498928 550350
rect 498608 550226 498928 550294
rect 498608 550170 498678 550226
rect 498734 550170 498802 550226
rect 498858 550170 498928 550226
rect 498608 550102 498928 550170
rect 498608 550046 498678 550102
rect 498734 550046 498802 550102
rect 498858 550046 498928 550102
rect 498608 549978 498928 550046
rect 498608 549922 498678 549978
rect 498734 549922 498802 549978
rect 498858 549922 498928 549978
rect 498608 549888 498928 549922
rect 529328 550350 529648 550384
rect 529328 550294 529398 550350
rect 529454 550294 529522 550350
rect 529578 550294 529648 550350
rect 529328 550226 529648 550294
rect 529328 550170 529398 550226
rect 529454 550170 529522 550226
rect 529578 550170 529648 550226
rect 529328 550102 529648 550170
rect 529328 550046 529398 550102
rect 529454 550046 529522 550102
rect 529578 550046 529648 550102
rect 529328 549978 529648 550046
rect 529328 549922 529398 549978
rect 529454 549922 529522 549978
rect 529578 549922 529648 549978
rect 529328 549888 529648 549922
rect 53168 544350 53488 544384
rect 53168 544294 53238 544350
rect 53294 544294 53362 544350
rect 53418 544294 53488 544350
rect 53168 544226 53488 544294
rect 53168 544170 53238 544226
rect 53294 544170 53362 544226
rect 53418 544170 53488 544226
rect 53168 544102 53488 544170
rect 53168 544046 53238 544102
rect 53294 544046 53362 544102
rect 53418 544046 53488 544102
rect 53168 543978 53488 544046
rect 53168 543922 53238 543978
rect 53294 543922 53362 543978
rect 53418 543922 53488 543978
rect 53168 543888 53488 543922
rect 83888 544350 84208 544384
rect 83888 544294 83958 544350
rect 84014 544294 84082 544350
rect 84138 544294 84208 544350
rect 83888 544226 84208 544294
rect 83888 544170 83958 544226
rect 84014 544170 84082 544226
rect 84138 544170 84208 544226
rect 83888 544102 84208 544170
rect 83888 544046 83958 544102
rect 84014 544046 84082 544102
rect 84138 544046 84208 544102
rect 83888 543978 84208 544046
rect 83888 543922 83958 543978
rect 84014 543922 84082 543978
rect 84138 543922 84208 543978
rect 83888 543888 84208 543922
rect 114608 544350 114928 544384
rect 114608 544294 114678 544350
rect 114734 544294 114802 544350
rect 114858 544294 114928 544350
rect 114608 544226 114928 544294
rect 114608 544170 114678 544226
rect 114734 544170 114802 544226
rect 114858 544170 114928 544226
rect 114608 544102 114928 544170
rect 114608 544046 114678 544102
rect 114734 544046 114802 544102
rect 114858 544046 114928 544102
rect 114608 543978 114928 544046
rect 114608 543922 114678 543978
rect 114734 543922 114802 543978
rect 114858 543922 114928 543978
rect 114608 543888 114928 543922
rect 145328 544350 145648 544384
rect 145328 544294 145398 544350
rect 145454 544294 145522 544350
rect 145578 544294 145648 544350
rect 145328 544226 145648 544294
rect 145328 544170 145398 544226
rect 145454 544170 145522 544226
rect 145578 544170 145648 544226
rect 145328 544102 145648 544170
rect 145328 544046 145398 544102
rect 145454 544046 145522 544102
rect 145578 544046 145648 544102
rect 145328 543978 145648 544046
rect 145328 543922 145398 543978
rect 145454 543922 145522 543978
rect 145578 543922 145648 543978
rect 145328 543888 145648 543922
rect 176048 544350 176368 544384
rect 176048 544294 176118 544350
rect 176174 544294 176242 544350
rect 176298 544294 176368 544350
rect 176048 544226 176368 544294
rect 176048 544170 176118 544226
rect 176174 544170 176242 544226
rect 176298 544170 176368 544226
rect 176048 544102 176368 544170
rect 176048 544046 176118 544102
rect 176174 544046 176242 544102
rect 176298 544046 176368 544102
rect 176048 543978 176368 544046
rect 176048 543922 176118 543978
rect 176174 543922 176242 543978
rect 176298 543922 176368 543978
rect 176048 543888 176368 543922
rect 206768 544350 207088 544384
rect 206768 544294 206838 544350
rect 206894 544294 206962 544350
rect 207018 544294 207088 544350
rect 206768 544226 207088 544294
rect 206768 544170 206838 544226
rect 206894 544170 206962 544226
rect 207018 544170 207088 544226
rect 206768 544102 207088 544170
rect 206768 544046 206838 544102
rect 206894 544046 206962 544102
rect 207018 544046 207088 544102
rect 206768 543978 207088 544046
rect 206768 543922 206838 543978
rect 206894 543922 206962 543978
rect 207018 543922 207088 543978
rect 206768 543888 207088 543922
rect 237488 544350 237808 544384
rect 237488 544294 237558 544350
rect 237614 544294 237682 544350
rect 237738 544294 237808 544350
rect 237488 544226 237808 544294
rect 237488 544170 237558 544226
rect 237614 544170 237682 544226
rect 237738 544170 237808 544226
rect 237488 544102 237808 544170
rect 237488 544046 237558 544102
rect 237614 544046 237682 544102
rect 237738 544046 237808 544102
rect 237488 543978 237808 544046
rect 237488 543922 237558 543978
rect 237614 543922 237682 543978
rect 237738 543922 237808 543978
rect 237488 543888 237808 543922
rect 268208 544350 268528 544384
rect 268208 544294 268278 544350
rect 268334 544294 268402 544350
rect 268458 544294 268528 544350
rect 268208 544226 268528 544294
rect 268208 544170 268278 544226
rect 268334 544170 268402 544226
rect 268458 544170 268528 544226
rect 268208 544102 268528 544170
rect 268208 544046 268278 544102
rect 268334 544046 268402 544102
rect 268458 544046 268528 544102
rect 268208 543978 268528 544046
rect 268208 543922 268278 543978
rect 268334 543922 268402 543978
rect 268458 543922 268528 543978
rect 268208 543888 268528 543922
rect 298928 544350 299248 544384
rect 298928 544294 298998 544350
rect 299054 544294 299122 544350
rect 299178 544294 299248 544350
rect 298928 544226 299248 544294
rect 298928 544170 298998 544226
rect 299054 544170 299122 544226
rect 299178 544170 299248 544226
rect 298928 544102 299248 544170
rect 298928 544046 298998 544102
rect 299054 544046 299122 544102
rect 299178 544046 299248 544102
rect 298928 543978 299248 544046
rect 298928 543922 298998 543978
rect 299054 543922 299122 543978
rect 299178 543922 299248 543978
rect 298928 543888 299248 543922
rect 329648 544350 329968 544384
rect 329648 544294 329718 544350
rect 329774 544294 329842 544350
rect 329898 544294 329968 544350
rect 329648 544226 329968 544294
rect 329648 544170 329718 544226
rect 329774 544170 329842 544226
rect 329898 544170 329968 544226
rect 329648 544102 329968 544170
rect 329648 544046 329718 544102
rect 329774 544046 329842 544102
rect 329898 544046 329968 544102
rect 329648 543978 329968 544046
rect 329648 543922 329718 543978
rect 329774 543922 329842 543978
rect 329898 543922 329968 543978
rect 329648 543888 329968 543922
rect 360368 544350 360688 544384
rect 360368 544294 360438 544350
rect 360494 544294 360562 544350
rect 360618 544294 360688 544350
rect 360368 544226 360688 544294
rect 360368 544170 360438 544226
rect 360494 544170 360562 544226
rect 360618 544170 360688 544226
rect 360368 544102 360688 544170
rect 360368 544046 360438 544102
rect 360494 544046 360562 544102
rect 360618 544046 360688 544102
rect 360368 543978 360688 544046
rect 360368 543922 360438 543978
rect 360494 543922 360562 543978
rect 360618 543922 360688 543978
rect 360368 543888 360688 543922
rect 391088 544350 391408 544384
rect 391088 544294 391158 544350
rect 391214 544294 391282 544350
rect 391338 544294 391408 544350
rect 391088 544226 391408 544294
rect 391088 544170 391158 544226
rect 391214 544170 391282 544226
rect 391338 544170 391408 544226
rect 391088 544102 391408 544170
rect 391088 544046 391158 544102
rect 391214 544046 391282 544102
rect 391338 544046 391408 544102
rect 391088 543978 391408 544046
rect 391088 543922 391158 543978
rect 391214 543922 391282 543978
rect 391338 543922 391408 543978
rect 391088 543888 391408 543922
rect 421808 544350 422128 544384
rect 421808 544294 421878 544350
rect 421934 544294 422002 544350
rect 422058 544294 422128 544350
rect 421808 544226 422128 544294
rect 421808 544170 421878 544226
rect 421934 544170 422002 544226
rect 422058 544170 422128 544226
rect 421808 544102 422128 544170
rect 421808 544046 421878 544102
rect 421934 544046 422002 544102
rect 422058 544046 422128 544102
rect 421808 543978 422128 544046
rect 421808 543922 421878 543978
rect 421934 543922 422002 543978
rect 422058 543922 422128 543978
rect 421808 543888 422128 543922
rect 452528 544350 452848 544384
rect 452528 544294 452598 544350
rect 452654 544294 452722 544350
rect 452778 544294 452848 544350
rect 452528 544226 452848 544294
rect 452528 544170 452598 544226
rect 452654 544170 452722 544226
rect 452778 544170 452848 544226
rect 452528 544102 452848 544170
rect 452528 544046 452598 544102
rect 452654 544046 452722 544102
rect 452778 544046 452848 544102
rect 452528 543978 452848 544046
rect 452528 543922 452598 543978
rect 452654 543922 452722 543978
rect 452778 543922 452848 543978
rect 452528 543888 452848 543922
rect 483248 544350 483568 544384
rect 483248 544294 483318 544350
rect 483374 544294 483442 544350
rect 483498 544294 483568 544350
rect 483248 544226 483568 544294
rect 483248 544170 483318 544226
rect 483374 544170 483442 544226
rect 483498 544170 483568 544226
rect 483248 544102 483568 544170
rect 483248 544046 483318 544102
rect 483374 544046 483442 544102
rect 483498 544046 483568 544102
rect 483248 543978 483568 544046
rect 483248 543922 483318 543978
rect 483374 543922 483442 543978
rect 483498 543922 483568 543978
rect 483248 543888 483568 543922
rect 513968 544350 514288 544384
rect 513968 544294 514038 544350
rect 514094 544294 514162 544350
rect 514218 544294 514288 544350
rect 513968 544226 514288 544294
rect 513968 544170 514038 544226
rect 514094 544170 514162 544226
rect 514218 544170 514288 544226
rect 513968 544102 514288 544170
rect 513968 544046 514038 544102
rect 514094 544046 514162 544102
rect 514218 544046 514288 544102
rect 513968 543978 514288 544046
rect 513968 543922 514038 543978
rect 514094 543922 514162 543978
rect 514218 543922 514288 543978
rect 513968 543888 514288 543922
rect 544688 544350 545008 544384
rect 544688 544294 544758 544350
rect 544814 544294 544882 544350
rect 544938 544294 545008 544350
rect 544688 544226 545008 544294
rect 544688 544170 544758 544226
rect 544814 544170 544882 544226
rect 544938 544170 545008 544226
rect 544688 544102 545008 544170
rect 544688 544046 544758 544102
rect 544814 544046 544882 544102
rect 544938 544046 545008 544102
rect 544688 543978 545008 544046
rect 544688 543922 544758 543978
rect 544814 543922 544882 543978
rect 544938 543922 545008 543978
rect 544688 543888 545008 543922
rect 37808 532350 38128 532384
rect 37808 532294 37878 532350
rect 37934 532294 38002 532350
rect 38058 532294 38128 532350
rect 37808 532226 38128 532294
rect 37808 532170 37878 532226
rect 37934 532170 38002 532226
rect 38058 532170 38128 532226
rect 37808 532102 38128 532170
rect 37808 532046 37878 532102
rect 37934 532046 38002 532102
rect 38058 532046 38128 532102
rect 37808 531978 38128 532046
rect 37808 531922 37878 531978
rect 37934 531922 38002 531978
rect 38058 531922 38128 531978
rect 37808 531888 38128 531922
rect 68528 532350 68848 532384
rect 68528 532294 68598 532350
rect 68654 532294 68722 532350
rect 68778 532294 68848 532350
rect 68528 532226 68848 532294
rect 68528 532170 68598 532226
rect 68654 532170 68722 532226
rect 68778 532170 68848 532226
rect 68528 532102 68848 532170
rect 68528 532046 68598 532102
rect 68654 532046 68722 532102
rect 68778 532046 68848 532102
rect 68528 531978 68848 532046
rect 68528 531922 68598 531978
rect 68654 531922 68722 531978
rect 68778 531922 68848 531978
rect 68528 531888 68848 531922
rect 99248 532350 99568 532384
rect 99248 532294 99318 532350
rect 99374 532294 99442 532350
rect 99498 532294 99568 532350
rect 99248 532226 99568 532294
rect 99248 532170 99318 532226
rect 99374 532170 99442 532226
rect 99498 532170 99568 532226
rect 99248 532102 99568 532170
rect 99248 532046 99318 532102
rect 99374 532046 99442 532102
rect 99498 532046 99568 532102
rect 99248 531978 99568 532046
rect 99248 531922 99318 531978
rect 99374 531922 99442 531978
rect 99498 531922 99568 531978
rect 99248 531888 99568 531922
rect 129968 532350 130288 532384
rect 129968 532294 130038 532350
rect 130094 532294 130162 532350
rect 130218 532294 130288 532350
rect 129968 532226 130288 532294
rect 129968 532170 130038 532226
rect 130094 532170 130162 532226
rect 130218 532170 130288 532226
rect 129968 532102 130288 532170
rect 129968 532046 130038 532102
rect 130094 532046 130162 532102
rect 130218 532046 130288 532102
rect 129968 531978 130288 532046
rect 129968 531922 130038 531978
rect 130094 531922 130162 531978
rect 130218 531922 130288 531978
rect 129968 531888 130288 531922
rect 160688 532350 161008 532384
rect 160688 532294 160758 532350
rect 160814 532294 160882 532350
rect 160938 532294 161008 532350
rect 160688 532226 161008 532294
rect 160688 532170 160758 532226
rect 160814 532170 160882 532226
rect 160938 532170 161008 532226
rect 160688 532102 161008 532170
rect 160688 532046 160758 532102
rect 160814 532046 160882 532102
rect 160938 532046 161008 532102
rect 160688 531978 161008 532046
rect 160688 531922 160758 531978
rect 160814 531922 160882 531978
rect 160938 531922 161008 531978
rect 160688 531888 161008 531922
rect 191408 532350 191728 532384
rect 191408 532294 191478 532350
rect 191534 532294 191602 532350
rect 191658 532294 191728 532350
rect 191408 532226 191728 532294
rect 191408 532170 191478 532226
rect 191534 532170 191602 532226
rect 191658 532170 191728 532226
rect 191408 532102 191728 532170
rect 191408 532046 191478 532102
rect 191534 532046 191602 532102
rect 191658 532046 191728 532102
rect 191408 531978 191728 532046
rect 191408 531922 191478 531978
rect 191534 531922 191602 531978
rect 191658 531922 191728 531978
rect 191408 531888 191728 531922
rect 222128 532350 222448 532384
rect 222128 532294 222198 532350
rect 222254 532294 222322 532350
rect 222378 532294 222448 532350
rect 222128 532226 222448 532294
rect 222128 532170 222198 532226
rect 222254 532170 222322 532226
rect 222378 532170 222448 532226
rect 222128 532102 222448 532170
rect 222128 532046 222198 532102
rect 222254 532046 222322 532102
rect 222378 532046 222448 532102
rect 222128 531978 222448 532046
rect 222128 531922 222198 531978
rect 222254 531922 222322 531978
rect 222378 531922 222448 531978
rect 222128 531888 222448 531922
rect 252848 532350 253168 532384
rect 252848 532294 252918 532350
rect 252974 532294 253042 532350
rect 253098 532294 253168 532350
rect 252848 532226 253168 532294
rect 252848 532170 252918 532226
rect 252974 532170 253042 532226
rect 253098 532170 253168 532226
rect 252848 532102 253168 532170
rect 252848 532046 252918 532102
rect 252974 532046 253042 532102
rect 253098 532046 253168 532102
rect 252848 531978 253168 532046
rect 252848 531922 252918 531978
rect 252974 531922 253042 531978
rect 253098 531922 253168 531978
rect 252848 531888 253168 531922
rect 283568 532350 283888 532384
rect 283568 532294 283638 532350
rect 283694 532294 283762 532350
rect 283818 532294 283888 532350
rect 283568 532226 283888 532294
rect 283568 532170 283638 532226
rect 283694 532170 283762 532226
rect 283818 532170 283888 532226
rect 283568 532102 283888 532170
rect 283568 532046 283638 532102
rect 283694 532046 283762 532102
rect 283818 532046 283888 532102
rect 283568 531978 283888 532046
rect 283568 531922 283638 531978
rect 283694 531922 283762 531978
rect 283818 531922 283888 531978
rect 283568 531888 283888 531922
rect 314288 532350 314608 532384
rect 314288 532294 314358 532350
rect 314414 532294 314482 532350
rect 314538 532294 314608 532350
rect 314288 532226 314608 532294
rect 314288 532170 314358 532226
rect 314414 532170 314482 532226
rect 314538 532170 314608 532226
rect 314288 532102 314608 532170
rect 314288 532046 314358 532102
rect 314414 532046 314482 532102
rect 314538 532046 314608 532102
rect 314288 531978 314608 532046
rect 314288 531922 314358 531978
rect 314414 531922 314482 531978
rect 314538 531922 314608 531978
rect 314288 531888 314608 531922
rect 345008 532350 345328 532384
rect 345008 532294 345078 532350
rect 345134 532294 345202 532350
rect 345258 532294 345328 532350
rect 345008 532226 345328 532294
rect 345008 532170 345078 532226
rect 345134 532170 345202 532226
rect 345258 532170 345328 532226
rect 345008 532102 345328 532170
rect 345008 532046 345078 532102
rect 345134 532046 345202 532102
rect 345258 532046 345328 532102
rect 345008 531978 345328 532046
rect 345008 531922 345078 531978
rect 345134 531922 345202 531978
rect 345258 531922 345328 531978
rect 345008 531888 345328 531922
rect 375728 532350 376048 532384
rect 375728 532294 375798 532350
rect 375854 532294 375922 532350
rect 375978 532294 376048 532350
rect 375728 532226 376048 532294
rect 375728 532170 375798 532226
rect 375854 532170 375922 532226
rect 375978 532170 376048 532226
rect 375728 532102 376048 532170
rect 375728 532046 375798 532102
rect 375854 532046 375922 532102
rect 375978 532046 376048 532102
rect 375728 531978 376048 532046
rect 375728 531922 375798 531978
rect 375854 531922 375922 531978
rect 375978 531922 376048 531978
rect 375728 531888 376048 531922
rect 406448 532350 406768 532384
rect 406448 532294 406518 532350
rect 406574 532294 406642 532350
rect 406698 532294 406768 532350
rect 406448 532226 406768 532294
rect 406448 532170 406518 532226
rect 406574 532170 406642 532226
rect 406698 532170 406768 532226
rect 406448 532102 406768 532170
rect 406448 532046 406518 532102
rect 406574 532046 406642 532102
rect 406698 532046 406768 532102
rect 406448 531978 406768 532046
rect 406448 531922 406518 531978
rect 406574 531922 406642 531978
rect 406698 531922 406768 531978
rect 406448 531888 406768 531922
rect 437168 532350 437488 532384
rect 437168 532294 437238 532350
rect 437294 532294 437362 532350
rect 437418 532294 437488 532350
rect 437168 532226 437488 532294
rect 437168 532170 437238 532226
rect 437294 532170 437362 532226
rect 437418 532170 437488 532226
rect 437168 532102 437488 532170
rect 437168 532046 437238 532102
rect 437294 532046 437362 532102
rect 437418 532046 437488 532102
rect 437168 531978 437488 532046
rect 437168 531922 437238 531978
rect 437294 531922 437362 531978
rect 437418 531922 437488 531978
rect 437168 531888 437488 531922
rect 467888 532350 468208 532384
rect 467888 532294 467958 532350
rect 468014 532294 468082 532350
rect 468138 532294 468208 532350
rect 467888 532226 468208 532294
rect 467888 532170 467958 532226
rect 468014 532170 468082 532226
rect 468138 532170 468208 532226
rect 467888 532102 468208 532170
rect 467888 532046 467958 532102
rect 468014 532046 468082 532102
rect 468138 532046 468208 532102
rect 467888 531978 468208 532046
rect 467888 531922 467958 531978
rect 468014 531922 468082 531978
rect 468138 531922 468208 531978
rect 467888 531888 468208 531922
rect 498608 532350 498928 532384
rect 498608 532294 498678 532350
rect 498734 532294 498802 532350
rect 498858 532294 498928 532350
rect 498608 532226 498928 532294
rect 498608 532170 498678 532226
rect 498734 532170 498802 532226
rect 498858 532170 498928 532226
rect 498608 532102 498928 532170
rect 498608 532046 498678 532102
rect 498734 532046 498802 532102
rect 498858 532046 498928 532102
rect 498608 531978 498928 532046
rect 498608 531922 498678 531978
rect 498734 531922 498802 531978
rect 498858 531922 498928 531978
rect 498608 531888 498928 531922
rect 529328 532350 529648 532384
rect 529328 532294 529398 532350
rect 529454 532294 529522 532350
rect 529578 532294 529648 532350
rect 529328 532226 529648 532294
rect 529328 532170 529398 532226
rect 529454 532170 529522 532226
rect 529578 532170 529648 532226
rect 529328 532102 529648 532170
rect 529328 532046 529398 532102
rect 529454 532046 529522 532102
rect 529578 532046 529648 532102
rect 529328 531978 529648 532046
rect 529328 531922 529398 531978
rect 529454 531922 529522 531978
rect 529578 531922 529648 531978
rect 529328 531888 529648 531922
rect 53168 526350 53488 526384
rect 53168 526294 53238 526350
rect 53294 526294 53362 526350
rect 53418 526294 53488 526350
rect 53168 526226 53488 526294
rect 53168 526170 53238 526226
rect 53294 526170 53362 526226
rect 53418 526170 53488 526226
rect 53168 526102 53488 526170
rect 53168 526046 53238 526102
rect 53294 526046 53362 526102
rect 53418 526046 53488 526102
rect 53168 525978 53488 526046
rect 53168 525922 53238 525978
rect 53294 525922 53362 525978
rect 53418 525922 53488 525978
rect 53168 525888 53488 525922
rect 83888 526350 84208 526384
rect 83888 526294 83958 526350
rect 84014 526294 84082 526350
rect 84138 526294 84208 526350
rect 83888 526226 84208 526294
rect 83888 526170 83958 526226
rect 84014 526170 84082 526226
rect 84138 526170 84208 526226
rect 83888 526102 84208 526170
rect 83888 526046 83958 526102
rect 84014 526046 84082 526102
rect 84138 526046 84208 526102
rect 83888 525978 84208 526046
rect 83888 525922 83958 525978
rect 84014 525922 84082 525978
rect 84138 525922 84208 525978
rect 83888 525888 84208 525922
rect 114608 526350 114928 526384
rect 114608 526294 114678 526350
rect 114734 526294 114802 526350
rect 114858 526294 114928 526350
rect 114608 526226 114928 526294
rect 114608 526170 114678 526226
rect 114734 526170 114802 526226
rect 114858 526170 114928 526226
rect 114608 526102 114928 526170
rect 114608 526046 114678 526102
rect 114734 526046 114802 526102
rect 114858 526046 114928 526102
rect 114608 525978 114928 526046
rect 114608 525922 114678 525978
rect 114734 525922 114802 525978
rect 114858 525922 114928 525978
rect 114608 525888 114928 525922
rect 145328 526350 145648 526384
rect 145328 526294 145398 526350
rect 145454 526294 145522 526350
rect 145578 526294 145648 526350
rect 145328 526226 145648 526294
rect 145328 526170 145398 526226
rect 145454 526170 145522 526226
rect 145578 526170 145648 526226
rect 145328 526102 145648 526170
rect 145328 526046 145398 526102
rect 145454 526046 145522 526102
rect 145578 526046 145648 526102
rect 145328 525978 145648 526046
rect 145328 525922 145398 525978
rect 145454 525922 145522 525978
rect 145578 525922 145648 525978
rect 145328 525888 145648 525922
rect 176048 526350 176368 526384
rect 176048 526294 176118 526350
rect 176174 526294 176242 526350
rect 176298 526294 176368 526350
rect 176048 526226 176368 526294
rect 176048 526170 176118 526226
rect 176174 526170 176242 526226
rect 176298 526170 176368 526226
rect 176048 526102 176368 526170
rect 176048 526046 176118 526102
rect 176174 526046 176242 526102
rect 176298 526046 176368 526102
rect 176048 525978 176368 526046
rect 176048 525922 176118 525978
rect 176174 525922 176242 525978
rect 176298 525922 176368 525978
rect 176048 525888 176368 525922
rect 206768 526350 207088 526384
rect 206768 526294 206838 526350
rect 206894 526294 206962 526350
rect 207018 526294 207088 526350
rect 206768 526226 207088 526294
rect 206768 526170 206838 526226
rect 206894 526170 206962 526226
rect 207018 526170 207088 526226
rect 206768 526102 207088 526170
rect 206768 526046 206838 526102
rect 206894 526046 206962 526102
rect 207018 526046 207088 526102
rect 206768 525978 207088 526046
rect 206768 525922 206838 525978
rect 206894 525922 206962 525978
rect 207018 525922 207088 525978
rect 206768 525888 207088 525922
rect 237488 526350 237808 526384
rect 237488 526294 237558 526350
rect 237614 526294 237682 526350
rect 237738 526294 237808 526350
rect 237488 526226 237808 526294
rect 237488 526170 237558 526226
rect 237614 526170 237682 526226
rect 237738 526170 237808 526226
rect 237488 526102 237808 526170
rect 237488 526046 237558 526102
rect 237614 526046 237682 526102
rect 237738 526046 237808 526102
rect 237488 525978 237808 526046
rect 237488 525922 237558 525978
rect 237614 525922 237682 525978
rect 237738 525922 237808 525978
rect 237488 525888 237808 525922
rect 268208 526350 268528 526384
rect 268208 526294 268278 526350
rect 268334 526294 268402 526350
rect 268458 526294 268528 526350
rect 268208 526226 268528 526294
rect 268208 526170 268278 526226
rect 268334 526170 268402 526226
rect 268458 526170 268528 526226
rect 268208 526102 268528 526170
rect 268208 526046 268278 526102
rect 268334 526046 268402 526102
rect 268458 526046 268528 526102
rect 268208 525978 268528 526046
rect 268208 525922 268278 525978
rect 268334 525922 268402 525978
rect 268458 525922 268528 525978
rect 268208 525888 268528 525922
rect 298928 526350 299248 526384
rect 298928 526294 298998 526350
rect 299054 526294 299122 526350
rect 299178 526294 299248 526350
rect 298928 526226 299248 526294
rect 298928 526170 298998 526226
rect 299054 526170 299122 526226
rect 299178 526170 299248 526226
rect 298928 526102 299248 526170
rect 298928 526046 298998 526102
rect 299054 526046 299122 526102
rect 299178 526046 299248 526102
rect 298928 525978 299248 526046
rect 298928 525922 298998 525978
rect 299054 525922 299122 525978
rect 299178 525922 299248 525978
rect 298928 525888 299248 525922
rect 329648 526350 329968 526384
rect 329648 526294 329718 526350
rect 329774 526294 329842 526350
rect 329898 526294 329968 526350
rect 329648 526226 329968 526294
rect 329648 526170 329718 526226
rect 329774 526170 329842 526226
rect 329898 526170 329968 526226
rect 329648 526102 329968 526170
rect 329648 526046 329718 526102
rect 329774 526046 329842 526102
rect 329898 526046 329968 526102
rect 329648 525978 329968 526046
rect 329648 525922 329718 525978
rect 329774 525922 329842 525978
rect 329898 525922 329968 525978
rect 329648 525888 329968 525922
rect 360368 526350 360688 526384
rect 360368 526294 360438 526350
rect 360494 526294 360562 526350
rect 360618 526294 360688 526350
rect 360368 526226 360688 526294
rect 360368 526170 360438 526226
rect 360494 526170 360562 526226
rect 360618 526170 360688 526226
rect 360368 526102 360688 526170
rect 360368 526046 360438 526102
rect 360494 526046 360562 526102
rect 360618 526046 360688 526102
rect 360368 525978 360688 526046
rect 360368 525922 360438 525978
rect 360494 525922 360562 525978
rect 360618 525922 360688 525978
rect 360368 525888 360688 525922
rect 391088 526350 391408 526384
rect 391088 526294 391158 526350
rect 391214 526294 391282 526350
rect 391338 526294 391408 526350
rect 391088 526226 391408 526294
rect 391088 526170 391158 526226
rect 391214 526170 391282 526226
rect 391338 526170 391408 526226
rect 391088 526102 391408 526170
rect 391088 526046 391158 526102
rect 391214 526046 391282 526102
rect 391338 526046 391408 526102
rect 391088 525978 391408 526046
rect 391088 525922 391158 525978
rect 391214 525922 391282 525978
rect 391338 525922 391408 525978
rect 391088 525888 391408 525922
rect 421808 526350 422128 526384
rect 421808 526294 421878 526350
rect 421934 526294 422002 526350
rect 422058 526294 422128 526350
rect 421808 526226 422128 526294
rect 421808 526170 421878 526226
rect 421934 526170 422002 526226
rect 422058 526170 422128 526226
rect 421808 526102 422128 526170
rect 421808 526046 421878 526102
rect 421934 526046 422002 526102
rect 422058 526046 422128 526102
rect 421808 525978 422128 526046
rect 421808 525922 421878 525978
rect 421934 525922 422002 525978
rect 422058 525922 422128 525978
rect 421808 525888 422128 525922
rect 452528 526350 452848 526384
rect 452528 526294 452598 526350
rect 452654 526294 452722 526350
rect 452778 526294 452848 526350
rect 452528 526226 452848 526294
rect 452528 526170 452598 526226
rect 452654 526170 452722 526226
rect 452778 526170 452848 526226
rect 452528 526102 452848 526170
rect 452528 526046 452598 526102
rect 452654 526046 452722 526102
rect 452778 526046 452848 526102
rect 452528 525978 452848 526046
rect 452528 525922 452598 525978
rect 452654 525922 452722 525978
rect 452778 525922 452848 525978
rect 452528 525888 452848 525922
rect 483248 526350 483568 526384
rect 483248 526294 483318 526350
rect 483374 526294 483442 526350
rect 483498 526294 483568 526350
rect 483248 526226 483568 526294
rect 483248 526170 483318 526226
rect 483374 526170 483442 526226
rect 483498 526170 483568 526226
rect 483248 526102 483568 526170
rect 483248 526046 483318 526102
rect 483374 526046 483442 526102
rect 483498 526046 483568 526102
rect 483248 525978 483568 526046
rect 483248 525922 483318 525978
rect 483374 525922 483442 525978
rect 483498 525922 483568 525978
rect 483248 525888 483568 525922
rect 513968 526350 514288 526384
rect 513968 526294 514038 526350
rect 514094 526294 514162 526350
rect 514218 526294 514288 526350
rect 513968 526226 514288 526294
rect 513968 526170 514038 526226
rect 514094 526170 514162 526226
rect 514218 526170 514288 526226
rect 513968 526102 514288 526170
rect 513968 526046 514038 526102
rect 514094 526046 514162 526102
rect 514218 526046 514288 526102
rect 513968 525978 514288 526046
rect 513968 525922 514038 525978
rect 514094 525922 514162 525978
rect 514218 525922 514288 525978
rect 513968 525888 514288 525922
rect 544688 526350 545008 526384
rect 544688 526294 544758 526350
rect 544814 526294 544882 526350
rect 544938 526294 545008 526350
rect 544688 526226 545008 526294
rect 544688 526170 544758 526226
rect 544814 526170 544882 526226
rect 544938 526170 545008 526226
rect 544688 526102 545008 526170
rect 544688 526046 544758 526102
rect 544814 526046 544882 526102
rect 544938 526046 545008 526102
rect 544688 525978 545008 526046
rect 544688 525922 544758 525978
rect 544814 525922 544882 525978
rect 544938 525922 545008 525978
rect 544688 525888 545008 525922
rect 37808 514350 38128 514384
rect 37808 514294 37878 514350
rect 37934 514294 38002 514350
rect 38058 514294 38128 514350
rect 37808 514226 38128 514294
rect 37808 514170 37878 514226
rect 37934 514170 38002 514226
rect 38058 514170 38128 514226
rect 37808 514102 38128 514170
rect 37808 514046 37878 514102
rect 37934 514046 38002 514102
rect 38058 514046 38128 514102
rect 37808 513978 38128 514046
rect 37808 513922 37878 513978
rect 37934 513922 38002 513978
rect 38058 513922 38128 513978
rect 37808 513888 38128 513922
rect 68528 514350 68848 514384
rect 68528 514294 68598 514350
rect 68654 514294 68722 514350
rect 68778 514294 68848 514350
rect 68528 514226 68848 514294
rect 68528 514170 68598 514226
rect 68654 514170 68722 514226
rect 68778 514170 68848 514226
rect 68528 514102 68848 514170
rect 68528 514046 68598 514102
rect 68654 514046 68722 514102
rect 68778 514046 68848 514102
rect 68528 513978 68848 514046
rect 68528 513922 68598 513978
rect 68654 513922 68722 513978
rect 68778 513922 68848 513978
rect 68528 513888 68848 513922
rect 99248 514350 99568 514384
rect 99248 514294 99318 514350
rect 99374 514294 99442 514350
rect 99498 514294 99568 514350
rect 99248 514226 99568 514294
rect 99248 514170 99318 514226
rect 99374 514170 99442 514226
rect 99498 514170 99568 514226
rect 99248 514102 99568 514170
rect 99248 514046 99318 514102
rect 99374 514046 99442 514102
rect 99498 514046 99568 514102
rect 99248 513978 99568 514046
rect 99248 513922 99318 513978
rect 99374 513922 99442 513978
rect 99498 513922 99568 513978
rect 99248 513888 99568 513922
rect 129968 514350 130288 514384
rect 129968 514294 130038 514350
rect 130094 514294 130162 514350
rect 130218 514294 130288 514350
rect 129968 514226 130288 514294
rect 129968 514170 130038 514226
rect 130094 514170 130162 514226
rect 130218 514170 130288 514226
rect 129968 514102 130288 514170
rect 129968 514046 130038 514102
rect 130094 514046 130162 514102
rect 130218 514046 130288 514102
rect 129968 513978 130288 514046
rect 129968 513922 130038 513978
rect 130094 513922 130162 513978
rect 130218 513922 130288 513978
rect 129968 513888 130288 513922
rect 160688 514350 161008 514384
rect 160688 514294 160758 514350
rect 160814 514294 160882 514350
rect 160938 514294 161008 514350
rect 160688 514226 161008 514294
rect 160688 514170 160758 514226
rect 160814 514170 160882 514226
rect 160938 514170 161008 514226
rect 160688 514102 161008 514170
rect 160688 514046 160758 514102
rect 160814 514046 160882 514102
rect 160938 514046 161008 514102
rect 160688 513978 161008 514046
rect 160688 513922 160758 513978
rect 160814 513922 160882 513978
rect 160938 513922 161008 513978
rect 160688 513888 161008 513922
rect 191408 514350 191728 514384
rect 191408 514294 191478 514350
rect 191534 514294 191602 514350
rect 191658 514294 191728 514350
rect 191408 514226 191728 514294
rect 191408 514170 191478 514226
rect 191534 514170 191602 514226
rect 191658 514170 191728 514226
rect 191408 514102 191728 514170
rect 191408 514046 191478 514102
rect 191534 514046 191602 514102
rect 191658 514046 191728 514102
rect 191408 513978 191728 514046
rect 191408 513922 191478 513978
rect 191534 513922 191602 513978
rect 191658 513922 191728 513978
rect 191408 513888 191728 513922
rect 222128 514350 222448 514384
rect 222128 514294 222198 514350
rect 222254 514294 222322 514350
rect 222378 514294 222448 514350
rect 222128 514226 222448 514294
rect 222128 514170 222198 514226
rect 222254 514170 222322 514226
rect 222378 514170 222448 514226
rect 222128 514102 222448 514170
rect 222128 514046 222198 514102
rect 222254 514046 222322 514102
rect 222378 514046 222448 514102
rect 222128 513978 222448 514046
rect 222128 513922 222198 513978
rect 222254 513922 222322 513978
rect 222378 513922 222448 513978
rect 222128 513888 222448 513922
rect 252848 514350 253168 514384
rect 252848 514294 252918 514350
rect 252974 514294 253042 514350
rect 253098 514294 253168 514350
rect 252848 514226 253168 514294
rect 252848 514170 252918 514226
rect 252974 514170 253042 514226
rect 253098 514170 253168 514226
rect 252848 514102 253168 514170
rect 252848 514046 252918 514102
rect 252974 514046 253042 514102
rect 253098 514046 253168 514102
rect 252848 513978 253168 514046
rect 252848 513922 252918 513978
rect 252974 513922 253042 513978
rect 253098 513922 253168 513978
rect 252848 513888 253168 513922
rect 283568 514350 283888 514384
rect 283568 514294 283638 514350
rect 283694 514294 283762 514350
rect 283818 514294 283888 514350
rect 283568 514226 283888 514294
rect 283568 514170 283638 514226
rect 283694 514170 283762 514226
rect 283818 514170 283888 514226
rect 283568 514102 283888 514170
rect 283568 514046 283638 514102
rect 283694 514046 283762 514102
rect 283818 514046 283888 514102
rect 283568 513978 283888 514046
rect 283568 513922 283638 513978
rect 283694 513922 283762 513978
rect 283818 513922 283888 513978
rect 283568 513888 283888 513922
rect 314288 514350 314608 514384
rect 314288 514294 314358 514350
rect 314414 514294 314482 514350
rect 314538 514294 314608 514350
rect 314288 514226 314608 514294
rect 314288 514170 314358 514226
rect 314414 514170 314482 514226
rect 314538 514170 314608 514226
rect 314288 514102 314608 514170
rect 314288 514046 314358 514102
rect 314414 514046 314482 514102
rect 314538 514046 314608 514102
rect 314288 513978 314608 514046
rect 314288 513922 314358 513978
rect 314414 513922 314482 513978
rect 314538 513922 314608 513978
rect 314288 513888 314608 513922
rect 345008 514350 345328 514384
rect 345008 514294 345078 514350
rect 345134 514294 345202 514350
rect 345258 514294 345328 514350
rect 345008 514226 345328 514294
rect 345008 514170 345078 514226
rect 345134 514170 345202 514226
rect 345258 514170 345328 514226
rect 345008 514102 345328 514170
rect 345008 514046 345078 514102
rect 345134 514046 345202 514102
rect 345258 514046 345328 514102
rect 345008 513978 345328 514046
rect 345008 513922 345078 513978
rect 345134 513922 345202 513978
rect 345258 513922 345328 513978
rect 345008 513888 345328 513922
rect 375728 514350 376048 514384
rect 375728 514294 375798 514350
rect 375854 514294 375922 514350
rect 375978 514294 376048 514350
rect 375728 514226 376048 514294
rect 375728 514170 375798 514226
rect 375854 514170 375922 514226
rect 375978 514170 376048 514226
rect 375728 514102 376048 514170
rect 375728 514046 375798 514102
rect 375854 514046 375922 514102
rect 375978 514046 376048 514102
rect 375728 513978 376048 514046
rect 375728 513922 375798 513978
rect 375854 513922 375922 513978
rect 375978 513922 376048 513978
rect 375728 513888 376048 513922
rect 406448 514350 406768 514384
rect 406448 514294 406518 514350
rect 406574 514294 406642 514350
rect 406698 514294 406768 514350
rect 406448 514226 406768 514294
rect 406448 514170 406518 514226
rect 406574 514170 406642 514226
rect 406698 514170 406768 514226
rect 406448 514102 406768 514170
rect 406448 514046 406518 514102
rect 406574 514046 406642 514102
rect 406698 514046 406768 514102
rect 406448 513978 406768 514046
rect 406448 513922 406518 513978
rect 406574 513922 406642 513978
rect 406698 513922 406768 513978
rect 406448 513888 406768 513922
rect 437168 514350 437488 514384
rect 437168 514294 437238 514350
rect 437294 514294 437362 514350
rect 437418 514294 437488 514350
rect 437168 514226 437488 514294
rect 437168 514170 437238 514226
rect 437294 514170 437362 514226
rect 437418 514170 437488 514226
rect 437168 514102 437488 514170
rect 437168 514046 437238 514102
rect 437294 514046 437362 514102
rect 437418 514046 437488 514102
rect 437168 513978 437488 514046
rect 437168 513922 437238 513978
rect 437294 513922 437362 513978
rect 437418 513922 437488 513978
rect 437168 513888 437488 513922
rect 467888 514350 468208 514384
rect 467888 514294 467958 514350
rect 468014 514294 468082 514350
rect 468138 514294 468208 514350
rect 467888 514226 468208 514294
rect 467888 514170 467958 514226
rect 468014 514170 468082 514226
rect 468138 514170 468208 514226
rect 467888 514102 468208 514170
rect 467888 514046 467958 514102
rect 468014 514046 468082 514102
rect 468138 514046 468208 514102
rect 467888 513978 468208 514046
rect 467888 513922 467958 513978
rect 468014 513922 468082 513978
rect 468138 513922 468208 513978
rect 467888 513888 468208 513922
rect 498608 514350 498928 514384
rect 498608 514294 498678 514350
rect 498734 514294 498802 514350
rect 498858 514294 498928 514350
rect 498608 514226 498928 514294
rect 498608 514170 498678 514226
rect 498734 514170 498802 514226
rect 498858 514170 498928 514226
rect 498608 514102 498928 514170
rect 498608 514046 498678 514102
rect 498734 514046 498802 514102
rect 498858 514046 498928 514102
rect 498608 513978 498928 514046
rect 498608 513922 498678 513978
rect 498734 513922 498802 513978
rect 498858 513922 498928 513978
rect 498608 513888 498928 513922
rect 529328 514350 529648 514384
rect 529328 514294 529398 514350
rect 529454 514294 529522 514350
rect 529578 514294 529648 514350
rect 529328 514226 529648 514294
rect 529328 514170 529398 514226
rect 529454 514170 529522 514226
rect 529578 514170 529648 514226
rect 529328 514102 529648 514170
rect 529328 514046 529398 514102
rect 529454 514046 529522 514102
rect 529578 514046 529648 514102
rect 529328 513978 529648 514046
rect 529328 513922 529398 513978
rect 529454 513922 529522 513978
rect 529578 513922 529648 513978
rect 529328 513888 529648 513922
rect 53168 508350 53488 508384
rect 53168 508294 53238 508350
rect 53294 508294 53362 508350
rect 53418 508294 53488 508350
rect 53168 508226 53488 508294
rect 53168 508170 53238 508226
rect 53294 508170 53362 508226
rect 53418 508170 53488 508226
rect 53168 508102 53488 508170
rect 53168 508046 53238 508102
rect 53294 508046 53362 508102
rect 53418 508046 53488 508102
rect 53168 507978 53488 508046
rect 53168 507922 53238 507978
rect 53294 507922 53362 507978
rect 53418 507922 53488 507978
rect 53168 507888 53488 507922
rect 83888 508350 84208 508384
rect 83888 508294 83958 508350
rect 84014 508294 84082 508350
rect 84138 508294 84208 508350
rect 83888 508226 84208 508294
rect 83888 508170 83958 508226
rect 84014 508170 84082 508226
rect 84138 508170 84208 508226
rect 83888 508102 84208 508170
rect 83888 508046 83958 508102
rect 84014 508046 84082 508102
rect 84138 508046 84208 508102
rect 83888 507978 84208 508046
rect 83888 507922 83958 507978
rect 84014 507922 84082 507978
rect 84138 507922 84208 507978
rect 83888 507888 84208 507922
rect 114608 508350 114928 508384
rect 114608 508294 114678 508350
rect 114734 508294 114802 508350
rect 114858 508294 114928 508350
rect 114608 508226 114928 508294
rect 114608 508170 114678 508226
rect 114734 508170 114802 508226
rect 114858 508170 114928 508226
rect 114608 508102 114928 508170
rect 114608 508046 114678 508102
rect 114734 508046 114802 508102
rect 114858 508046 114928 508102
rect 114608 507978 114928 508046
rect 114608 507922 114678 507978
rect 114734 507922 114802 507978
rect 114858 507922 114928 507978
rect 114608 507888 114928 507922
rect 145328 508350 145648 508384
rect 145328 508294 145398 508350
rect 145454 508294 145522 508350
rect 145578 508294 145648 508350
rect 145328 508226 145648 508294
rect 145328 508170 145398 508226
rect 145454 508170 145522 508226
rect 145578 508170 145648 508226
rect 145328 508102 145648 508170
rect 145328 508046 145398 508102
rect 145454 508046 145522 508102
rect 145578 508046 145648 508102
rect 145328 507978 145648 508046
rect 145328 507922 145398 507978
rect 145454 507922 145522 507978
rect 145578 507922 145648 507978
rect 145328 507888 145648 507922
rect 176048 508350 176368 508384
rect 176048 508294 176118 508350
rect 176174 508294 176242 508350
rect 176298 508294 176368 508350
rect 176048 508226 176368 508294
rect 176048 508170 176118 508226
rect 176174 508170 176242 508226
rect 176298 508170 176368 508226
rect 176048 508102 176368 508170
rect 176048 508046 176118 508102
rect 176174 508046 176242 508102
rect 176298 508046 176368 508102
rect 176048 507978 176368 508046
rect 176048 507922 176118 507978
rect 176174 507922 176242 507978
rect 176298 507922 176368 507978
rect 176048 507888 176368 507922
rect 206768 508350 207088 508384
rect 206768 508294 206838 508350
rect 206894 508294 206962 508350
rect 207018 508294 207088 508350
rect 206768 508226 207088 508294
rect 206768 508170 206838 508226
rect 206894 508170 206962 508226
rect 207018 508170 207088 508226
rect 206768 508102 207088 508170
rect 206768 508046 206838 508102
rect 206894 508046 206962 508102
rect 207018 508046 207088 508102
rect 206768 507978 207088 508046
rect 206768 507922 206838 507978
rect 206894 507922 206962 507978
rect 207018 507922 207088 507978
rect 206768 507888 207088 507922
rect 237488 508350 237808 508384
rect 237488 508294 237558 508350
rect 237614 508294 237682 508350
rect 237738 508294 237808 508350
rect 237488 508226 237808 508294
rect 237488 508170 237558 508226
rect 237614 508170 237682 508226
rect 237738 508170 237808 508226
rect 237488 508102 237808 508170
rect 237488 508046 237558 508102
rect 237614 508046 237682 508102
rect 237738 508046 237808 508102
rect 237488 507978 237808 508046
rect 237488 507922 237558 507978
rect 237614 507922 237682 507978
rect 237738 507922 237808 507978
rect 237488 507888 237808 507922
rect 268208 508350 268528 508384
rect 268208 508294 268278 508350
rect 268334 508294 268402 508350
rect 268458 508294 268528 508350
rect 268208 508226 268528 508294
rect 268208 508170 268278 508226
rect 268334 508170 268402 508226
rect 268458 508170 268528 508226
rect 268208 508102 268528 508170
rect 268208 508046 268278 508102
rect 268334 508046 268402 508102
rect 268458 508046 268528 508102
rect 268208 507978 268528 508046
rect 268208 507922 268278 507978
rect 268334 507922 268402 507978
rect 268458 507922 268528 507978
rect 268208 507888 268528 507922
rect 298928 508350 299248 508384
rect 298928 508294 298998 508350
rect 299054 508294 299122 508350
rect 299178 508294 299248 508350
rect 298928 508226 299248 508294
rect 298928 508170 298998 508226
rect 299054 508170 299122 508226
rect 299178 508170 299248 508226
rect 298928 508102 299248 508170
rect 298928 508046 298998 508102
rect 299054 508046 299122 508102
rect 299178 508046 299248 508102
rect 298928 507978 299248 508046
rect 298928 507922 298998 507978
rect 299054 507922 299122 507978
rect 299178 507922 299248 507978
rect 298928 507888 299248 507922
rect 329648 508350 329968 508384
rect 329648 508294 329718 508350
rect 329774 508294 329842 508350
rect 329898 508294 329968 508350
rect 329648 508226 329968 508294
rect 329648 508170 329718 508226
rect 329774 508170 329842 508226
rect 329898 508170 329968 508226
rect 329648 508102 329968 508170
rect 329648 508046 329718 508102
rect 329774 508046 329842 508102
rect 329898 508046 329968 508102
rect 329648 507978 329968 508046
rect 329648 507922 329718 507978
rect 329774 507922 329842 507978
rect 329898 507922 329968 507978
rect 329648 507888 329968 507922
rect 360368 508350 360688 508384
rect 360368 508294 360438 508350
rect 360494 508294 360562 508350
rect 360618 508294 360688 508350
rect 360368 508226 360688 508294
rect 360368 508170 360438 508226
rect 360494 508170 360562 508226
rect 360618 508170 360688 508226
rect 360368 508102 360688 508170
rect 360368 508046 360438 508102
rect 360494 508046 360562 508102
rect 360618 508046 360688 508102
rect 360368 507978 360688 508046
rect 360368 507922 360438 507978
rect 360494 507922 360562 507978
rect 360618 507922 360688 507978
rect 360368 507888 360688 507922
rect 391088 508350 391408 508384
rect 391088 508294 391158 508350
rect 391214 508294 391282 508350
rect 391338 508294 391408 508350
rect 391088 508226 391408 508294
rect 391088 508170 391158 508226
rect 391214 508170 391282 508226
rect 391338 508170 391408 508226
rect 391088 508102 391408 508170
rect 391088 508046 391158 508102
rect 391214 508046 391282 508102
rect 391338 508046 391408 508102
rect 391088 507978 391408 508046
rect 391088 507922 391158 507978
rect 391214 507922 391282 507978
rect 391338 507922 391408 507978
rect 391088 507888 391408 507922
rect 421808 508350 422128 508384
rect 421808 508294 421878 508350
rect 421934 508294 422002 508350
rect 422058 508294 422128 508350
rect 421808 508226 422128 508294
rect 421808 508170 421878 508226
rect 421934 508170 422002 508226
rect 422058 508170 422128 508226
rect 421808 508102 422128 508170
rect 421808 508046 421878 508102
rect 421934 508046 422002 508102
rect 422058 508046 422128 508102
rect 421808 507978 422128 508046
rect 421808 507922 421878 507978
rect 421934 507922 422002 507978
rect 422058 507922 422128 507978
rect 421808 507888 422128 507922
rect 452528 508350 452848 508384
rect 452528 508294 452598 508350
rect 452654 508294 452722 508350
rect 452778 508294 452848 508350
rect 452528 508226 452848 508294
rect 452528 508170 452598 508226
rect 452654 508170 452722 508226
rect 452778 508170 452848 508226
rect 452528 508102 452848 508170
rect 452528 508046 452598 508102
rect 452654 508046 452722 508102
rect 452778 508046 452848 508102
rect 452528 507978 452848 508046
rect 452528 507922 452598 507978
rect 452654 507922 452722 507978
rect 452778 507922 452848 507978
rect 452528 507888 452848 507922
rect 483248 508350 483568 508384
rect 483248 508294 483318 508350
rect 483374 508294 483442 508350
rect 483498 508294 483568 508350
rect 483248 508226 483568 508294
rect 483248 508170 483318 508226
rect 483374 508170 483442 508226
rect 483498 508170 483568 508226
rect 483248 508102 483568 508170
rect 483248 508046 483318 508102
rect 483374 508046 483442 508102
rect 483498 508046 483568 508102
rect 483248 507978 483568 508046
rect 483248 507922 483318 507978
rect 483374 507922 483442 507978
rect 483498 507922 483568 507978
rect 483248 507888 483568 507922
rect 513968 508350 514288 508384
rect 513968 508294 514038 508350
rect 514094 508294 514162 508350
rect 514218 508294 514288 508350
rect 513968 508226 514288 508294
rect 513968 508170 514038 508226
rect 514094 508170 514162 508226
rect 514218 508170 514288 508226
rect 513968 508102 514288 508170
rect 513968 508046 514038 508102
rect 514094 508046 514162 508102
rect 514218 508046 514288 508102
rect 513968 507978 514288 508046
rect 513968 507922 514038 507978
rect 514094 507922 514162 507978
rect 514218 507922 514288 507978
rect 513968 507888 514288 507922
rect 544688 508350 545008 508384
rect 544688 508294 544758 508350
rect 544814 508294 544882 508350
rect 544938 508294 545008 508350
rect 544688 508226 545008 508294
rect 544688 508170 544758 508226
rect 544814 508170 544882 508226
rect 544938 508170 545008 508226
rect 544688 508102 545008 508170
rect 544688 508046 544758 508102
rect 544814 508046 544882 508102
rect 544938 508046 545008 508102
rect 544688 507978 545008 508046
rect 544688 507922 544758 507978
rect 544814 507922 544882 507978
rect 544938 507922 545008 507978
rect 544688 507888 545008 507922
rect 37808 496350 38128 496384
rect 37808 496294 37878 496350
rect 37934 496294 38002 496350
rect 38058 496294 38128 496350
rect 37808 496226 38128 496294
rect 37808 496170 37878 496226
rect 37934 496170 38002 496226
rect 38058 496170 38128 496226
rect 37808 496102 38128 496170
rect 37808 496046 37878 496102
rect 37934 496046 38002 496102
rect 38058 496046 38128 496102
rect 37808 495978 38128 496046
rect 37808 495922 37878 495978
rect 37934 495922 38002 495978
rect 38058 495922 38128 495978
rect 37808 495888 38128 495922
rect 68528 496350 68848 496384
rect 68528 496294 68598 496350
rect 68654 496294 68722 496350
rect 68778 496294 68848 496350
rect 68528 496226 68848 496294
rect 68528 496170 68598 496226
rect 68654 496170 68722 496226
rect 68778 496170 68848 496226
rect 68528 496102 68848 496170
rect 68528 496046 68598 496102
rect 68654 496046 68722 496102
rect 68778 496046 68848 496102
rect 68528 495978 68848 496046
rect 68528 495922 68598 495978
rect 68654 495922 68722 495978
rect 68778 495922 68848 495978
rect 68528 495888 68848 495922
rect 99248 496350 99568 496384
rect 99248 496294 99318 496350
rect 99374 496294 99442 496350
rect 99498 496294 99568 496350
rect 99248 496226 99568 496294
rect 99248 496170 99318 496226
rect 99374 496170 99442 496226
rect 99498 496170 99568 496226
rect 99248 496102 99568 496170
rect 99248 496046 99318 496102
rect 99374 496046 99442 496102
rect 99498 496046 99568 496102
rect 99248 495978 99568 496046
rect 99248 495922 99318 495978
rect 99374 495922 99442 495978
rect 99498 495922 99568 495978
rect 99248 495888 99568 495922
rect 129968 496350 130288 496384
rect 129968 496294 130038 496350
rect 130094 496294 130162 496350
rect 130218 496294 130288 496350
rect 129968 496226 130288 496294
rect 129968 496170 130038 496226
rect 130094 496170 130162 496226
rect 130218 496170 130288 496226
rect 129968 496102 130288 496170
rect 129968 496046 130038 496102
rect 130094 496046 130162 496102
rect 130218 496046 130288 496102
rect 129968 495978 130288 496046
rect 129968 495922 130038 495978
rect 130094 495922 130162 495978
rect 130218 495922 130288 495978
rect 129968 495888 130288 495922
rect 160688 496350 161008 496384
rect 160688 496294 160758 496350
rect 160814 496294 160882 496350
rect 160938 496294 161008 496350
rect 160688 496226 161008 496294
rect 160688 496170 160758 496226
rect 160814 496170 160882 496226
rect 160938 496170 161008 496226
rect 160688 496102 161008 496170
rect 160688 496046 160758 496102
rect 160814 496046 160882 496102
rect 160938 496046 161008 496102
rect 160688 495978 161008 496046
rect 160688 495922 160758 495978
rect 160814 495922 160882 495978
rect 160938 495922 161008 495978
rect 160688 495888 161008 495922
rect 191408 496350 191728 496384
rect 191408 496294 191478 496350
rect 191534 496294 191602 496350
rect 191658 496294 191728 496350
rect 191408 496226 191728 496294
rect 191408 496170 191478 496226
rect 191534 496170 191602 496226
rect 191658 496170 191728 496226
rect 191408 496102 191728 496170
rect 191408 496046 191478 496102
rect 191534 496046 191602 496102
rect 191658 496046 191728 496102
rect 191408 495978 191728 496046
rect 191408 495922 191478 495978
rect 191534 495922 191602 495978
rect 191658 495922 191728 495978
rect 191408 495888 191728 495922
rect 222128 496350 222448 496384
rect 222128 496294 222198 496350
rect 222254 496294 222322 496350
rect 222378 496294 222448 496350
rect 222128 496226 222448 496294
rect 222128 496170 222198 496226
rect 222254 496170 222322 496226
rect 222378 496170 222448 496226
rect 222128 496102 222448 496170
rect 222128 496046 222198 496102
rect 222254 496046 222322 496102
rect 222378 496046 222448 496102
rect 222128 495978 222448 496046
rect 222128 495922 222198 495978
rect 222254 495922 222322 495978
rect 222378 495922 222448 495978
rect 222128 495888 222448 495922
rect 252848 496350 253168 496384
rect 252848 496294 252918 496350
rect 252974 496294 253042 496350
rect 253098 496294 253168 496350
rect 252848 496226 253168 496294
rect 252848 496170 252918 496226
rect 252974 496170 253042 496226
rect 253098 496170 253168 496226
rect 252848 496102 253168 496170
rect 252848 496046 252918 496102
rect 252974 496046 253042 496102
rect 253098 496046 253168 496102
rect 252848 495978 253168 496046
rect 252848 495922 252918 495978
rect 252974 495922 253042 495978
rect 253098 495922 253168 495978
rect 252848 495888 253168 495922
rect 283568 496350 283888 496384
rect 283568 496294 283638 496350
rect 283694 496294 283762 496350
rect 283818 496294 283888 496350
rect 283568 496226 283888 496294
rect 283568 496170 283638 496226
rect 283694 496170 283762 496226
rect 283818 496170 283888 496226
rect 283568 496102 283888 496170
rect 283568 496046 283638 496102
rect 283694 496046 283762 496102
rect 283818 496046 283888 496102
rect 283568 495978 283888 496046
rect 283568 495922 283638 495978
rect 283694 495922 283762 495978
rect 283818 495922 283888 495978
rect 283568 495888 283888 495922
rect 314288 496350 314608 496384
rect 314288 496294 314358 496350
rect 314414 496294 314482 496350
rect 314538 496294 314608 496350
rect 314288 496226 314608 496294
rect 314288 496170 314358 496226
rect 314414 496170 314482 496226
rect 314538 496170 314608 496226
rect 314288 496102 314608 496170
rect 314288 496046 314358 496102
rect 314414 496046 314482 496102
rect 314538 496046 314608 496102
rect 314288 495978 314608 496046
rect 314288 495922 314358 495978
rect 314414 495922 314482 495978
rect 314538 495922 314608 495978
rect 314288 495888 314608 495922
rect 345008 496350 345328 496384
rect 345008 496294 345078 496350
rect 345134 496294 345202 496350
rect 345258 496294 345328 496350
rect 345008 496226 345328 496294
rect 345008 496170 345078 496226
rect 345134 496170 345202 496226
rect 345258 496170 345328 496226
rect 345008 496102 345328 496170
rect 345008 496046 345078 496102
rect 345134 496046 345202 496102
rect 345258 496046 345328 496102
rect 345008 495978 345328 496046
rect 345008 495922 345078 495978
rect 345134 495922 345202 495978
rect 345258 495922 345328 495978
rect 345008 495888 345328 495922
rect 375728 496350 376048 496384
rect 375728 496294 375798 496350
rect 375854 496294 375922 496350
rect 375978 496294 376048 496350
rect 375728 496226 376048 496294
rect 375728 496170 375798 496226
rect 375854 496170 375922 496226
rect 375978 496170 376048 496226
rect 375728 496102 376048 496170
rect 375728 496046 375798 496102
rect 375854 496046 375922 496102
rect 375978 496046 376048 496102
rect 375728 495978 376048 496046
rect 375728 495922 375798 495978
rect 375854 495922 375922 495978
rect 375978 495922 376048 495978
rect 375728 495888 376048 495922
rect 406448 496350 406768 496384
rect 406448 496294 406518 496350
rect 406574 496294 406642 496350
rect 406698 496294 406768 496350
rect 406448 496226 406768 496294
rect 406448 496170 406518 496226
rect 406574 496170 406642 496226
rect 406698 496170 406768 496226
rect 406448 496102 406768 496170
rect 406448 496046 406518 496102
rect 406574 496046 406642 496102
rect 406698 496046 406768 496102
rect 406448 495978 406768 496046
rect 406448 495922 406518 495978
rect 406574 495922 406642 495978
rect 406698 495922 406768 495978
rect 406448 495888 406768 495922
rect 437168 496350 437488 496384
rect 437168 496294 437238 496350
rect 437294 496294 437362 496350
rect 437418 496294 437488 496350
rect 437168 496226 437488 496294
rect 437168 496170 437238 496226
rect 437294 496170 437362 496226
rect 437418 496170 437488 496226
rect 437168 496102 437488 496170
rect 437168 496046 437238 496102
rect 437294 496046 437362 496102
rect 437418 496046 437488 496102
rect 437168 495978 437488 496046
rect 437168 495922 437238 495978
rect 437294 495922 437362 495978
rect 437418 495922 437488 495978
rect 437168 495888 437488 495922
rect 467888 496350 468208 496384
rect 467888 496294 467958 496350
rect 468014 496294 468082 496350
rect 468138 496294 468208 496350
rect 467888 496226 468208 496294
rect 467888 496170 467958 496226
rect 468014 496170 468082 496226
rect 468138 496170 468208 496226
rect 467888 496102 468208 496170
rect 467888 496046 467958 496102
rect 468014 496046 468082 496102
rect 468138 496046 468208 496102
rect 467888 495978 468208 496046
rect 467888 495922 467958 495978
rect 468014 495922 468082 495978
rect 468138 495922 468208 495978
rect 467888 495888 468208 495922
rect 498608 496350 498928 496384
rect 498608 496294 498678 496350
rect 498734 496294 498802 496350
rect 498858 496294 498928 496350
rect 498608 496226 498928 496294
rect 498608 496170 498678 496226
rect 498734 496170 498802 496226
rect 498858 496170 498928 496226
rect 498608 496102 498928 496170
rect 498608 496046 498678 496102
rect 498734 496046 498802 496102
rect 498858 496046 498928 496102
rect 498608 495978 498928 496046
rect 498608 495922 498678 495978
rect 498734 495922 498802 495978
rect 498858 495922 498928 495978
rect 498608 495888 498928 495922
rect 529328 496350 529648 496384
rect 529328 496294 529398 496350
rect 529454 496294 529522 496350
rect 529578 496294 529648 496350
rect 529328 496226 529648 496294
rect 529328 496170 529398 496226
rect 529454 496170 529522 496226
rect 529578 496170 529648 496226
rect 529328 496102 529648 496170
rect 529328 496046 529398 496102
rect 529454 496046 529522 496102
rect 529578 496046 529648 496102
rect 529328 495978 529648 496046
rect 529328 495922 529398 495978
rect 529454 495922 529522 495978
rect 529578 495922 529648 495978
rect 529328 495888 529648 495922
rect 53168 490350 53488 490384
rect 53168 490294 53238 490350
rect 53294 490294 53362 490350
rect 53418 490294 53488 490350
rect 53168 490226 53488 490294
rect 53168 490170 53238 490226
rect 53294 490170 53362 490226
rect 53418 490170 53488 490226
rect 53168 490102 53488 490170
rect 53168 490046 53238 490102
rect 53294 490046 53362 490102
rect 53418 490046 53488 490102
rect 53168 489978 53488 490046
rect 53168 489922 53238 489978
rect 53294 489922 53362 489978
rect 53418 489922 53488 489978
rect 53168 489888 53488 489922
rect 83888 490350 84208 490384
rect 83888 490294 83958 490350
rect 84014 490294 84082 490350
rect 84138 490294 84208 490350
rect 83888 490226 84208 490294
rect 83888 490170 83958 490226
rect 84014 490170 84082 490226
rect 84138 490170 84208 490226
rect 83888 490102 84208 490170
rect 83888 490046 83958 490102
rect 84014 490046 84082 490102
rect 84138 490046 84208 490102
rect 83888 489978 84208 490046
rect 83888 489922 83958 489978
rect 84014 489922 84082 489978
rect 84138 489922 84208 489978
rect 83888 489888 84208 489922
rect 114608 490350 114928 490384
rect 114608 490294 114678 490350
rect 114734 490294 114802 490350
rect 114858 490294 114928 490350
rect 114608 490226 114928 490294
rect 114608 490170 114678 490226
rect 114734 490170 114802 490226
rect 114858 490170 114928 490226
rect 114608 490102 114928 490170
rect 114608 490046 114678 490102
rect 114734 490046 114802 490102
rect 114858 490046 114928 490102
rect 114608 489978 114928 490046
rect 114608 489922 114678 489978
rect 114734 489922 114802 489978
rect 114858 489922 114928 489978
rect 114608 489888 114928 489922
rect 145328 490350 145648 490384
rect 145328 490294 145398 490350
rect 145454 490294 145522 490350
rect 145578 490294 145648 490350
rect 145328 490226 145648 490294
rect 145328 490170 145398 490226
rect 145454 490170 145522 490226
rect 145578 490170 145648 490226
rect 145328 490102 145648 490170
rect 145328 490046 145398 490102
rect 145454 490046 145522 490102
rect 145578 490046 145648 490102
rect 145328 489978 145648 490046
rect 145328 489922 145398 489978
rect 145454 489922 145522 489978
rect 145578 489922 145648 489978
rect 145328 489888 145648 489922
rect 176048 490350 176368 490384
rect 176048 490294 176118 490350
rect 176174 490294 176242 490350
rect 176298 490294 176368 490350
rect 176048 490226 176368 490294
rect 176048 490170 176118 490226
rect 176174 490170 176242 490226
rect 176298 490170 176368 490226
rect 176048 490102 176368 490170
rect 176048 490046 176118 490102
rect 176174 490046 176242 490102
rect 176298 490046 176368 490102
rect 176048 489978 176368 490046
rect 176048 489922 176118 489978
rect 176174 489922 176242 489978
rect 176298 489922 176368 489978
rect 176048 489888 176368 489922
rect 206768 490350 207088 490384
rect 206768 490294 206838 490350
rect 206894 490294 206962 490350
rect 207018 490294 207088 490350
rect 206768 490226 207088 490294
rect 206768 490170 206838 490226
rect 206894 490170 206962 490226
rect 207018 490170 207088 490226
rect 206768 490102 207088 490170
rect 206768 490046 206838 490102
rect 206894 490046 206962 490102
rect 207018 490046 207088 490102
rect 206768 489978 207088 490046
rect 206768 489922 206838 489978
rect 206894 489922 206962 489978
rect 207018 489922 207088 489978
rect 206768 489888 207088 489922
rect 237488 490350 237808 490384
rect 237488 490294 237558 490350
rect 237614 490294 237682 490350
rect 237738 490294 237808 490350
rect 237488 490226 237808 490294
rect 237488 490170 237558 490226
rect 237614 490170 237682 490226
rect 237738 490170 237808 490226
rect 237488 490102 237808 490170
rect 237488 490046 237558 490102
rect 237614 490046 237682 490102
rect 237738 490046 237808 490102
rect 237488 489978 237808 490046
rect 237488 489922 237558 489978
rect 237614 489922 237682 489978
rect 237738 489922 237808 489978
rect 237488 489888 237808 489922
rect 268208 490350 268528 490384
rect 268208 490294 268278 490350
rect 268334 490294 268402 490350
rect 268458 490294 268528 490350
rect 268208 490226 268528 490294
rect 268208 490170 268278 490226
rect 268334 490170 268402 490226
rect 268458 490170 268528 490226
rect 268208 490102 268528 490170
rect 268208 490046 268278 490102
rect 268334 490046 268402 490102
rect 268458 490046 268528 490102
rect 268208 489978 268528 490046
rect 268208 489922 268278 489978
rect 268334 489922 268402 489978
rect 268458 489922 268528 489978
rect 268208 489888 268528 489922
rect 298928 490350 299248 490384
rect 298928 490294 298998 490350
rect 299054 490294 299122 490350
rect 299178 490294 299248 490350
rect 298928 490226 299248 490294
rect 298928 490170 298998 490226
rect 299054 490170 299122 490226
rect 299178 490170 299248 490226
rect 298928 490102 299248 490170
rect 298928 490046 298998 490102
rect 299054 490046 299122 490102
rect 299178 490046 299248 490102
rect 298928 489978 299248 490046
rect 298928 489922 298998 489978
rect 299054 489922 299122 489978
rect 299178 489922 299248 489978
rect 298928 489888 299248 489922
rect 329648 490350 329968 490384
rect 329648 490294 329718 490350
rect 329774 490294 329842 490350
rect 329898 490294 329968 490350
rect 329648 490226 329968 490294
rect 329648 490170 329718 490226
rect 329774 490170 329842 490226
rect 329898 490170 329968 490226
rect 329648 490102 329968 490170
rect 329648 490046 329718 490102
rect 329774 490046 329842 490102
rect 329898 490046 329968 490102
rect 329648 489978 329968 490046
rect 329648 489922 329718 489978
rect 329774 489922 329842 489978
rect 329898 489922 329968 489978
rect 329648 489888 329968 489922
rect 360368 490350 360688 490384
rect 360368 490294 360438 490350
rect 360494 490294 360562 490350
rect 360618 490294 360688 490350
rect 360368 490226 360688 490294
rect 360368 490170 360438 490226
rect 360494 490170 360562 490226
rect 360618 490170 360688 490226
rect 360368 490102 360688 490170
rect 360368 490046 360438 490102
rect 360494 490046 360562 490102
rect 360618 490046 360688 490102
rect 360368 489978 360688 490046
rect 360368 489922 360438 489978
rect 360494 489922 360562 489978
rect 360618 489922 360688 489978
rect 360368 489888 360688 489922
rect 391088 490350 391408 490384
rect 391088 490294 391158 490350
rect 391214 490294 391282 490350
rect 391338 490294 391408 490350
rect 391088 490226 391408 490294
rect 391088 490170 391158 490226
rect 391214 490170 391282 490226
rect 391338 490170 391408 490226
rect 391088 490102 391408 490170
rect 391088 490046 391158 490102
rect 391214 490046 391282 490102
rect 391338 490046 391408 490102
rect 391088 489978 391408 490046
rect 391088 489922 391158 489978
rect 391214 489922 391282 489978
rect 391338 489922 391408 489978
rect 391088 489888 391408 489922
rect 421808 490350 422128 490384
rect 421808 490294 421878 490350
rect 421934 490294 422002 490350
rect 422058 490294 422128 490350
rect 421808 490226 422128 490294
rect 421808 490170 421878 490226
rect 421934 490170 422002 490226
rect 422058 490170 422128 490226
rect 421808 490102 422128 490170
rect 421808 490046 421878 490102
rect 421934 490046 422002 490102
rect 422058 490046 422128 490102
rect 421808 489978 422128 490046
rect 421808 489922 421878 489978
rect 421934 489922 422002 489978
rect 422058 489922 422128 489978
rect 421808 489888 422128 489922
rect 452528 490350 452848 490384
rect 452528 490294 452598 490350
rect 452654 490294 452722 490350
rect 452778 490294 452848 490350
rect 452528 490226 452848 490294
rect 452528 490170 452598 490226
rect 452654 490170 452722 490226
rect 452778 490170 452848 490226
rect 452528 490102 452848 490170
rect 452528 490046 452598 490102
rect 452654 490046 452722 490102
rect 452778 490046 452848 490102
rect 452528 489978 452848 490046
rect 452528 489922 452598 489978
rect 452654 489922 452722 489978
rect 452778 489922 452848 489978
rect 452528 489888 452848 489922
rect 483248 490350 483568 490384
rect 483248 490294 483318 490350
rect 483374 490294 483442 490350
rect 483498 490294 483568 490350
rect 483248 490226 483568 490294
rect 483248 490170 483318 490226
rect 483374 490170 483442 490226
rect 483498 490170 483568 490226
rect 483248 490102 483568 490170
rect 483248 490046 483318 490102
rect 483374 490046 483442 490102
rect 483498 490046 483568 490102
rect 483248 489978 483568 490046
rect 483248 489922 483318 489978
rect 483374 489922 483442 489978
rect 483498 489922 483568 489978
rect 483248 489888 483568 489922
rect 513968 490350 514288 490384
rect 513968 490294 514038 490350
rect 514094 490294 514162 490350
rect 514218 490294 514288 490350
rect 513968 490226 514288 490294
rect 513968 490170 514038 490226
rect 514094 490170 514162 490226
rect 514218 490170 514288 490226
rect 513968 490102 514288 490170
rect 513968 490046 514038 490102
rect 514094 490046 514162 490102
rect 514218 490046 514288 490102
rect 513968 489978 514288 490046
rect 513968 489922 514038 489978
rect 514094 489922 514162 489978
rect 514218 489922 514288 489978
rect 513968 489888 514288 489922
rect 544688 490350 545008 490384
rect 544688 490294 544758 490350
rect 544814 490294 544882 490350
rect 544938 490294 545008 490350
rect 544688 490226 545008 490294
rect 544688 490170 544758 490226
rect 544814 490170 544882 490226
rect 544938 490170 545008 490226
rect 544688 490102 545008 490170
rect 544688 490046 544758 490102
rect 544814 490046 544882 490102
rect 544938 490046 545008 490102
rect 544688 489978 545008 490046
rect 544688 489922 544758 489978
rect 544814 489922 544882 489978
rect 544938 489922 545008 489978
rect 544688 489888 545008 489922
rect 37808 478350 38128 478384
rect 37808 478294 37878 478350
rect 37934 478294 38002 478350
rect 38058 478294 38128 478350
rect 37808 478226 38128 478294
rect 37808 478170 37878 478226
rect 37934 478170 38002 478226
rect 38058 478170 38128 478226
rect 37808 478102 38128 478170
rect 37808 478046 37878 478102
rect 37934 478046 38002 478102
rect 38058 478046 38128 478102
rect 37808 477978 38128 478046
rect 37808 477922 37878 477978
rect 37934 477922 38002 477978
rect 38058 477922 38128 477978
rect 37808 477888 38128 477922
rect 68528 478350 68848 478384
rect 68528 478294 68598 478350
rect 68654 478294 68722 478350
rect 68778 478294 68848 478350
rect 68528 478226 68848 478294
rect 68528 478170 68598 478226
rect 68654 478170 68722 478226
rect 68778 478170 68848 478226
rect 68528 478102 68848 478170
rect 68528 478046 68598 478102
rect 68654 478046 68722 478102
rect 68778 478046 68848 478102
rect 68528 477978 68848 478046
rect 68528 477922 68598 477978
rect 68654 477922 68722 477978
rect 68778 477922 68848 477978
rect 68528 477888 68848 477922
rect 99248 478350 99568 478384
rect 99248 478294 99318 478350
rect 99374 478294 99442 478350
rect 99498 478294 99568 478350
rect 99248 478226 99568 478294
rect 99248 478170 99318 478226
rect 99374 478170 99442 478226
rect 99498 478170 99568 478226
rect 99248 478102 99568 478170
rect 99248 478046 99318 478102
rect 99374 478046 99442 478102
rect 99498 478046 99568 478102
rect 99248 477978 99568 478046
rect 99248 477922 99318 477978
rect 99374 477922 99442 477978
rect 99498 477922 99568 477978
rect 99248 477888 99568 477922
rect 129968 478350 130288 478384
rect 129968 478294 130038 478350
rect 130094 478294 130162 478350
rect 130218 478294 130288 478350
rect 129968 478226 130288 478294
rect 129968 478170 130038 478226
rect 130094 478170 130162 478226
rect 130218 478170 130288 478226
rect 129968 478102 130288 478170
rect 129968 478046 130038 478102
rect 130094 478046 130162 478102
rect 130218 478046 130288 478102
rect 129968 477978 130288 478046
rect 129968 477922 130038 477978
rect 130094 477922 130162 477978
rect 130218 477922 130288 477978
rect 129968 477888 130288 477922
rect 160688 478350 161008 478384
rect 160688 478294 160758 478350
rect 160814 478294 160882 478350
rect 160938 478294 161008 478350
rect 160688 478226 161008 478294
rect 160688 478170 160758 478226
rect 160814 478170 160882 478226
rect 160938 478170 161008 478226
rect 160688 478102 161008 478170
rect 160688 478046 160758 478102
rect 160814 478046 160882 478102
rect 160938 478046 161008 478102
rect 160688 477978 161008 478046
rect 160688 477922 160758 477978
rect 160814 477922 160882 477978
rect 160938 477922 161008 477978
rect 160688 477888 161008 477922
rect 191408 478350 191728 478384
rect 191408 478294 191478 478350
rect 191534 478294 191602 478350
rect 191658 478294 191728 478350
rect 191408 478226 191728 478294
rect 191408 478170 191478 478226
rect 191534 478170 191602 478226
rect 191658 478170 191728 478226
rect 191408 478102 191728 478170
rect 191408 478046 191478 478102
rect 191534 478046 191602 478102
rect 191658 478046 191728 478102
rect 191408 477978 191728 478046
rect 191408 477922 191478 477978
rect 191534 477922 191602 477978
rect 191658 477922 191728 477978
rect 191408 477888 191728 477922
rect 222128 478350 222448 478384
rect 222128 478294 222198 478350
rect 222254 478294 222322 478350
rect 222378 478294 222448 478350
rect 222128 478226 222448 478294
rect 222128 478170 222198 478226
rect 222254 478170 222322 478226
rect 222378 478170 222448 478226
rect 222128 478102 222448 478170
rect 222128 478046 222198 478102
rect 222254 478046 222322 478102
rect 222378 478046 222448 478102
rect 222128 477978 222448 478046
rect 222128 477922 222198 477978
rect 222254 477922 222322 477978
rect 222378 477922 222448 477978
rect 222128 477888 222448 477922
rect 252848 478350 253168 478384
rect 252848 478294 252918 478350
rect 252974 478294 253042 478350
rect 253098 478294 253168 478350
rect 252848 478226 253168 478294
rect 252848 478170 252918 478226
rect 252974 478170 253042 478226
rect 253098 478170 253168 478226
rect 252848 478102 253168 478170
rect 252848 478046 252918 478102
rect 252974 478046 253042 478102
rect 253098 478046 253168 478102
rect 252848 477978 253168 478046
rect 252848 477922 252918 477978
rect 252974 477922 253042 477978
rect 253098 477922 253168 477978
rect 252848 477888 253168 477922
rect 283568 478350 283888 478384
rect 283568 478294 283638 478350
rect 283694 478294 283762 478350
rect 283818 478294 283888 478350
rect 283568 478226 283888 478294
rect 283568 478170 283638 478226
rect 283694 478170 283762 478226
rect 283818 478170 283888 478226
rect 283568 478102 283888 478170
rect 283568 478046 283638 478102
rect 283694 478046 283762 478102
rect 283818 478046 283888 478102
rect 283568 477978 283888 478046
rect 283568 477922 283638 477978
rect 283694 477922 283762 477978
rect 283818 477922 283888 477978
rect 283568 477888 283888 477922
rect 314288 478350 314608 478384
rect 314288 478294 314358 478350
rect 314414 478294 314482 478350
rect 314538 478294 314608 478350
rect 314288 478226 314608 478294
rect 314288 478170 314358 478226
rect 314414 478170 314482 478226
rect 314538 478170 314608 478226
rect 314288 478102 314608 478170
rect 314288 478046 314358 478102
rect 314414 478046 314482 478102
rect 314538 478046 314608 478102
rect 314288 477978 314608 478046
rect 314288 477922 314358 477978
rect 314414 477922 314482 477978
rect 314538 477922 314608 477978
rect 314288 477888 314608 477922
rect 345008 478350 345328 478384
rect 345008 478294 345078 478350
rect 345134 478294 345202 478350
rect 345258 478294 345328 478350
rect 345008 478226 345328 478294
rect 345008 478170 345078 478226
rect 345134 478170 345202 478226
rect 345258 478170 345328 478226
rect 345008 478102 345328 478170
rect 345008 478046 345078 478102
rect 345134 478046 345202 478102
rect 345258 478046 345328 478102
rect 345008 477978 345328 478046
rect 345008 477922 345078 477978
rect 345134 477922 345202 477978
rect 345258 477922 345328 477978
rect 345008 477888 345328 477922
rect 375728 478350 376048 478384
rect 375728 478294 375798 478350
rect 375854 478294 375922 478350
rect 375978 478294 376048 478350
rect 375728 478226 376048 478294
rect 375728 478170 375798 478226
rect 375854 478170 375922 478226
rect 375978 478170 376048 478226
rect 375728 478102 376048 478170
rect 375728 478046 375798 478102
rect 375854 478046 375922 478102
rect 375978 478046 376048 478102
rect 375728 477978 376048 478046
rect 375728 477922 375798 477978
rect 375854 477922 375922 477978
rect 375978 477922 376048 477978
rect 375728 477888 376048 477922
rect 406448 478350 406768 478384
rect 406448 478294 406518 478350
rect 406574 478294 406642 478350
rect 406698 478294 406768 478350
rect 406448 478226 406768 478294
rect 406448 478170 406518 478226
rect 406574 478170 406642 478226
rect 406698 478170 406768 478226
rect 406448 478102 406768 478170
rect 406448 478046 406518 478102
rect 406574 478046 406642 478102
rect 406698 478046 406768 478102
rect 406448 477978 406768 478046
rect 406448 477922 406518 477978
rect 406574 477922 406642 477978
rect 406698 477922 406768 477978
rect 406448 477888 406768 477922
rect 437168 478350 437488 478384
rect 437168 478294 437238 478350
rect 437294 478294 437362 478350
rect 437418 478294 437488 478350
rect 437168 478226 437488 478294
rect 437168 478170 437238 478226
rect 437294 478170 437362 478226
rect 437418 478170 437488 478226
rect 437168 478102 437488 478170
rect 437168 478046 437238 478102
rect 437294 478046 437362 478102
rect 437418 478046 437488 478102
rect 437168 477978 437488 478046
rect 437168 477922 437238 477978
rect 437294 477922 437362 477978
rect 437418 477922 437488 477978
rect 437168 477888 437488 477922
rect 467888 478350 468208 478384
rect 467888 478294 467958 478350
rect 468014 478294 468082 478350
rect 468138 478294 468208 478350
rect 467888 478226 468208 478294
rect 467888 478170 467958 478226
rect 468014 478170 468082 478226
rect 468138 478170 468208 478226
rect 467888 478102 468208 478170
rect 467888 478046 467958 478102
rect 468014 478046 468082 478102
rect 468138 478046 468208 478102
rect 467888 477978 468208 478046
rect 467888 477922 467958 477978
rect 468014 477922 468082 477978
rect 468138 477922 468208 477978
rect 467888 477888 468208 477922
rect 498608 478350 498928 478384
rect 498608 478294 498678 478350
rect 498734 478294 498802 478350
rect 498858 478294 498928 478350
rect 498608 478226 498928 478294
rect 498608 478170 498678 478226
rect 498734 478170 498802 478226
rect 498858 478170 498928 478226
rect 498608 478102 498928 478170
rect 498608 478046 498678 478102
rect 498734 478046 498802 478102
rect 498858 478046 498928 478102
rect 498608 477978 498928 478046
rect 498608 477922 498678 477978
rect 498734 477922 498802 477978
rect 498858 477922 498928 477978
rect 498608 477888 498928 477922
rect 529328 478350 529648 478384
rect 529328 478294 529398 478350
rect 529454 478294 529522 478350
rect 529578 478294 529648 478350
rect 529328 478226 529648 478294
rect 529328 478170 529398 478226
rect 529454 478170 529522 478226
rect 529578 478170 529648 478226
rect 529328 478102 529648 478170
rect 529328 478046 529398 478102
rect 529454 478046 529522 478102
rect 529578 478046 529648 478102
rect 529328 477978 529648 478046
rect 529328 477922 529398 477978
rect 529454 477922 529522 477978
rect 529578 477922 529648 477978
rect 529328 477888 529648 477922
rect 53168 472350 53488 472384
rect 53168 472294 53238 472350
rect 53294 472294 53362 472350
rect 53418 472294 53488 472350
rect 53168 472226 53488 472294
rect 53168 472170 53238 472226
rect 53294 472170 53362 472226
rect 53418 472170 53488 472226
rect 53168 472102 53488 472170
rect 53168 472046 53238 472102
rect 53294 472046 53362 472102
rect 53418 472046 53488 472102
rect 53168 471978 53488 472046
rect 53168 471922 53238 471978
rect 53294 471922 53362 471978
rect 53418 471922 53488 471978
rect 53168 471888 53488 471922
rect 83888 472350 84208 472384
rect 83888 472294 83958 472350
rect 84014 472294 84082 472350
rect 84138 472294 84208 472350
rect 83888 472226 84208 472294
rect 83888 472170 83958 472226
rect 84014 472170 84082 472226
rect 84138 472170 84208 472226
rect 83888 472102 84208 472170
rect 83888 472046 83958 472102
rect 84014 472046 84082 472102
rect 84138 472046 84208 472102
rect 83888 471978 84208 472046
rect 83888 471922 83958 471978
rect 84014 471922 84082 471978
rect 84138 471922 84208 471978
rect 83888 471888 84208 471922
rect 114608 472350 114928 472384
rect 114608 472294 114678 472350
rect 114734 472294 114802 472350
rect 114858 472294 114928 472350
rect 114608 472226 114928 472294
rect 114608 472170 114678 472226
rect 114734 472170 114802 472226
rect 114858 472170 114928 472226
rect 114608 472102 114928 472170
rect 114608 472046 114678 472102
rect 114734 472046 114802 472102
rect 114858 472046 114928 472102
rect 114608 471978 114928 472046
rect 114608 471922 114678 471978
rect 114734 471922 114802 471978
rect 114858 471922 114928 471978
rect 114608 471888 114928 471922
rect 145328 472350 145648 472384
rect 145328 472294 145398 472350
rect 145454 472294 145522 472350
rect 145578 472294 145648 472350
rect 145328 472226 145648 472294
rect 145328 472170 145398 472226
rect 145454 472170 145522 472226
rect 145578 472170 145648 472226
rect 145328 472102 145648 472170
rect 145328 472046 145398 472102
rect 145454 472046 145522 472102
rect 145578 472046 145648 472102
rect 145328 471978 145648 472046
rect 145328 471922 145398 471978
rect 145454 471922 145522 471978
rect 145578 471922 145648 471978
rect 145328 471888 145648 471922
rect 176048 472350 176368 472384
rect 176048 472294 176118 472350
rect 176174 472294 176242 472350
rect 176298 472294 176368 472350
rect 176048 472226 176368 472294
rect 176048 472170 176118 472226
rect 176174 472170 176242 472226
rect 176298 472170 176368 472226
rect 176048 472102 176368 472170
rect 176048 472046 176118 472102
rect 176174 472046 176242 472102
rect 176298 472046 176368 472102
rect 176048 471978 176368 472046
rect 176048 471922 176118 471978
rect 176174 471922 176242 471978
rect 176298 471922 176368 471978
rect 176048 471888 176368 471922
rect 206768 472350 207088 472384
rect 206768 472294 206838 472350
rect 206894 472294 206962 472350
rect 207018 472294 207088 472350
rect 206768 472226 207088 472294
rect 206768 472170 206838 472226
rect 206894 472170 206962 472226
rect 207018 472170 207088 472226
rect 206768 472102 207088 472170
rect 206768 472046 206838 472102
rect 206894 472046 206962 472102
rect 207018 472046 207088 472102
rect 206768 471978 207088 472046
rect 206768 471922 206838 471978
rect 206894 471922 206962 471978
rect 207018 471922 207088 471978
rect 206768 471888 207088 471922
rect 237488 472350 237808 472384
rect 237488 472294 237558 472350
rect 237614 472294 237682 472350
rect 237738 472294 237808 472350
rect 237488 472226 237808 472294
rect 237488 472170 237558 472226
rect 237614 472170 237682 472226
rect 237738 472170 237808 472226
rect 237488 472102 237808 472170
rect 237488 472046 237558 472102
rect 237614 472046 237682 472102
rect 237738 472046 237808 472102
rect 237488 471978 237808 472046
rect 237488 471922 237558 471978
rect 237614 471922 237682 471978
rect 237738 471922 237808 471978
rect 237488 471888 237808 471922
rect 268208 472350 268528 472384
rect 268208 472294 268278 472350
rect 268334 472294 268402 472350
rect 268458 472294 268528 472350
rect 268208 472226 268528 472294
rect 268208 472170 268278 472226
rect 268334 472170 268402 472226
rect 268458 472170 268528 472226
rect 268208 472102 268528 472170
rect 268208 472046 268278 472102
rect 268334 472046 268402 472102
rect 268458 472046 268528 472102
rect 268208 471978 268528 472046
rect 268208 471922 268278 471978
rect 268334 471922 268402 471978
rect 268458 471922 268528 471978
rect 268208 471888 268528 471922
rect 298928 472350 299248 472384
rect 298928 472294 298998 472350
rect 299054 472294 299122 472350
rect 299178 472294 299248 472350
rect 298928 472226 299248 472294
rect 298928 472170 298998 472226
rect 299054 472170 299122 472226
rect 299178 472170 299248 472226
rect 298928 472102 299248 472170
rect 298928 472046 298998 472102
rect 299054 472046 299122 472102
rect 299178 472046 299248 472102
rect 298928 471978 299248 472046
rect 298928 471922 298998 471978
rect 299054 471922 299122 471978
rect 299178 471922 299248 471978
rect 298928 471888 299248 471922
rect 329648 472350 329968 472384
rect 329648 472294 329718 472350
rect 329774 472294 329842 472350
rect 329898 472294 329968 472350
rect 329648 472226 329968 472294
rect 329648 472170 329718 472226
rect 329774 472170 329842 472226
rect 329898 472170 329968 472226
rect 329648 472102 329968 472170
rect 329648 472046 329718 472102
rect 329774 472046 329842 472102
rect 329898 472046 329968 472102
rect 329648 471978 329968 472046
rect 329648 471922 329718 471978
rect 329774 471922 329842 471978
rect 329898 471922 329968 471978
rect 329648 471888 329968 471922
rect 360368 472350 360688 472384
rect 360368 472294 360438 472350
rect 360494 472294 360562 472350
rect 360618 472294 360688 472350
rect 360368 472226 360688 472294
rect 360368 472170 360438 472226
rect 360494 472170 360562 472226
rect 360618 472170 360688 472226
rect 360368 472102 360688 472170
rect 360368 472046 360438 472102
rect 360494 472046 360562 472102
rect 360618 472046 360688 472102
rect 360368 471978 360688 472046
rect 360368 471922 360438 471978
rect 360494 471922 360562 471978
rect 360618 471922 360688 471978
rect 360368 471888 360688 471922
rect 391088 472350 391408 472384
rect 391088 472294 391158 472350
rect 391214 472294 391282 472350
rect 391338 472294 391408 472350
rect 391088 472226 391408 472294
rect 391088 472170 391158 472226
rect 391214 472170 391282 472226
rect 391338 472170 391408 472226
rect 391088 472102 391408 472170
rect 391088 472046 391158 472102
rect 391214 472046 391282 472102
rect 391338 472046 391408 472102
rect 391088 471978 391408 472046
rect 391088 471922 391158 471978
rect 391214 471922 391282 471978
rect 391338 471922 391408 471978
rect 391088 471888 391408 471922
rect 421808 472350 422128 472384
rect 421808 472294 421878 472350
rect 421934 472294 422002 472350
rect 422058 472294 422128 472350
rect 421808 472226 422128 472294
rect 421808 472170 421878 472226
rect 421934 472170 422002 472226
rect 422058 472170 422128 472226
rect 421808 472102 422128 472170
rect 421808 472046 421878 472102
rect 421934 472046 422002 472102
rect 422058 472046 422128 472102
rect 421808 471978 422128 472046
rect 421808 471922 421878 471978
rect 421934 471922 422002 471978
rect 422058 471922 422128 471978
rect 421808 471888 422128 471922
rect 452528 472350 452848 472384
rect 452528 472294 452598 472350
rect 452654 472294 452722 472350
rect 452778 472294 452848 472350
rect 452528 472226 452848 472294
rect 452528 472170 452598 472226
rect 452654 472170 452722 472226
rect 452778 472170 452848 472226
rect 452528 472102 452848 472170
rect 452528 472046 452598 472102
rect 452654 472046 452722 472102
rect 452778 472046 452848 472102
rect 452528 471978 452848 472046
rect 452528 471922 452598 471978
rect 452654 471922 452722 471978
rect 452778 471922 452848 471978
rect 452528 471888 452848 471922
rect 483248 472350 483568 472384
rect 483248 472294 483318 472350
rect 483374 472294 483442 472350
rect 483498 472294 483568 472350
rect 483248 472226 483568 472294
rect 483248 472170 483318 472226
rect 483374 472170 483442 472226
rect 483498 472170 483568 472226
rect 483248 472102 483568 472170
rect 483248 472046 483318 472102
rect 483374 472046 483442 472102
rect 483498 472046 483568 472102
rect 483248 471978 483568 472046
rect 483248 471922 483318 471978
rect 483374 471922 483442 471978
rect 483498 471922 483568 471978
rect 483248 471888 483568 471922
rect 513968 472350 514288 472384
rect 513968 472294 514038 472350
rect 514094 472294 514162 472350
rect 514218 472294 514288 472350
rect 513968 472226 514288 472294
rect 513968 472170 514038 472226
rect 514094 472170 514162 472226
rect 514218 472170 514288 472226
rect 513968 472102 514288 472170
rect 513968 472046 514038 472102
rect 514094 472046 514162 472102
rect 514218 472046 514288 472102
rect 513968 471978 514288 472046
rect 513968 471922 514038 471978
rect 514094 471922 514162 471978
rect 514218 471922 514288 471978
rect 513968 471888 514288 471922
rect 544688 472350 545008 472384
rect 544688 472294 544758 472350
rect 544814 472294 544882 472350
rect 544938 472294 545008 472350
rect 544688 472226 545008 472294
rect 544688 472170 544758 472226
rect 544814 472170 544882 472226
rect 544938 472170 545008 472226
rect 544688 472102 545008 472170
rect 544688 472046 544758 472102
rect 544814 472046 544882 472102
rect 544938 472046 545008 472102
rect 544688 471978 545008 472046
rect 544688 471922 544758 471978
rect 544814 471922 544882 471978
rect 544938 471922 545008 471978
rect 544688 471888 545008 471922
rect 37808 460350 38128 460384
rect 37808 460294 37878 460350
rect 37934 460294 38002 460350
rect 38058 460294 38128 460350
rect 37808 460226 38128 460294
rect 37808 460170 37878 460226
rect 37934 460170 38002 460226
rect 38058 460170 38128 460226
rect 37808 460102 38128 460170
rect 37808 460046 37878 460102
rect 37934 460046 38002 460102
rect 38058 460046 38128 460102
rect 37808 459978 38128 460046
rect 37808 459922 37878 459978
rect 37934 459922 38002 459978
rect 38058 459922 38128 459978
rect 37808 459888 38128 459922
rect 68528 460350 68848 460384
rect 68528 460294 68598 460350
rect 68654 460294 68722 460350
rect 68778 460294 68848 460350
rect 68528 460226 68848 460294
rect 68528 460170 68598 460226
rect 68654 460170 68722 460226
rect 68778 460170 68848 460226
rect 68528 460102 68848 460170
rect 68528 460046 68598 460102
rect 68654 460046 68722 460102
rect 68778 460046 68848 460102
rect 68528 459978 68848 460046
rect 68528 459922 68598 459978
rect 68654 459922 68722 459978
rect 68778 459922 68848 459978
rect 68528 459888 68848 459922
rect 99248 460350 99568 460384
rect 99248 460294 99318 460350
rect 99374 460294 99442 460350
rect 99498 460294 99568 460350
rect 99248 460226 99568 460294
rect 99248 460170 99318 460226
rect 99374 460170 99442 460226
rect 99498 460170 99568 460226
rect 99248 460102 99568 460170
rect 99248 460046 99318 460102
rect 99374 460046 99442 460102
rect 99498 460046 99568 460102
rect 99248 459978 99568 460046
rect 99248 459922 99318 459978
rect 99374 459922 99442 459978
rect 99498 459922 99568 459978
rect 99248 459888 99568 459922
rect 129968 460350 130288 460384
rect 129968 460294 130038 460350
rect 130094 460294 130162 460350
rect 130218 460294 130288 460350
rect 129968 460226 130288 460294
rect 129968 460170 130038 460226
rect 130094 460170 130162 460226
rect 130218 460170 130288 460226
rect 129968 460102 130288 460170
rect 129968 460046 130038 460102
rect 130094 460046 130162 460102
rect 130218 460046 130288 460102
rect 129968 459978 130288 460046
rect 129968 459922 130038 459978
rect 130094 459922 130162 459978
rect 130218 459922 130288 459978
rect 129968 459888 130288 459922
rect 160688 460350 161008 460384
rect 160688 460294 160758 460350
rect 160814 460294 160882 460350
rect 160938 460294 161008 460350
rect 160688 460226 161008 460294
rect 160688 460170 160758 460226
rect 160814 460170 160882 460226
rect 160938 460170 161008 460226
rect 160688 460102 161008 460170
rect 160688 460046 160758 460102
rect 160814 460046 160882 460102
rect 160938 460046 161008 460102
rect 160688 459978 161008 460046
rect 160688 459922 160758 459978
rect 160814 459922 160882 459978
rect 160938 459922 161008 459978
rect 160688 459888 161008 459922
rect 191408 460350 191728 460384
rect 191408 460294 191478 460350
rect 191534 460294 191602 460350
rect 191658 460294 191728 460350
rect 191408 460226 191728 460294
rect 191408 460170 191478 460226
rect 191534 460170 191602 460226
rect 191658 460170 191728 460226
rect 191408 460102 191728 460170
rect 191408 460046 191478 460102
rect 191534 460046 191602 460102
rect 191658 460046 191728 460102
rect 191408 459978 191728 460046
rect 191408 459922 191478 459978
rect 191534 459922 191602 459978
rect 191658 459922 191728 459978
rect 191408 459888 191728 459922
rect 222128 460350 222448 460384
rect 222128 460294 222198 460350
rect 222254 460294 222322 460350
rect 222378 460294 222448 460350
rect 222128 460226 222448 460294
rect 222128 460170 222198 460226
rect 222254 460170 222322 460226
rect 222378 460170 222448 460226
rect 222128 460102 222448 460170
rect 222128 460046 222198 460102
rect 222254 460046 222322 460102
rect 222378 460046 222448 460102
rect 222128 459978 222448 460046
rect 222128 459922 222198 459978
rect 222254 459922 222322 459978
rect 222378 459922 222448 459978
rect 222128 459888 222448 459922
rect 252848 460350 253168 460384
rect 252848 460294 252918 460350
rect 252974 460294 253042 460350
rect 253098 460294 253168 460350
rect 252848 460226 253168 460294
rect 252848 460170 252918 460226
rect 252974 460170 253042 460226
rect 253098 460170 253168 460226
rect 252848 460102 253168 460170
rect 252848 460046 252918 460102
rect 252974 460046 253042 460102
rect 253098 460046 253168 460102
rect 252848 459978 253168 460046
rect 252848 459922 252918 459978
rect 252974 459922 253042 459978
rect 253098 459922 253168 459978
rect 252848 459888 253168 459922
rect 283568 460350 283888 460384
rect 283568 460294 283638 460350
rect 283694 460294 283762 460350
rect 283818 460294 283888 460350
rect 283568 460226 283888 460294
rect 283568 460170 283638 460226
rect 283694 460170 283762 460226
rect 283818 460170 283888 460226
rect 283568 460102 283888 460170
rect 283568 460046 283638 460102
rect 283694 460046 283762 460102
rect 283818 460046 283888 460102
rect 283568 459978 283888 460046
rect 283568 459922 283638 459978
rect 283694 459922 283762 459978
rect 283818 459922 283888 459978
rect 283568 459888 283888 459922
rect 314288 460350 314608 460384
rect 314288 460294 314358 460350
rect 314414 460294 314482 460350
rect 314538 460294 314608 460350
rect 314288 460226 314608 460294
rect 314288 460170 314358 460226
rect 314414 460170 314482 460226
rect 314538 460170 314608 460226
rect 314288 460102 314608 460170
rect 314288 460046 314358 460102
rect 314414 460046 314482 460102
rect 314538 460046 314608 460102
rect 314288 459978 314608 460046
rect 314288 459922 314358 459978
rect 314414 459922 314482 459978
rect 314538 459922 314608 459978
rect 314288 459888 314608 459922
rect 345008 460350 345328 460384
rect 345008 460294 345078 460350
rect 345134 460294 345202 460350
rect 345258 460294 345328 460350
rect 345008 460226 345328 460294
rect 345008 460170 345078 460226
rect 345134 460170 345202 460226
rect 345258 460170 345328 460226
rect 345008 460102 345328 460170
rect 345008 460046 345078 460102
rect 345134 460046 345202 460102
rect 345258 460046 345328 460102
rect 345008 459978 345328 460046
rect 345008 459922 345078 459978
rect 345134 459922 345202 459978
rect 345258 459922 345328 459978
rect 345008 459888 345328 459922
rect 375728 460350 376048 460384
rect 375728 460294 375798 460350
rect 375854 460294 375922 460350
rect 375978 460294 376048 460350
rect 375728 460226 376048 460294
rect 375728 460170 375798 460226
rect 375854 460170 375922 460226
rect 375978 460170 376048 460226
rect 375728 460102 376048 460170
rect 375728 460046 375798 460102
rect 375854 460046 375922 460102
rect 375978 460046 376048 460102
rect 375728 459978 376048 460046
rect 375728 459922 375798 459978
rect 375854 459922 375922 459978
rect 375978 459922 376048 459978
rect 375728 459888 376048 459922
rect 406448 460350 406768 460384
rect 406448 460294 406518 460350
rect 406574 460294 406642 460350
rect 406698 460294 406768 460350
rect 406448 460226 406768 460294
rect 406448 460170 406518 460226
rect 406574 460170 406642 460226
rect 406698 460170 406768 460226
rect 406448 460102 406768 460170
rect 406448 460046 406518 460102
rect 406574 460046 406642 460102
rect 406698 460046 406768 460102
rect 406448 459978 406768 460046
rect 406448 459922 406518 459978
rect 406574 459922 406642 459978
rect 406698 459922 406768 459978
rect 406448 459888 406768 459922
rect 437168 460350 437488 460384
rect 437168 460294 437238 460350
rect 437294 460294 437362 460350
rect 437418 460294 437488 460350
rect 437168 460226 437488 460294
rect 437168 460170 437238 460226
rect 437294 460170 437362 460226
rect 437418 460170 437488 460226
rect 437168 460102 437488 460170
rect 437168 460046 437238 460102
rect 437294 460046 437362 460102
rect 437418 460046 437488 460102
rect 437168 459978 437488 460046
rect 437168 459922 437238 459978
rect 437294 459922 437362 459978
rect 437418 459922 437488 459978
rect 437168 459888 437488 459922
rect 467888 460350 468208 460384
rect 467888 460294 467958 460350
rect 468014 460294 468082 460350
rect 468138 460294 468208 460350
rect 467888 460226 468208 460294
rect 467888 460170 467958 460226
rect 468014 460170 468082 460226
rect 468138 460170 468208 460226
rect 467888 460102 468208 460170
rect 467888 460046 467958 460102
rect 468014 460046 468082 460102
rect 468138 460046 468208 460102
rect 467888 459978 468208 460046
rect 467888 459922 467958 459978
rect 468014 459922 468082 459978
rect 468138 459922 468208 459978
rect 467888 459888 468208 459922
rect 498608 460350 498928 460384
rect 498608 460294 498678 460350
rect 498734 460294 498802 460350
rect 498858 460294 498928 460350
rect 498608 460226 498928 460294
rect 498608 460170 498678 460226
rect 498734 460170 498802 460226
rect 498858 460170 498928 460226
rect 498608 460102 498928 460170
rect 498608 460046 498678 460102
rect 498734 460046 498802 460102
rect 498858 460046 498928 460102
rect 498608 459978 498928 460046
rect 498608 459922 498678 459978
rect 498734 459922 498802 459978
rect 498858 459922 498928 459978
rect 498608 459888 498928 459922
rect 529328 460350 529648 460384
rect 529328 460294 529398 460350
rect 529454 460294 529522 460350
rect 529578 460294 529648 460350
rect 529328 460226 529648 460294
rect 529328 460170 529398 460226
rect 529454 460170 529522 460226
rect 529578 460170 529648 460226
rect 529328 460102 529648 460170
rect 529328 460046 529398 460102
rect 529454 460046 529522 460102
rect 529578 460046 529648 460102
rect 529328 459978 529648 460046
rect 529328 459922 529398 459978
rect 529454 459922 529522 459978
rect 529578 459922 529648 459978
rect 529328 459888 529648 459922
rect 53168 454350 53488 454384
rect 53168 454294 53238 454350
rect 53294 454294 53362 454350
rect 53418 454294 53488 454350
rect 53168 454226 53488 454294
rect 53168 454170 53238 454226
rect 53294 454170 53362 454226
rect 53418 454170 53488 454226
rect 53168 454102 53488 454170
rect 53168 454046 53238 454102
rect 53294 454046 53362 454102
rect 53418 454046 53488 454102
rect 53168 453978 53488 454046
rect 53168 453922 53238 453978
rect 53294 453922 53362 453978
rect 53418 453922 53488 453978
rect 53168 453888 53488 453922
rect 83888 454350 84208 454384
rect 83888 454294 83958 454350
rect 84014 454294 84082 454350
rect 84138 454294 84208 454350
rect 83888 454226 84208 454294
rect 83888 454170 83958 454226
rect 84014 454170 84082 454226
rect 84138 454170 84208 454226
rect 83888 454102 84208 454170
rect 83888 454046 83958 454102
rect 84014 454046 84082 454102
rect 84138 454046 84208 454102
rect 83888 453978 84208 454046
rect 83888 453922 83958 453978
rect 84014 453922 84082 453978
rect 84138 453922 84208 453978
rect 83888 453888 84208 453922
rect 114608 454350 114928 454384
rect 114608 454294 114678 454350
rect 114734 454294 114802 454350
rect 114858 454294 114928 454350
rect 114608 454226 114928 454294
rect 114608 454170 114678 454226
rect 114734 454170 114802 454226
rect 114858 454170 114928 454226
rect 114608 454102 114928 454170
rect 114608 454046 114678 454102
rect 114734 454046 114802 454102
rect 114858 454046 114928 454102
rect 114608 453978 114928 454046
rect 114608 453922 114678 453978
rect 114734 453922 114802 453978
rect 114858 453922 114928 453978
rect 114608 453888 114928 453922
rect 145328 454350 145648 454384
rect 145328 454294 145398 454350
rect 145454 454294 145522 454350
rect 145578 454294 145648 454350
rect 145328 454226 145648 454294
rect 145328 454170 145398 454226
rect 145454 454170 145522 454226
rect 145578 454170 145648 454226
rect 145328 454102 145648 454170
rect 145328 454046 145398 454102
rect 145454 454046 145522 454102
rect 145578 454046 145648 454102
rect 145328 453978 145648 454046
rect 145328 453922 145398 453978
rect 145454 453922 145522 453978
rect 145578 453922 145648 453978
rect 145328 453888 145648 453922
rect 176048 454350 176368 454384
rect 176048 454294 176118 454350
rect 176174 454294 176242 454350
rect 176298 454294 176368 454350
rect 176048 454226 176368 454294
rect 176048 454170 176118 454226
rect 176174 454170 176242 454226
rect 176298 454170 176368 454226
rect 176048 454102 176368 454170
rect 176048 454046 176118 454102
rect 176174 454046 176242 454102
rect 176298 454046 176368 454102
rect 176048 453978 176368 454046
rect 176048 453922 176118 453978
rect 176174 453922 176242 453978
rect 176298 453922 176368 453978
rect 176048 453888 176368 453922
rect 206768 454350 207088 454384
rect 206768 454294 206838 454350
rect 206894 454294 206962 454350
rect 207018 454294 207088 454350
rect 206768 454226 207088 454294
rect 206768 454170 206838 454226
rect 206894 454170 206962 454226
rect 207018 454170 207088 454226
rect 206768 454102 207088 454170
rect 206768 454046 206838 454102
rect 206894 454046 206962 454102
rect 207018 454046 207088 454102
rect 206768 453978 207088 454046
rect 206768 453922 206838 453978
rect 206894 453922 206962 453978
rect 207018 453922 207088 453978
rect 206768 453888 207088 453922
rect 237488 454350 237808 454384
rect 237488 454294 237558 454350
rect 237614 454294 237682 454350
rect 237738 454294 237808 454350
rect 237488 454226 237808 454294
rect 237488 454170 237558 454226
rect 237614 454170 237682 454226
rect 237738 454170 237808 454226
rect 237488 454102 237808 454170
rect 237488 454046 237558 454102
rect 237614 454046 237682 454102
rect 237738 454046 237808 454102
rect 237488 453978 237808 454046
rect 237488 453922 237558 453978
rect 237614 453922 237682 453978
rect 237738 453922 237808 453978
rect 237488 453888 237808 453922
rect 268208 454350 268528 454384
rect 268208 454294 268278 454350
rect 268334 454294 268402 454350
rect 268458 454294 268528 454350
rect 268208 454226 268528 454294
rect 268208 454170 268278 454226
rect 268334 454170 268402 454226
rect 268458 454170 268528 454226
rect 268208 454102 268528 454170
rect 268208 454046 268278 454102
rect 268334 454046 268402 454102
rect 268458 454046 268528 454102
rect 268208 453978 268528 454046
rect 268208 453922 268278 453978
rect 268334 453922 268402 453978
rect 268458 453922 268528 453978
rect 268208 453888 268528 453922
rect 298928 454350 299248 454384
rect 298928 454294 298998 454350
rect 299054 454294 299122 454350
rect 299178 454294 299248 454350
rect 298928 454226 299248 454294
rect 298928 454170 298998 454226
rect 299054 454170 299122 454226
rect 299178 454170 299248 454226
rect 298928 454102 299248 454170
rect 298928 454046 298998 454102
rect 299054 454046 299122 454102
rect 299178 454046 299248 454102
rect 298928 453978 299248 454046
rect 298928 453922 298998 453978
rect 299054 453922 299122 453978
rect 299178 453922 299248 453978
rect 298928 453888 299248 453922
rect 329648 454350 329968 454384
rect 329648 454294 329718 454350
rect 329774 454294 329842 454350
rect 329898 454294 329968 454350
rect 329648 454226 329968 454294
rect 329648 454170 329718 454226
rect 329774 454170 329842 454226
rect 329898 454170 329968 454226
rect 329648 454102 329968 454170
rect 329648 454046 329718 454102
rect 329774 454046 329842 454102
rect 329898 454046 329968 454102
rect 329648 453978 329968 454046
rect 329648 453922 329718 453978
rect 329774 453922 329842 453978
rect 329898 453922 329968 453978
rect 329648 453888 329968 453922
rect 360368 454350 360688 454384
rect 360368 454294 360438 454350
rect 360494 454294 360562 454350
rect 360618 454294 360688 454350
rect 360368 454226 360688 454294
rect 360368 454170 360438 454226
rect 360494 454170 360562 454226
rect 360618 454170 360688 454226
rect 360368 454102 360688 454170
rect 360368 454046 360438 454102
rect 360494 454046 360562 454102
rect 360618 454046 360688 454102
rect 360368 453978 360688 454046
rect 360368 453922 360438 453978
rect 360494 453922 360562 453978
rect 360618 453922 360688 453978
rect 360368 453888 360688 453922
rect 391088 454350 391408 454384
rect 391088 454294 391158 454350
rect 391214 454294 391282 454350
rect 391338 454294 391408 454350
rect 391088 454226 391408 454294
rect 391088 454170 391158 454226
rect 391214 454170 391282 454226
rect 391338 454170 391408 454226
rect 391088 454102 391408 454170
rect 391088 454046 391158 454102
rect 391214 454046 391282 454102
rect 391338 454046 391408 454102
rect 391088 453978 391408 454046
rect 391088 453922 391158 453978
rect 391214 453922 391282 453978
rect 391338 453922 391408 453978
rect 391088 453888 391408 453922
rect 421808 454350 422128 454384
rect 421808 454294 421878 454350
rect 421934 454294 422002 454350
rect 422058 454294 422128 454350
rect 421808 454226 422128 454294
rect 421808 454170 421878 454226
rect 421934 454170 422002 454226
rect 422058 454170 422128 454226
rect 421808 454102 422128 454170
rect 421808 454046 421878 454102
rect 421934 454046 422002 454102
rect 422058 454046 422128 454102
rect 421808 453978 422128 454046
rect 421808 453922 421878 453978
rect 421934 453922 422002 453978
rect 422058 453922 422128 453978
rect 421808 453888 422128 453922
rect 452528 454350 452848 454384
rect 452528 454294 452598 454350
rect 452654 454294 452722 454350
rect 452778 454294 452848 454350
rect 452528 454226 452848 454294
rect 452528 454170 452598 454226
rect 452654 454170 452722 454226
rect 452778 454170 452848 454226
rect 452528 454102 452848 454170
rect 452528 454046 452598 454102
rect 452654 454046 452722 454102
rect 452778 454046 452848 454102
rect 452528 453978 452848 454046
rect 452528 453922 452598 453978
rect 452654 453922 452722 453978
rect 452778 453922 452848 453978
rect 452528 453888 452848 453922
rect 483248 454350 483568 454384
rect 483248 454294 483318 454350
rect 483374 454294 483442 454350
rect 483498 454294 483568 454350
rect 483248 454226 483568 454294
rect 483248 454170 483318 454226
rect 483374 454170 483442 454226
rect 483498 454170 483568 454226
rect 483248 454102 483568 454170
rect 483248 454046 483318 454102
rect 483374 454046 483442 454102
rect 483498 454046 483568 454102
rect 483248 453978 483568 454046
rect 483248 453922 483318 453978
rect 483374 453922 483442 453978
rect 483498 453922 483568 453978
rect 483248 453888 483568 453922
rect 513968 454350 514288 454384
rect 513968 454294 514038 454350
rect 514094 454294 514162 454350
rect 514218 454294 514288 454350
rect 513968 454226 514288 454294
rect 513968 454170 514038 454226
rect 514094 454170 514162 454226
rect 514218 454170 514288 454226
rect 513968 454102 514288 454170
rect 513968 454046 514038 454102
rect 514094 454046 514162 454102
rect 514218 454046 514288 454102
rect 513968 453978 514288 454046
rect 513968 453922 514038 453978
rect 514094 453922 514162 453978
rect 514218 453922 514288 453978
rect 513968 453888 514288 453922
rect 544688 454350 545008 454384
rect 544688 454294 544758 454350
rect 544814 454294 544882 454350
rect 544938 454294 545008 454350
rect 544688 454226 545008 454294
rect 544688 454170 544758 454226
rect 544814 454170 544882 454226
rect 544938 454170 545008 454226
rect 544688 454102 545008 454170
rect 544688 454046 544758 454102
rect 544814 454046 544882 454102
rect 544938 454046 545008 454102
rect 544688 453978 545008 454046
rect 544688 453922 544758 453978
rect 544814 453922 544882 453978
rect 544938 453922 545008 453978
rect 544688 453888 545008 453922
rect 37808 442350 38128 442384
rect 37808 442294 37878 442350
rect 37934 442294 38002 442350
rect 38058 442294 38128 442350
rect 37808 442226 38128 442294
rect 37808 442170 37878 442226
rect 37934 442170 38002 442226
rect 38058 442170 38128 442226
rect 37808 442102 38128 442170
rect 37808 442046 37878 442102
rect 37934 442046 38002 442102
rect 38058 442046 38128 442102
rect 37808 441978 38128 442046
rect 37808 441922 37878 441978
rect 37934 441922 38002 441978
rect 38058 441922 38128 441978
rect 37808 441888 38128 441922
rect 68528 442350 68848 442384
rect 68528 442294 68598 442350
rect 68654 442294 68722 442350
rect 68778 442294 68848 442350
rect 68528 442226 68848 442294
rect 68528 442170 68598 442226
rect 68654 442170 68722 442226
rect 68778 442170 68848 442226
rect 68528 442102 68848 442170
rect 68528 442046 68598 442102
rect 68654 442046 68722 442102
rect 68778 442046 68848 442102
rect 68528 441978 68848 442046
rect 68528 441922 68598 441978
rect 68654 441922 68722 441978
rect 68778 441922 68848 441978
rect 68528 441888 68848 441922
rect 99248 442350 99568 442384
rect 99248 442294 99318 442350
rect 99374 442294 99442 442350
rect 99498 442294 99568 442350
rect 99248 442226 99568 442294
rect 99248 442170 99318 442226
rect 99374 442170 99442 442226
rect 99498 442170 99568 442226
rect 99248 442102 99568 442170
rect 99248 442046 99318 442102
rect 99374 442046 99442 442102
rect 99498 442046 99568 442102
rect 99248 441978 99568 442046
rect 99248 441922 99318 441978
rect 99374 441922 99442 441978
rect 99498 441922 99568 441978
rect 99248 441888 99568 441922
rect 129968 442350 130288 442384
rect 129968 442294 130038 442350
rect 130094 442294 130162 442350
rect 130218 442294 130288 442350
rect 129968 442226 130288 442294
rect 129968 442170 130038 442226
rect 130094 442170 130162 442226
rect 130218 442170 130288 442226
rect 129968 442102 130288 442170
rect 129968 442046 130038 442102
rect 130094 442046 130162 442102
rect 130218 442046 130288 442102
rect 129968 441978 130288 442046
rect 129968 441922 130038 441978
rect 130094 441922 130162 441978
rect 130218 441922 130288 441978
rect 129968 441888 130288 441922
rect 160688 442350 161008 442384
rect 160688 442294 160758 442350
rect 160814 442294 160882 442350
rect 160938 442294 161008 442350
rect 160688 442226 161008 442294
rect 160688 442170 160758 442226
rect 160814 442170 160882 442226
rect 160938 442170 161008 442226
rect 160688 442102 161008 442170
rect 160688 442046 160758 442102
rect 160814 442046 160882 442102
rect 160938 442046 161008 442102
rect 160688 441978 161008 442046
rect 160688 441922 160758 441978
rect 160814 441922 160882 441978
rect 160938 441922 161008 441978
rect 160688 441888 161008 441922
rect 191408 442350 191728 442384
rect 191408 442294 191478 442350
rect 191534 442294 191602 442350
rect 191658 442294 191728 442350
rect 191408 442226 191728 442294
rect 191408 442170 191478 442226
rect 191534 442170 191602 442226
rect 191658 442170 191728 442226
rect 191408 442102 191728 442170
rect 191408 442046 191478 442102
rect 191534 442046 191602 442102
rect 191658 442046 191728 442102
rect 191408 441978 191728 442046
rect 191408 441922 191478 441978
rect 191534 441922 191602 441978
rect 191658 441922 191728 441978
rect 191408 441888 191728 441922
rect 222128 442350 222448 442384
rect 222128 442294 222198 442350
rect 222254 442294 222322 442350
rect 222378 442294 222448 442350
rect 222128 442226 222448 442294
rect 222128 442170 222198 442226
rect 222254 442170 222322 442226
rect 222378 442170 222448 442226
rect 222128 442102 222448 442170
rect 222128 442046 222198 442102
rect 222254 442046 222322 442102
rect 222378 442046 222448 442102
rect 222128 441978 222448 442046
rect 222128 441922 222198 441978
rect 222254 441922 222322 441978
rect 222378 441922 222448 441978
rect 222128 441888 222448 441922
rect 252848 442350 253168 442384
rect 252848 442294 252918 442350
rect 252974 442294 253042 442350
rect 253098 442294 253168 442350
rect 252848 442226 253168 442294
rect 252848 442170 252918 442226
rect 252974 442170 253042 442226
rect 253098 442170 253168 442226
rect 252848 442102 253168 442170
rect 252848 442046 252918 442102
rect 252974 442046 253042 442102
rect 253098 442046 253168 442102
rect 252848 441978 253168 442046
rect 252848 441922 252918 441978
rect 252974 441922 253042 441978
rect 253098 441922 253168 441978
rect 252848 441888 253168 441922
rect 283568 442350 283888 442384
rect 283568 442294 283638 442350
rect 283694 442294 283762 442350
rect 283818 442294 283888 442350
rect 283568 442226 283888 442294
rect 283568 442170 283638 442226
rect 283694 442170 283762 442226
rect 283818 442170 283888 442226
rect 283568 442102 283888 442170
rect 283568 442046 283638 442102
rect 283694 442046 283762 442102
rect 283818 442046 283888 442102
rect 283568 441978 283888 442046
rect 283568 441922 283638 441978
rect 283694 441922 283762 441978
rect 283818 441922 283888 441978
rect 283568 441888 283888 441922
rect 314288 442350 314608 442384
rect 314288 442294 314358 442350
rect 314414 442294 314482 442350
rect 314538 442294 314608 442350
rect 314288 442226 314608 442294
rect 314288 442170 314358 442226
rect 314414 442170 314482 442226
rect 314538 442170 314608 442226
rect 314288 442102 314608 442170
rect 314288 442046 314358 442102
rect 314414 442046 314482 442102
rect 314538 442046 314608 442102
rect 314288 441978 314608 442046
rect 314288 441922 314358 441978
rect 314414 441922 314482 441978
rect 314538 441922 314608 441978
rect 314288 441888 314608 441922
rect 345008 442350 345328 442384
rect 345008 442294 345078 442350
rect 345134 442294 345202 442350
rect 345258 442294 345328 442350
rect 345008 442226 345328 442294
rect 345008 442170 345078 442226
rect 345134 442170 345202 442226
rect 345258 442170 345328 442226
rect 345008 442102 345328 442170
rect 345008 442046 345078 442102
rect 345134 442046 345202 442102
rect 345258 442046 345328 442102
rect 345008 441978 345328 442046
rect 345008 441922 345078 441978
rect 345134 441922 345202 441978
rect 345258 441922 345328 441978
rect 345008 441888 345328 441922
rect 375728 442350 376048 442384
rect 375728 442294 375798 442350
rect 375854 442294 375922 442350
rect 375978 442294 376048 442350
rect 375728 442226 376048 442294
rect 375728 442170 375798 442226
rect 375854 442170 375922 442226
rect 375978 442170 376048 442226
rect 375728 442102 376048 442170
rect 375728 442046 375798 442102
rect 375854 442046 375922 442102
rect 375978 442046 376048 442102
rect 375728 441978 376048 442046
rect 375728 441922 375798 441978
rect 375854 441922 375922 441978
rect 375978 441922 376048 441978
rect 375728 441888 376048 441922
rect 406448 442350 406768 442384
rect 406448 442294 406518 442350
rect 406574 442294 406642 442350
rect 406698 442294 406768 442350
rect 406448 442226 406768 442294
rect 406448 442170 406518 442226
rect 406574 442170 406642 442226
rect 406698 442170 406768 442226
rect 406448 442102 406768 442170
rect 406448 442046 406518 442102
rect 406574 442046 406642 442102
rect 406698 442046 406768 442102
rect 406448 441978 406768 442046
rect 406448 441922 406518 441978
rect 406574 441922 406642 441978
rect 406698 441922 406768 441978
rect 406448 441888 406768 441922
rect 437168 442350 437488 442384
rect 437168 442294 437238 442350
rect 437294 442294 437362 442350
rect 437418 442294 437488 442350
rect 437168 442226 437488 442294
rect 437168 442170 437238 442226
rect 437294 442170 437362 442226
rect 437418 442170 437488 442226
rect 437168 442102 437488 442170
rect 437168 442046 437238 442102
rect 437294 442046 437362 442102
rect 437418 442046 437488 442102
rect 437168 441978 437488 442046
rect 437168 441922 437238 441978
rect 437294 441922 437362 441978
rect 437418 441922 437488 441978
rect 437168 441888 437488 441922
rect 467888 442350 468208 442384
rect 467888 442294 467958 442350
rect 468014 442294 468082 442350
rect 468138 442294 468208 442350
rect 467888 442226 468208 442294
rect 467888 442170 467958 442226
rect 468014 442170 468082 442226
rect 468138 442170 468208 442226
rect 467888 442102 468208 442170
rect 467888 442046 467958 442102
rect 468014 442046 468082 442102
rect 468138 442046 468208 442102
rect 467888 441978 468208 442046
rect 467888 441922 467958 441978
rect 468014 441922 468082 441978
rect 468138 441922 468208 441978
rect 467888 441888 468208 441922
rect 498608 442350 498928 442384
rect 498608 442294 498678 442350
rect 498734 442294 498802 442350
rect 498858 442294 498928 442350
rect 498608 442226 498928 442294
rect 498608 442170 498678 442226
rect 498734 442170 498802 442226
rect 498858 442170 498928 442226
rect 498608 442102 498928 442170
rect 498608 442046 498678 442102
rect 498734 442046 498802 442102
rect 498858 442046 498928 442102
rect 498608 441978 498928 442046
rect 498608 441922 498678 441978
rect 498734 441922 498802 441978
rect 498858 441922 498928 441978
rect 498608 441888 498928 441922
rect 529328 442350 529648 442384
rect 529328 442294 529398 442350
rect 529454 442294 529522 442350
rect 529578 442294 529648 442350
rect 529328 442226 529648 442294
rect 529328 442170 529398 442226
rect 529454 442170 529522 442226
rect 529578 442170 529648 442226
rect 529328 442102 529648 442170
rect 529328 442046 529398 442102
rect 529454 442046 529522 442102
rect 529578 442046 529648 442102
rect 529328 441978 529648 442046
rect 529328 441922 529398 441978
rect 529454 441922 529522 441978
rect 529578 441922 529648 441978
rect 529328 441888 529648 441922
rect 53168 436350 53488 436384
rect 53168 436294 53238 436350
rect 53294 436294 53362 436350
rect 53418 436294 53488 436350
rect 53168 436226 53488 436294
rect 53168 436170 53238 436226
rect 53294 436170 53362 436226
rect 53418 436170 53488 436226
rect 53168 436102 53488 436170
rect 53168 436046 53238 436102
rect 53294 436046 53362 436102
rect 53418 436046 53488 436102
rect 53168 435978 53488 436046
rect 53168 435922 53238 435978
rect 53294 435922 53362 435978
rect 53418 435922 53488 435978
rect 53168 435888 53488 435922
rect 83888 436350 84208 436384
rect 83888 436294 83958 436350
rect 84014 436294 84082 436350
rect 84138 436294 84208 436350
rect 83888 436226 84208 436294
rect 83888 436170 83958 436226
rect 84014 436170 84082 436226
rect 84138 436170 84208 436226
rect 83888 436102 84208 436170
rect 83888 436046 83958 436102
rect 84014 436046 84082 436102
rect 84138 436046 84208 436102
rect 83888 435978 84208 436046
rect 83888 435922 83958 435978
rect 84014 435922 84082 435978
rect 84138 435922 84208 435978
rect 83888 435888 84208 435922
rect 114608 436350 114928 436384
rect 114608 436294 114678 436350
rect 114734 436294 114802 436350
rect 114858 436294 114928 436350
rect 114608 436226 114928 436294
rect 114608 436170 114678 436226
rect 114734 436170 114802 436226
rect 114858 436170 114928 436226
rect 114608 436102 114928 436170
rect 114608 436046 114678 436102
rect 114734 436046 114802 436102
rect 114858 436046 114928 436102
rect 114608 435978 114928 436046
rect 114608 435922 114678 435978
rect 114734 435922 114802 435978
rect 114858 435922 114928 435978
rect 114608 435888 114928 435922
rect 145328 436350 145648 436384
rect 145328 436294 145398 436350
rect 145454 436294 145522 436350
rect 145578 436294 145648 436350
rect 145328 436226 145648 436294
rect 145328 436170 145398 436226
rect 145454 436170 145522 436226
rect 145578 436170 145648 436226
rect 145328 436102 145648 436170
rect 145328 436046 145398 436102
rect 145454 436046 145522 436102
rect 145578 436046 145648 436102
rect 145328 435978 145648 436046
rect 145328 435922 145398 435978
rect 145454 435922 145522 435978
rect 145578 435922 145648 435978
rect 145328 435888 145648 435922
rect 176048 436350 176368 436384
rect 176048 436294 176118 436350
rect 176174 436294 176242 436350
rect 176298 436294 176368 436350
rect 176048 436226 176368 436294
rect 176048 436170 176118 436226
rect 176174 436170 176242 436226
rect 176298 436170 176368 436226
rect 176048 436102 176368 436170
rect 176048 436046 176118 436102
rect 176174 436046 176242 436102
rect 176298 436046 176368 436102
rect 176048 435978 176368 436046
rect 176048 435922 176118 435978
rect 176174 435922 176242 435978
rect 176298 435922 176368 435978
rect 176048 435888 176368 435922
rect 206768 436350 207088 436384
rect 206768 436294 206838 436350
rect 206894 436294 206962 436350
rect 207018 436294 207088 436350
rect 206768 436226 207088 436294
rect 206768 436170 206838 436226
rect 206894 436170 206962 436226
rect 207018 436170 207088 436226
rect 206768 436102 207088 436170
rect 206768 436046 206838 436102
rect 206894 436046 206962 436102
rect 207018 436046 207088 436102
rect 206768 435978 207088 436046
rect 206768 435922 206838 435978
rect 206894 435922 206962 435978
rect 207018 435922 207088 435978
rect 206768 435888 207088 435922
rect 237488 436350 237808 436384
rect 237488 436294 237558 436350
rect 237614 436294 237682 436350
rect 237738 436294 237808 436350
rect 237488 436226 237808 436294
rect 237488 436170 237558 436226
rect 237614 436170 237682 436226
rect 237738 436170 237808 436226
rect 237488 436102 237808 436170
rect 237488 436046 237558 436102
rect 237614 436046 237682 436102
rect 237738 436046 237808 436102
rect 237488 435978 237808 436046
rect 237488 435922 237558 435978
rect 237614 435922 237682 435978
rect 237738 435922 237808 435978
rect 237488 435888 237808 435922
rect 268208 436350 268528 436384
rect 268208 436294 268278 436350
rect 268334 436294 268402 436350
rect 268458 436294 268528 436350
rect 268208 436226 268528 436294
rect 268208 436170 268278 436226
rect 268334 436170 268402 436226
rect 268458 436170 268528 436226
rect 268208 436102 268528 436170
rect 268208 436046 268278 436102
rect 268334 436046 268402 436102
rect 268458 436046 268528 436102
rect 268208 435978 268528 436046
rect 268208 435922 268278 435978
rect 268334 435922 268402 435978
rect 268458 435922 268528 435978
rect 268208 435888 268528 435922
rect 298928 436350 299248 436384
rect 298928 436294 298998 436350
rect 299054 436294 299122 436350
rect 299178 436294 299248 436350
rect 298928 436226 299248 436294
rect 298928 436170 298998 436226
rect 299054 436170 299122 436226
rect 299178 436170 299248 436226
rect 298928 436102 299248 436170
rect 298928 436046 298998 436102
rect 299054 436046 299122 436102
rect 299178 436046 299248 436102
rect 298928 435978 299248 436046
rect 298928 435922 298998 435978
rect 299054 435922 299122 435978
rect 299178 435922 299248 435978
rect 298928 435888 299248 435922
rect 329648 436350 329968 436384
rect 329648 436294 329718 436350
rect 329774 436294 329842 436350
rect 329898 436294 329968 436350
rect 329648 436226 329968 436294
rect 329648 436170 329718 436226
rect 329774 436170 329842 436226
rect 329898 436170 329968 436226
rect 329648 436102 329968 436170
rect 329648 436046 329718 436102
rect 329774 436046 329842 436102
rect 329898 436046 329968 436102
rect 329648 435978 329968 436046
rect 329648 435922 329718 435978
rect 329774 435922 329842 435978
rect 329898 435922 329968 435978
rect 329648 435888 329968 435922
rect 360368 436350 360688 436384
rect 360368 436294 360438 436350
rect 360494 436294 360562 436350
rect 360618 436294 360688 436350
rect 360368 436226 360688 436294
rect 360368 436170 360438 436226
rect 360494 436170 360562 436226
rect 360618 436170 360688 436226
rect 360368 436102 360688 436170
rect 360368 436046 360438 436102
rect 360494 436046 360562 436102
rect 360618 436046 360688 436102
rect 360368 435978 360688 436046
rect 360368 435922 360438 435978
rect 360494 435922 360562 435978
rect 360618 435922 360688 435978
rect 360368 435888 360688 435922
rect 391088 436350 391408 436384
rect 391088 436294 391158 436350
rect 391214 436294 391282 436350
rect 391338 436294 391408 436350
rect 391088 436226 391408 436294
rect 391088 436170 391158 436226
rect 391214 436170 391282 436226
rect 391338 436170 391408 436226
rect 391088 436102 391408 436170
rect 391088 436046 391158 436102
rect 391214 436046 391282 436102
rect 391338 436046 391408 436102
rect 391088 435978 391408 436046
rect 391088 435922 391158 435978
rect 391214 435922 391282 435978
rect 391338 435922 391408 435978
rect 391088 435888 391408 435922
rect 421808 436350 422128 436384
rect 421808 436294 421878 436350
rect 421934 436294 422002 436350
rect 422058 436294 422128 436350
rect 421808 436226 422128 436294
rect 421808 436170 421878 436226
rect 421934 436170 422002 436226
rect 422058 436170 422128 436226
rect 421808 436102 422128 436170
rect 421808 436046 421878 436102
rect 421934 436046 422002 436102
rect 422058 436046 422128 436102
rect 421808 435978 422128 436046
rect 421808 435922 421878 435978
rect 421934 435922 422002 435978
rect 422058 435922 422128 435978
rect 421808 435888 422128 435922
rect 452528 436350 452848 436384
rect 452528 436294 452598 436350
rect 452654 436294 452722 436350
rect 452778 436294 452848 436350
rect 452528 436226 452848 436294
rect 452528 436170 452598 436226
rect 452654 436170 452722 436226
rect 452778 436170 452848 436226
rect 452528 436102 452848 436170
rect 452528 436046 452598 436102
rect 452654 436046 452722 436102
rect 452778 436046 452848 436102
rect 452528 435978 452848 436046
rect 452528 435922 452598 435978
rect 452654 435922 452722 435978
rect 452778 435922 452848 435978
rect 452528 435888 452848 435922
rect 483248 436350 483568 436384
rect 483248 436294 483318 436350
rect 483374 436294 483442 436350
rect 483498 436294 483568 436350
rect 483248 436226 483568 436294
rect 483248 436170 483318 436226
rect 483374 436170 483442 436226
rect 483498 436170 483568 436226
rect 483248 436102 483568 436170
rect 483248 436046 483318 436102
rect 483374 436046 483442 436102
rect 483498 436046 483568 436102
rect 483248 435978 483568 436046
rect 483248 435922 483318 435978
rect 483374 435922 483442 435978
rect 483498 435922 483568 435978
rect 483248 435888 483568 435922
rect 513968 436350 514288 436384
rect 513968 436294 514038 436350
rect 514094 436294 514162 436350
rect 514218 436294 514288 436350
rect 513968 436226 514288 436294
rect 513968 436170 514038 436226
rect 514094 436170 514162 436226
rect 514218 436170 514288 436226
rect 513968 436102 514288 436170
rect 513968 436046 514038 436102
rect 514094 436046 514162 436102
rect 514218 436046 514288 436102
rect 513968 435978 514288 436046
rect 513968 435922 514038 435978
rect 514094 435922 514162 435978
rect 514218 435922 514288 435978
rect 513968 435888 514288 435922
rect 544688 436350 545008 436384
rect 544688 436294 544758 436350
rect 544814 436294 544882 436350
rect 544938 436294 545008 436350
rect 544688 436226 545008 436294
rect 544688 436170 544758 436226
rect 544814 436170 544882 436226
rect 544938 436170 545008 436226
rect 544688 436102 545008 436170
rect 544688 436046 544758 436102
rect 544814 436046 544882 436102
rect 544938 436046 545008 436102
rect 544688 435978 545008 436046
rect 544688 435922 544758 435978
rect 544814 435922 544882 435978
rect 544938 435922 545008 435978
rect 544688 435888 545008 435922
rect 37808 424350 38128 424384
rect 37808 424294 37878 424350
rect 37934 424294 38002 424350
rect 38058 424294 38128 424350
rect 37808 424226 38128 424294
rect 37808 424170 37878 424226
rect 37934 424170 38002 424226
rect 38058 424170 38128 424226
rect 37808 424102 38128 424170
rect 37808 424046 37878 424102
rect 37934 424046 38002 424102
rect 38058 424046 38128 424102
rect 37808 423978 38128 424046
rect 37808 423922 37878 423978
rect 37934 423922 38002 423978
rect 38058 423922 38128 423978
rect 37808 423888 38128 423922
rect 68528 424350 68848 424384
rect 68528 424294 68598 424350
rect 68654 424294 68722 424350
rect 68778 424294 68848 424350
rect 68528 424226 68848 424294
rect 68528 424170 68598 424226
rect 68654 424170 68722 424226
rect 68778 424170 68848 424226
rect 68528 424102 68848 424170
rect 68528 424046 68598 424102
rect 68654 424046 68722 424102
rect 68778 424046 68848 424102
rect 68528 423978 68848 424046
rect 68528 423922 68598 423978
rect 68654 423922 68722 423978
rect 68778 423922 68848 423978
rect 68528 423888 68848 423922
rect 99248 424350 99568 424384
rect 99248 424294 99318 424350
rect 99374 424294 99442 424350
rect 99498 424294 99568 424350
rect 99248 424226 99568 424294
rect 99248 424170 99318 424226
rect 99374 424170 99442 424226
rect 99498 424170 99568 424226
rect 99248 424102 99568 424170
rect 99248 424046 99318 424102
rect 99374 424046 99442 424102
rect 99498 424046 99568 424102
rect 99248 423978 99568 424046
rect 99248 423922 99318 423978
rect 99374 423922 99442 423978
rect 99498 423922 99568 423978
rect 99248 423888 99568 423922
rect 129968 424350 130288 424384
rect 129968 424294 130038 424350
rect 130094 424294 130162 424350
rect 130218 424294 130288 424350
rect 129968 424226 130288 424294
rect 129968 424170 130038 424226
rect 130094 424170 130162 424226
rect 130218 424170 130288 424226
rect 129968 424102 130288 424170
rect 129968 424046 130038 424102
rect 130094 424046 130162 424102
rect 130218 424046 130288 424102
rect 129968 423978 130288 424046
rect 129968 423922 130038 423978
rect 130094 423922 130162 423978
rect 130218 423922 130288 423978
rect 129968 423888 130288 423922
rect 160688 424350 161008 424384
rect 160688 424294 160758 424350
rect 160814 424294 160882 424350
rect 160938 424294 161008 424350
rect 160688 424226 161008 424294
rect 160688 424170 160758 424226
rect 160814 424170 160882 424226
rect 160938 424170 161008 424226
rect 160688 424102 161008 424170
rect 160688 424046 160758 424102
rect 160814 424046 160882 424102
rect 160938 424046 161008 424102
rect 160688 423978 161008 424046
rect 160688 423922 160758 423978
rect 160814 423922 160882 423978
rect 160938 423922 161008 423978
rect 160688 423888 161008 423922
rect 191408 424350 191728 424384
rect 191408 424294 191478 424350
rect 191534 424294 191602 424350
rect 191658 424294 191728 424350
rect 191408 424226 191728 424294
rect 191408 424170 191478 424226
rect 191534 424170 191602 424226
rect 191658 424170 191728 424226
rect 191408 424102 191728 424170
rect 191408 424046 191478 424102
rect 191534 424046 191602 424102
rect 191658 424046 191728 424102
rect 191408 423978 191728 424046
rect 191408 423922 191478 423978
rect 191534 423922 191602 423978
rect 191658 423922 191728 423978
rect 191408 423888 191728 423922
rect 222128 424350 222448 424384
rect 222128 424294 222198 424350
rect 222254 424294 222322 424350
rect 222378 424294 222448 424350
rect 222128 424226 222448 424294
rect 222128 424170 222198 424226
rect 222254 424170 222322 424226
rect 222378 424170 222448 424226
rect 222128 424102 222448 424170
rect 222128 424046 222198 424102
rect 222254 424046 222322 424102
rect 222378 424046 222448 424102
rect 222128 423978 222448 424046
rect 222128 423922 222198 423978
rect 222254 423922 222322 423978
rect 222378 423922 222448 423978
rect 222128 423888 222448 423922
rect 252848 424350 253168 424384
rect 252848 424294 252918 424350
rect 252974 424294 253042 424350
rect 253098 424294 253168 424350
rect 252848 424226 253168 424294
rect 252848 424170 252918 424226
rect 252974 424170 253042 424226
rect 253098 424170 253168 424226
rect 252848 424102 253168 424170
rect 252848 424046 252918 424102
rect 252974 424046 253042 424102
rect 253098 424046 253168 424102
rect 252848 423978 253168 424046
rect 252848 423922 252918 423978
rect 252974 423922 253042 423978
rect 253098 423922 253168 423978
rect 252848 423888 253168 423922
rect 283568 424350 283888 424384
rect 283568 424294 283638 424350
rect 283694 424294 283762 424350
rect 283818 424294 283888 424350
rect 283568 424226 283888 424294
rect 283568 424170 283638 424226
rect 283694 424170 283762 424226
rect 283818 424170 283888 424226
rect 283568 424102 283888 424170
rect 283568 424046 283638 424102
rect 283694 424046 283762 424102
rect 283818 424046 283888 424102
rect 283568 423978 283888 424046
rect 283568 423922 283638 423978
rect 283694 423922 283762 423978
rect 283818 423922 283888 423978
rect 283568 423888 283888 423922
rect 314288 424350 314608 424384
rect 314288 424294 314358 424350
rect 314414 424294 314482 424350
rect 314538 424294 314608 424350
rect 314288 424226 314608 424294
rect 314288 424170 314358 424226
rect 314414 424170 314482 424226
rect 314538 424170 314608 424226
rect 314288 424102 314608 424170
rect 314288 424046 314358 424102
rect 314414 424046 314482 424102
rect 314538 424046 314608 424102
rect 314288 423978 314608 424046
rect 314288 423922 314358 423978
rect 314414 423922 314482 423978
rect 314538 423922 314608 423978
rect 314288 423888 314608 423922
rect 345008 424350 345328 424384
rect 345008 424294 345078 424350
rect 345134 424294 345202 424350
rect 345258 424294 345328 424350
rect 345008 424226 345328 424294
rect 345008 424170 345078 424226
rect 345134 424170 345202 424226
rect 345258 424170 345328 424226
rect 345008 424102 345328 424170
rect 345008 424046 345078 424102
rect 345134 424046 345202 424102
rect 345258 424046 345328 424102
rect 345008 423978 345328 424046
rect 345008 423922 345078 423978
rect 345134 423922 345202 423978
rect 345258 423922 345328 423978
rect 345008 423888 345328 423922
rect 375728 424350 376048 424384
rect 375728 424294 375798 424350
rect 375854 424294 375922 424350
rect 375978 424294 376048 424350
rect 375728 424226 376048 424294
rect 375728 424170 375798 424226
rect 375854 424170 375922 424226
rect 375978 424170 376048 424226
rect 375728 424102 376048 424170
rect 375728 424046 375798 424102
rect 375854 424046 375922 424102
rect 375978 424046 376048 424102
rect 375728 423978 376048 424046
rect 375728 423922 375798 423978
rect 375854 423922 375922 423978
rect 375978 423922 376048 423978
rect 375728 423888 376048 423922
rect 406448 424350 406768 424384
rect 406448 424294 406518 424350
rect 406574 424294 406642 424350
rect 406698 424294 406768 424350
rect 406448 424226 406768 424294
rect 406448 424170 406518 424226
rect 406574 424170 406642 424226
rect 406698 424170 406768 424226
rect 406448 424102 406768 424170
rect 406448 424046 406518 424102
rect 406574 424046 406642 424102
rect 406698 424046 406768 424102
rect 406448 423978 406768 424046
rect 406448 423922 406518 423978
rect 406574 423922 406642 423978
rect 406698 423922 406768 423978
rect 406448 423888 406768 423922
rect 437168 424350 437488 424384
rect 437168 424294 437238 424350
rect 437294 424294 437362 424350
rect 437418 424294 437488 424350
rect 437168 424226 437488 424294
rect 437168 424170 437238 424226
rect 437294 424170 437362 424226
rect 437418 424170 437488 424226
rect 437168 424102 437488 424170
rect 437168 424046 437238 424102
rect 437294 424046 437362 424102
rect 437418 424046 437488 424102
rect 437168 423978 437488 424046
rect 437168 423922 437238 423978
rect 437294 423922 437362 423978
rect 437418 423922 437488 423978
rect 437168 423888 437488 423922
rect 467888 424350 468208 424384
rect 467888 424294 467958 424350
rect 468014 424294 468082 424350
rect 468138 424294 468208 424350
rect 467888 424226 468208 424294
rect 467888 424170 467958 424226
rect 468014 424170 468082 424226
rect 468138 424170 468208 424226
rect 467888 424102 468208 424170
rect 467888 424046 467958 424102
rect 468014 424046 468082 424102
rect 468138 424046 468208 424102
rect 467888 423978 468208 424046
rect 467888 423922 467958 423978
rect 468014 423922 468082 423978
rect 468138 423922 468208 423978
rect 467888 423888 468208 423922
rect 498608 424350 498928 424384
rect 498608 424294 498678 424350
rect 498734 424294 498802 424350
rect 498858 424294 498928 424350
rect 498608 424226 498928 424294
rect 498608 424170 498678 424226
rect 498734 424170 498802 424226
rect 498858 424170 498928 424226
rect 498608 424102 498928 424170
rect 498608 424046 498678 424102
rect 498734 424046 498802 424102
rect 498858 424046 498928 424102
rect 498608 423978 498928 424046
rect 498608 423922 498678 423978
rect 498734 423922 498802 423978
rect 498858 423922 498928 423978
rect 498608 423888 498928 423922
rect 529328 424350 529648 424384
rect 529328 424294 529398 424350
rect 529454 424294 529522 424350
rect 529578 424294 529648 424350
rect 529328 424226 529648 424294
rect 529328 424170 529398 424226
rect 529454 424170 529522 424226
rect 529578 424170 529648 424226
rect 529328 424102 529648 424170
rect 529328 424046 529398 424102
rect 529454 424046 529522 424102
rect 529578 424046 529648 424102
rect 529328 423978 529648 424046
rect 529328 423922 529398 423978
rect 529454 423922 529522 423978
rect 529578 423922 529648 423978
rect 529328 423888 529648 423922
rect 53168 418350 53488 418384
rect 53168 418294 53238 418350
rect 53294 418294 53362 418350
rect 53418 418294 53488 418350
rect 53168 418226 53488 418294
rect 53168 418170 53238 418226
rect 53294 418170 53362 418226
rect 53418 418170 53488 418226
rect 53168 418102 53488 418170
rect 53168 418046 53238 418102
rect 53294 418046 53362 418102
rect 53418 418046 53488 418102
rect 53168 417978 53488 418046
rect 53168 417922 53238 417978
rect 53294 417922 53362 417978
rect 53418 417922 53488 417978
rect 53168 417888 53488 417922
rect 83888 418350 84208 418384
rect 83888 418294 83958 418350
rect 84014 418294 84082 418350
rect 84138 418294 84208 418350
rect 83888 418226 84208 418294
rect 83888 418170 83958 418226
rect 84014 418170 84082 418226
rect 84138 418170 84208 418226
rect 83888 418102 84208 418170
rect 83888 418046 83958 418102
rect 84014 418046 84082 418102
rect 84138 418046 84208 418102
rect 83888 417978 84208 418046
rect 83888 417922 83958 417978
rect 84014 417922 84082 417978
rect 84138 417922 84208 417978
rect 83888 417888 84208 417922
rect 114608 418350 114928 418384
rect 114608 418294 114678 418350
rect 114734 418294 114802 418350
rect 114858 418294 114928 418350
rect 114608 418226 114928 418294
rect 114608 418170 114678 418226
rect 114734 418170 114802 418226
rect 114858 418170 114928 418226
rect 114608 418102 114928 418170
rect 114608 418046 114678 418102
rect 114734 418046 114802 418102
rect 114858 418046 114928 418102
rect 114608 417978 114928 418046
rect 114608 417922 114678 417978
rect 114734 417922 114802 417978
rect 114858 417922 114928 417978
rect 114608 417888 114928 417922
rect 145328 418350 145648 418384
rect 145328 418294 145398 418350
rect 145454 418294 145522 418350
rect 145578 418294 145648 418350
rect 145328 418226 145648 418294
rect 145328 418170 145398 418226
rect 145454 418170 145522 418226
rect 145578 418170 145648 418226
rect 145328 418102 145648 418170
rect 145328 418046 145398 418102
rect 145454 418046 145522 418102
rect 145578 418046 145648 418102
rect 145328 417978 145648 418046
rect 145328 417922 145398 417978
rect 145454 417922 145522 417978
rect 145578 417922 145648 417978
rect 145328 417888 145648 417922
rect 176048 418350 176368 418384
rect 176048 418294 176118 418350
rect 176174 418294 176242 418350
rect 176298 418294 176368 418350
rect 176048 418226 176368 418294
rect 176048 418170 176118 418226
rect 176174 418170 176242 418226
rect 176298 418170 176368 418226
rect 176048 418102 176368 418170
rect 176048 418046 176118 418102
rect 176174 418046 176242 418102
rect 176298 418046 176368 418102
rect 176048 417978 176368 418046
rect 176048 417922 176118 417978
rect 176174 417922 176242 417978
rect 176298 417922 176368 417978
rect 176048 417888 176368 417922
rect 206768 418350 207088 418384
rect 206768 418294 206838 418350
rect 206894 418294 206962 418350
rect 207018 418294 207088 418350
rect 206768 418226 207088 418294
rect 206768 418170 206838 418226
rect 206894 418170 206962 418226
rect 207018 418170 207088 418226
rect 206768 418102 207088 418170
rect 206768 418046 206838 418102
rect 206894 418046 206962 418102
rect 207018 418046 207088 418102
rect 206768 417978 207088 418046
rect 206768 417922 206838 417978
rect 206894 417922 206962 417978
rect 207018 417922 207088 417978
rect 206768 417888 207088 417922
rect 237488 418350 237808 418384
rect 237488 418294 237558 418350
rect 237614 418294 237682 418350
rect 237738 418294 237808 418350
rect 237488 418226 237808 418294
rect 237488 418170 237558 418226
rect 237614 418170 237682 418226
rect 237738 418170 237808 418226
rect 237488 418102 237808 418170
rect 237488 418046 237558 418102
rect 237614 418046 237682 418102
rect 237738 418046 237808 418102
rect 237488 417978 237808 418046
rect 237488 417922 237558 417978
rect 237614 417922 237682 417978
rect 237738 417922 237808 417978
rect 237488 417888 237808 417922
rect 268208 418350 268528 418384
rect 268208 418294 268278 418350
rect 268334 418294 268402 418350
rect 268458 418294 268528 418350
rect 268208 418226 268528 418294
rect 268208 418170 268278 418226
rect 268334 418170 268402 418226
rect 268458 418170 268528 418226
rect 268208 418102 268528 418170
rect 268208 418046 268278 418102
rect 268334 418046 268402 418102
rect 268458 418046 268528 418102
rect 268208 417978 268528 418046
rect 268208 417922 268278 417978
rect 268334 417922 268402 417978
rect 268458 417922 268528 417978
rect 268208 417888 268528 417922
rect 298928 418350 299248 418384
rect 298928 418294 298998 418350
rect 299054 418294 299122 418350
rect 299178 418294 299248 418350
rect 298928 418226 299248 418294
rect 298928 418170 298998 418226
rect 299054 418170 299122 418226
rect 299178 418170 299248 418226
rect 298928 418102 299248 418170
rect 298928 418046 298998 418102
rect 299054 418046 299122 418102
rect 299178 418046 299248 418102
rect 298928 417978 299248 418046
rect 298928 417922 298998 417978
rect 299054 417922 299122 417978
rect 299178 417922 299248 417978
rect 298928 417888 299248 417922
rect 329648 418350 329968 418384
rect 329648 418294 329718 418350
rect 329774 418294 329842 418350
rect 329898 418294 329968 418350
rect 329648 418226 329968 418294
rect 329648 418170 329718 418226
rect 329774 418170 329842 418226
rect 329898 418170 329968 418226
rect 329648 418102 329968 418170
rect 329648 418046 329718 418102
rect 329774 418046 329842 418102
rect 329898 418046 329968 418102
rect 329648 417978 329968 418046
rect 329648 417922 329718 417978
rect 329774 417922 329842 417978
rect 329898 417922 329968 417978
rect 329648 417888 329968 417922
rect 360368 418350 360688 418384
rect 360368 418294 360438 418350
rect 360494 418294 360562 418350
rect 360618 418294 360688 418350
rect 360368 418226 360688 418294
rect 360368 418170 360438 418226
rect 360494 418170 360562 418226
rect 360618 418170 360688 418226
rect 360368 418102 360688 418170
rect 360368 418046 360438 418102
rect 360494 418046 360562 418102
rect 360618 418046 360688 418102
rect 360368 417978 360688 418046
rect 360368 417922 360438 417978
rect 360494 417922 360562 417978
rect 360618 417922 360688 417978
rect 360368 417888 360688 417922
rect 391088 418350 391408 418384
rect 391088 418294 391158 418350
rect 391214 418294 391282 418350
rect 391338 418294 391408 418350
rect 391088 418226 391408 418294
rect 391088 418170 391158 418226
rect 391214 418170 391282 418226
rect 391338 418170 391408 418226
rect 391088 418102 391408 418170
rect 391088 418046 391158 418102
rect 391214 418046 391282 418102
rect 391338 418046 391408 418102
rect 391088 417978 391408 418046
rect 391088 417922 391158 417978
rect 391214 417922 391282 417978
rect 391338 417922 391408 417978
rect 391088 417888 391408 417922
rect 421808 418350 422128 418384
rect 421808 418294 421878 418350
rect 421934 418294 422002 418350
rect 422058 418294 422128 418350
rect 421808 418226 422128 418294
rect 421808 418170 421878 418226
rect 421934 418170 422002 418226
rect 422058 418170 422128 418226
rect 421808 418102 422128 418170
rect 421808 418046 421878 418102
rect 421934 418046 422002 418102
rect 422058 418046 422128 418102
rect 421808 417978 422128 418046
rect 421808 417922 421878 417978
rect 421934 417922 422002 417978
rect 422058 417922 422128 417978
rect 421808 417888 422128 417922
rect 452528 418350 452848 418384
rect 452528 418294 452598 418350
rect 452654 418294 452722 418350
rect 452778 418294 452848 418350
rect 452528 418226 452848 418294
rect 452528 418170 452598 418226
rect 452654 418170 452722 418226
rect 452778 418170 452848 418226
rect 452528 418102 452848 418170
rect 452528 418046 452598 418102
rect 452654 418046 452722 418102
rect 452778 418046 452848 418102
rect 452528 417978 452848 418046
rect 452528 417922 452598 417978
rect 452654 417922 452722 417978
rect 452778 417922 452848 417978
rect 452528 417888 452848 417922
rect 483248 418350 483568 418384
rect 483248 418294 483318 418350
rect 483374 418294 483442 418350
rect 483498 418294 483568 418350
rect 483248 418226 483568 418294
rect 483248 418170 483318 418226
rect 483374 418170 483442 418226
rect 483498 418170 483568 418226
rect 483248 418102 483568 418170
rect 483248 418046 483318 418102
rect 483374 418046 483442 418102
rect 483498 418046 483568 418102
rect 483248 417978 483568 418046
rect 483248 417922 483318 417978
rect 483374 417922 483442 417978
rect 483498 417922 483568 417978
rect 483248 417888 483568 417922
rect 513968 418350 514288 418384
rect 513968 418294 514038 418350
rect 514094 418294 514162 418350
rect 514218 418294 514288 418350
rect 513968 418226 514288 418294
rect 513968 418170 514038 418226
rect 514094 418170 514162 418226
rect 514218 418170 514288 418226
rect 513968 418102 514288 418170
rect 513968 418046 514038 418102
rect 514094 418046 514162 418102
rect 514218 418046 514288 418102
rect 513968 417978 514288 418046
rect 513968 417922 514038 417978
rect 514094 417922 514162 417978
rect 514218 417922 514288 417978
rect 513968 417888 514288 417922
rect 544688 418350 545008 418384
rect 544688 418294 544758 418350
rect 544814 418294 544882 418350
rect 544938 418294 545008 418350
rect 544688 418226 545008 418294
rect 544688 418170 544758 418226
rect 544814 418170 544882 418226
rect 544938 418170 545008 418226
rect 544688 418102 545008 418170
rect 544688 418046 544758 418102
rect 544814 418046 544882 418102
rect 544938 418046 545008 418102
rect 544688 417978 545008 418046
rect 544688 417922 544758 417978
rect 544814 417922 544882 417978
rect 544938 417922 545008 417978
rect 544688 417888 545008 417922
rect 37808 406350 38128 406384
rect 37808 406294 37878 406350
rect 37934 406294 38002 406350
rect 38058 406294 38128 406350
rect 37808 406226 38128 406294
rect 37808 406170 37878 406226
rect 37934 406170 38002 406226
rect 38058 406170 38128 406226
rect 37808 406102 38128 406170
rect 37808 406046 37878 406102
rect 37934 406046 38002 406102
rect 38058 406046 38128 406102
rect 37808 405978 38128 406046
rect 37808 405922 37878 405978
rect 37934 405922 38002 405978
rect 38058 405922 38128 405978
rect 37808 405888 38128 405922
rect 68528 406350 68848 406384
rect 68528 406294 68598 406350
rect 68654 406294 68722 406350
rect 68778 406294 68848 406350
rect 68528 406226 68848 406294
rect 68528 406170 68598 406226
rect 68654 406170 68722 406226
rect 68778 406170 68848 406226
rect 68528 406102 68848 406170
rect 68528 406046 68598 406102
rect 68654 406046 68722 406102
rect 68778 406046 68848 406102
rect 68528 405978 68848 406046
rect 68528 405922 68598 405978
rect 68654 405922 68722 405978
rect 68778 405922 68848 405978
rect 68528 405888 68848 405922
rect 99248 406350 99568 406384
rect 99248 406294 99318 406350
rect 99374 406294 99442 406350
rect 99498 406294 99568 406350
rect 99248 406226 99568 406294
rect 99248 406170 99318 406226
rect 99374 406170 99442 406226
rect 99498 406170 99568 406226
rect 99248 406102 99568 406170
rect 99248 406046 99318 406102
rect 99374 406046 99442 406102
rect 99498 406046 99568 406102
rect 99248 405978 99568 406046
rect 99248 405922 99318 405978
rect 99374 405922 99442 405978
rect 99498 405922 99568 405978
rect 99248 405888 99568 405922
rect 129968 406350 130288 406384
rect 129968 406294 130038 406350
rect 130094 406294 130162 406350
rect 130218 406294 130288 406350
rect 129968 406226 130288 406294
rect 129968 406170 130038 406226
rect 130094 406170 130162 406226
rect 130218 406170 130288 406226
rect 129968 406102 130288 406170
rect 129968 406046 130038 406102
rect 130094 406046 130162 406102
rect 130218 406046 130288 406102
rect 129968 405978 130288 406046
rect 129968 405922 130038 405978
rect 130094 405922 130162 405978
rect 130218 405922 130288 405978
rect 129968 405888 130288 405922
rect 160688 406350 161008 406384
rect 160688 406294 160758 406350
rect 160814 406294 160882 406350
rect 160938 406294 161008 406350
rect 160688 406226 161008 406294
rect 160688 406170 160758 406226
rect 160814 406170 160882 406226
rect 160938 406170 161008 406226
rect 160688 406102 161008 406170
rect 160688 406046 160758 406102
rect 160814 406046 160882 406102
rect 160938 406046 161008 406102
rect 160688 405978 161008 406046
rect 160688 405922 160758 405978
rect 160814 405922 160882 405978
rect 160938 405922 161008 405978
rect 160688 405888 161008 405922
rect 191408 406350 191728 406384
rect 191408 406294 191478 406350
rect 191534 406294 191602 406350
rect 191658 406294 191728 406350
rect 191408 406226 191728 406294
rect 191408 406170 191478 406226
rect 191534 406170 191602 406226
rect 191658 406170 191728 406226
rect 191408 406102 191728 406170
rect 191408 406046 191478 406102
rect 191534 406046 191602 406102
rect 191658 406046 191728 406102
rect 191408 405978 191728 406046
rect 191408 405922 191478 405978
rect 191534 405922 191602 405978
rect 191658 405922 191728 405978
rect 191408 405888 191728 405922
rect 222128 406350 222448 406384
rect 222128 406294 222198 406350
rect 222254 406294 222322 406350
rect 222378 406294 222448 406350
rect 222128 406226 222448 406294
rect 222128 406170 222198 406226
rect 222254 406170 222322 406226
rect 222378 406170 222448 406226
rect 222128 406102 222448 406170
rect 222128 406046 222198 406102
rect 222254 406046 222322 406102
rect 222378 406046 222448 406102
rect 222128 405978 222448 406046
rect 222128 405922 222198 405978
rect 222254 405922 222322 405978
rect 222378 405922 222448 405978
rect 222128 405888 222448 405922
rect 252848 406350 253168 406384
rect 252848 406294 252918 406350
rect 252974 406294 253042 406350
rect 253098 406294 253168 406350
rect 252848 406226 253168 406294
rect 252848 406170 252918 406226
rect 252974 406170 253042 406226
rect 253098 406170 253168 406226
rect 252848 406102 253168 406170
rect 252848 406046 252918 406102
rect 252974 406046 253042 406102
rect 253098 406046 253168 406102
rect 252848 405978 253168 406046
rect 252848 405922 252918 405978
rect 252974 405922 253042 405978
rect 253098 405922 253168 405978
rect 252848 405888 253168 405922
rect 283568 406350 283888 406384
rect 283568 406294 283638 406350
rect 283694 406294 283762 406350
rect 283818 406294 283888 406350
rect 283568 406226 283888 406294
rect 283568 406170 283638 406226
rect 283694 406170 283762 406226
rect 283818 406170 283888 406226
rect 283568 406102 283888 406170
rect 283568 406046 283638 406102
rect 283694 406046 283762 406102
rect 283818 406046 283888 406102
rect 283568 405978 283888 406046
rect 283568 405922 283638 405978
rect 283694 405922 283762 405978
rect 283818 405922 283888 405978
rect 283568 405888 283888 405922
rect 314288 406350 314608 406384
rect 314288 406294 314358 406350
rect 314414 406294 314482 406350
rect 314538 406294 314608 406350
rect 314288 406226 314608 406294
rect 314288 406170 314358 406226
rect 314414 406170 314482 406226
rect 314538 406170 314608 406226
rect 314288 406102 314608 406170
rect 314288 406046 314358 406102
rect 314414 406046 314482 406102
rect 314538 406046 314608 406102
rect 314288 405978 314608 406046
rect 314288 405922 314358 405978
rect 314414 405922 314482 405978
rect 314538 405922 314608 405978
rect 314288 405888 314608 405922
rect 345008 406350 345328 406384
rect 345008 406294 345078 406350
rect 345134 406294 345202 406350
rect 345258 406294 345328 406350
rect 345008 406226 345328 406294
rect 345008 406170 345078 406226
rect 345134 406170 345202 406226
rect 345258 406170 345328 406226
rect 345008 406102 345328 406170
rect 345008 406046 345078 406102
rect 345134 406046 345202 406102
rect 345258 406046 345328 406102
rect 345008 405978 345328 406046
rect 345008 405922 345078 405978
rect 345134 405922 345202 405978
rect 345258 405922 345328 405978
rect 345008 405888 345328 405922
rect 375728 406350 376048 406384
rect 375728 406294 375798 406350
rect 375854 406294 375922 406350
rect 375978 406294 376048 406350
rect 375728 406226 376048 406294
rect 375728 406170 375798 406226
rect 375854 406170 375922 406226
rect 375978 406170 376048 406226
rect 375728 406102 376048 406170
rect 375728 406046 375798 406102
rect 375854 406046 375922 406102
rect 375978 406046 376048 406102
rect 375728 405978 376048 406046
rect 375728 405922 375798 405978
rect 375854 405922 375922 405978
rect 375978 405922 376048 405978
rect 375728 405888 376048 405922
rect 406448 406350 406768 406384
rect 406448 406294 406518 406350
rect 406574 406294 406642 406350
rect 406698 406294 406768 406350
rect 406448 406226 406768 406294
rect 406448 406170 406518 406226
rect 406574 406170 406642 406226
rect 406698 406170 406768 406226
rect 406448 406102 406768 406170
rect 406448 406046 406518 406102
rect 406574 406046 406642 406102
rect 406698 406046 406768 406102
rect 406448 405978 406768 406046
rect 406448 405922 406518 405978
rect 406574 405922 406642 405978
rect 406698 405922 406768 405978
rect 406448 405888 406768 405922
rect 437168 406350 437488 406384
rect 437168 406294 437238 406350
rect 437294 406294 437362 406350
rect 437418 406294 437488 406350
rect 437168 406226 437488 406294
rect 437168 406170 437238 406226
rect 437294 406170 437362 406226
rect 437418 406170 437488 406226
rect 437168 406102 437488 406170
rect 437168 406046 437238 406102
rect 437294 406046 437362 406102
rect 437418 406046 437488 406102
rect 437168 405978 437488 406046
rect 437168 405922 437238 405978
rect 437294 405922 437362 405978
rect 437418 405922 437488 405978
rect 437168 405888 437488 405922
rect 467888 406350 468208 406384
rect 467888 406294 467958 406350
rect 468014 406294 468082 406350
rect 468138 406294 468208 406350
rect 467888 406226 468208 406294
rect 467888 406170 467958 406226
rect 468014 406170 468082 406226
rect 468138 406170 468208 406226
rect 467888 406102 468208 406170
rect 467888 406046 467958 406102
rect 468014 406046 468082 406102
rect 468138 406046 468208 406102
rect 467888 405978 468208 406046
rect 467888 405922 467958 405978
rect 468014 405922 468082 405978
rect 468138 405922 468208 405978
rect 467888 405888 468208 405922
rect 498608 406350 498928 406384
rect 498608 406294 498678 406350
rect 498734 406294 498802 406350
rect 498858 406294 498928 406350
rect 498608 406226 498928 406294
rect 498608 406170 498678 406226
rect 498734 406170 498802 406226
rect 498858 406170 498928 406226
rect 498608 406102 498928 406170
rect 498608 406046 498678 406102
rect 498734 406046 498802 406102
rect 498858 406046 498928 406102
rect 498608 405978 498928 406046
rect 498608 405922 498678 405978
rect 498734 405922 498802 405978
rect 498858 405922 498928 405978
rect 498608 405888 498928 405922
rect 529328 406350 529648 406384
rect 529328 406294 529398 406350
rect 529454 406294 529522 406350
rect 529578 406294 529648 406350
rect 529328 406226 529648 406294
rect 529328 406170 529398 406226
rect 529454 406170 529522 406226
rect 529578 406170 529648 406226
rect 529328 406102 529648 406170
rect 529328 406046 529398 406102
rect 529454 406046 529522 406102
rect 529578 406046 529648 406102
rect 529328 405978 529648 406046
rect 529328 405922 529398 405978
rect 529454 405922 529522 405978
rect 529578 405922 529648 405978
rect 529328 405888 529648 405922
rect 53168 400350 53488 400384
rect 53168 400294 53238 400350
rect 53294 400294 53362 400350
rect 53418 400294 53488 400350
rect 53168 400226 53488 400294
rect 53168 400170 53238 400226
rect 53294 400170 53362 400226
rect 53418 400170 53488 400226
rect 53168 400102 53488 400170
rect 53168 400046 53238 400102
rect 53294 400046 53362 400102
rect 53418 400046 53488 400102
rect 53168 399978 53488 400046
rect 53168 399922 53238 399978
rect 53294 399922 53362 399978
rect 53418 399922 53488 399978
rect 53168 399888 53488 399922
rect 83888 400350 84208 400384
rect 83888 400294 83958 400350
rect 84014 400294 84082 400350
rect 84138 400294 84208 400350
rect 83888 400226 84208 400294
rect 83888 400170 83958 400226
rect 84014 400170 84082 400226
rect 84138 400170 84208 400226
rect 83888 400102 84208 400170
rect 83888 400046 83958 400102
rect 84014 400046 84082 400102
rect 84138 400046 84208 400102
rect 83888 399978 84208 400046
rect 83888 399922 83958 399978
rect 84014 399922 84082 399978
rect 84138 399922 84208 399978
rect 83888 399888 84208 399922
rect 114608 400350 114928 400384
rect 114608 400294 114678 400350
rect 114734 400294 114802 400350
rect 114858 400294 114928 400350
rect 114608 400226 114928 400294
rect 114608 400170 114678 400226
rect 114734 400170 114802 400226
rect 114858 400170 114928 400226
rect 114608 400102 114928 400170
rect 114608 400046 114678 400102
rect 114734 400046 114802 400102
rect 114858 400046 114928 400102
rect 114608 399978 114928 400046
rect 114608 399922 114678 399978
rect 114734 399922 114802 399978
rect 114858 399922 114928 399978
rect 114608 399888 114928 399922
rect 145328 400350 145648 400384
rect 145328 400294 145398 400350
rect 145454 400294 145522 400350
rect 145578 400294 145648 400350
rect 145328 400226 145648 400294
rect 145328 400170 145398 400226
rect 145454 400170 145522 400226
rect 145578 400170 145648 400226
rect 145328 400102 145648 400170
rect 145328 400046 145398 400102
rect 145454 400046 145522 400102
rect 145578 400046 145648 400102
rect 145328 399978 145648 400046
rect 145328 399922 145398 399978
rect 145454 399922 145522 399978
rect 145578 399922 145648 399978
rect 145328 399888 145648 399922
rect 176048 400350 176368 400384
rect 176048 400294 176118 400350
rect 176174 400294 176242 400350
rect 176298 400294 176368 400350
rect 176048 400226 176368 400294
rect 176048 400170 176118 400226
rect 176174 400170 176242 400226
rect 176298 400170 176368 400226
rect 176048 400102 176368 400170
rect 176048 400046 176118 400102
rect 176174 400046 176242 400102
rect 176298 400046 176368 400102
rect 176048 399978 176368 400046
rect 176048 399922 176118 399978
rect 176174 399922 176242 399978
rect 176298 399922 176368 399978
rect 176048 399888 176368 399922
rect 206768 400350 207088 400384
rect 206768 400294 206838 400350
rect 206894 400294 206962 400350
rect 207018 400294 207088 400350
rect 206768 400226 207088 400294
rect 206768 400170 206838 400226
rect 206894 400170 206962 400226
rect 207018 400170 207088 400226
rect 206768 400102 207088 400170
rect 206768 400046 206838 400102
rect 206894 400046 206962 400102
rect 207018 400046 207088 400102
rect 206768 399978 207088 400046
rect 206768 399922 206838 399978
rect 206894 399922 206962 399978
rect 207018 399922 207088 399978
rect 206768 399888 207088 399922
rect 237488 400350 237808 400384
rect 237488 400294 237558 400350
rect 237614 400294 237682 400350
rect 237738 400294 237808 400350
rect 237488 400226 237808 400294
rect 237488 400170 237558 400226
rect 237614 400170 237682 400226
rect 237738 400170 237808 400226
rect 237488 400102 237808 400170
rect 237488 400046 237558 400102
rect 237614 400046 237682 400102
rect 237738 400046 237808 400102
rect 237488 399978 237808 400046
rect 237488 399922 237558 399978
rect 237614 399922 237682 399978
rect 237738 399922 237808 399978
rect 237488 399888 237808 399922
rect 268208 400350 268528 400384
rect 268208 400294 268278 400350
rect 268334 400294 268402 400350
rect 268458 400294 268528 400350
rect 268208 400226 268528 400294
rect 268208 400170 268278 400226
rect 268334 400170 268402 400226
rect 268458 400170 268528 400226
rect 268208 400102 268528 400170
rect 268208 400046 268278 400102
rect 268334 400046 268402 400102
rect 268458 400046 268528 400102
rect 268208 399978 268528 400046
rect 268208 399922 268278 399978
rect 268334 399922 268402 399978
rect 268458 399922 268528 399978
rect 268208 399888 268528 399922
rect 298928 400350 299248 400384
rect 298928 400294 298998 400350
rect 299054 400294 299122 400350
rect 299178 400294 299248 400350
rect 298928 400226 299248 400294
rect 298928 400170 298998 400226
rect 299054 400170 299122 400226
rect 299178 400170 299248 400226
rect 298928 400102 299248 400170
rect 298928 400046 298998 400102
rect 299054 400046 299122 400102
rect 299178 400046 299248 400102
rect 298928 399978 299248 400046
rect 298928 399922 298998 399978
rect 299054 399922 299122 399978
rect 299178 399922 299248 399978
rect 298928 399888 299248 399922
rect 329648 400350 329968 400384
rect 329648 400294 329718 400350
rect 329774 400294 329842 400350
rect 329898 400294 329968 400350
rect 329648 400226 329968 400294
rect 329648 400170 329718 400226
rect 329774 400170 329842 400226
rect 329898 400170 329968 400226
rect 329648 400102 329968 400170
rect 329648 400046 329718 400102
rect 329774 400046 329842 400102
rect 329898 400046 329968 400102
rect 329648 399978 329968 400046
rect 329648 399922 329718 399978
rect 329774 399922 329842 399978
rect 329898 399922 329968 399978
rect 329648 399888 329968 399922
rect 360368 400350 360688 400384
rect 360368 400294 360438 400350
rect 360494 400294 360562 400350
rect 360618 400294 360688 400350
rect 360368 400226 360688 400294
rect 360368 400170 360438 400226
rect 360494 400170 360562 400226
rect 360618 400170 360688 400226
rect 360368 400102 360688 400170
rect 360368 400046 360438 400102
rect 360494 400046 360562 400102
rect 360618 400046 360688 400102
rect 360368 399978 360688 400046
rect 360368 399922 360438 399978
rect 360494 399922 360562 399978
rect 360618 399922 360688 399978
rect 360368 399888 360688 399922
rect 391088 400350 391408 400384
rect 391088 400294 391158 400350
rect 391214 400294 391282 400350
rect 391338 400294 391408 400350
rect 391088 400226 391408 400294
rect 391088 400170 391158 400226
rect 391214 400170 391282 400226
rect 391338 400170 391408 400226
rect 391088 400102 391408 400170
rect 391088 400046 391158 400102
rect 391214 400046 391282 400102
rect 391338 400046 391408 400102
rect 391088 399978 391408 400046
rect 391088 399922 391158 399978
rect 391214 399922 391282 399978
rect 391338 399922 391408 399978
rect 391088 399888 391408 399922
rect 421808 400350 422128 400384
rect 421808 400294 421878 400350
rect 421934 400294 422002 400350
rect 422058 400294 422128 400350
rect 421808 400226 422128 400294
rect 421808 400170 421878 400226
rect 421934 400170 422002 400226
rect 422058 400170 422128 400226
rect 421808 400102 422128 400170
rect 421808 400046 421878 400102
rect 421934 400046 422002 400102
rect 422058 400046 422128 400102
rect 421808 399978 422128 400046
rect 421808 399922 421878 399978
rect 421934 399922 422002 399978
rect 422058 399922 422128 399978
rect 421808 399888 422128 399922
rect 452528 400350 452848 400384
rect 452528 400294 452598 400350
rect 452654 400294 452722 400350
rect 452778 400294 452848 400350
rect 452528 400226 452848 400294
rect 452528 400170 452598 400226
rect 452654 400170 452722 400226
rect 452778 400170 452848 400226
rect 452528 400102 452848 400170
rect 452528 400046 452598 400102
rect 452654 400046 452722 400102
rect 452778 400046 452848 400102
rect 452528 399978 452848 400046
rect 452528 399922 452598 399978
rect 452654 399922 452722 399978
rect 452778 399922 452848 399978
rect 452528 399888 452848 399922
rect 483248 400350 483568 400384
rect 483248 400294 483318 400350
rect 483374 400294 483442 400350
rect 483498 400294 483568 400350
rect 483248 400226 483568 400294
rect 483248 400170 483318 400226
rect 483374 400170 483442 400226
rect 483498 400170 483568 400226
rect 483248 400102 483568 400170
rect 483248 400046 483318 400102
rect 483374 400046 483442 400102
rect 483498 400046 483568 400102
rect 483248 399978 483568 400046
rect 483248 399922 483318 399978
rect 483374 399922 483442 399978
rect 483498 399922 483568 399978
rect 483248 399888 483568 399922
rect 513968 400350 514288 400384
rect 513968 400294 514038 400350
rect 514094 400294 514162 400350
rect 514218 400294 514288 400350
rect 513968 400226 514288 400294
rect 513968 400170 514038 400226
rect 514094 400170 514162 400226
rect 514218 400170 514288 400226
rect 513968 400102 514288 400170
rect 513968 400046 514038 400102
rect 514094 400046 514162 400102
rect 514218 400046 514288 400102
rect 513968 399978 514288 400046
rect 513968 399922 514038 399978
rect 514094 399922 514162 399978
rect 514218 399922 514288 399978
rect 513968 399888 514288 399922
rect 544688 400350 545008 400384
rect 544688 400294 544758 400350
rect 544814 400294 544882 400350
rect 544938 400294 545008 400350
rect 544688 400226 545008 400294
rect 544688 400170 544758 400226
rect 544814 400170 544882 400226
rect 544938 400170 545008 400226
rect 544688 400102 545008 400170
rect 544688 400046 544758 400102
rect 544814 400046 544882 400102
rect 544938 400046 545008 400102
rect 544688 399978 545008 400046
rect 544688 399922 544758 399978
rect 544814 399922 544882 399978
rect 544938 399922 545008 399978
rect 544688 399888 545008 399922
rect 29484 375554 29540 375564
rect 152012 394324 152068 394334
rect 29372 374546 29428 374556
rect 28476 372306 28532 372316
rect 17612 372082 17668 372092
rect 150780 372260 150836 372270
rect 150332 371476 150388 371486
rect 37712 370350 38032 370384
rect 37712 370294 37782 370350
rect 37838 370294 37906 370350
rect 37962 370294 38032 370350
rect 37712 370226 38032 370294
rect 37712 370170 37782 370226
rect 37838 370170 37906 370226
rect 37962 370170 38032 370226
rect 37712 370102 38032 370170
rect 37712 370046 37782 370102
rect 37838 370046 37906 370102
rect 37962 370046 38032 370102
rect 37712 369978 38032 370046
rect 37712 369922 37782 369978
rect 37838 369922 37906 369978
rect 37962 369922 38032 369978
rect 37712 369888 38032 369922
rect 68432 370350 68752 370384
rect 68432 370294 68502 370350
rect 68558 370294 68626 370350
rect 68682 370294 68752 370350
rect 68432 370226 68752 370294
rect 68432 370170 68502 370226
rect 68558 370170 68626 370226
rect 68682 370170 68752 370226
rect 68432 370102 68752 370170
rect 68432 370046 68502 370102
rect 68558 370046 68626 370102
rect 68682 370046 68752 370102
rect 68432 369978 68752 370046
rect 68432 369922 68502 369978
rect 68558 369922 68626 369978
rect 68682 369922 68752 369978
rect 68432 369888 68752 369922
rect 99152 370350 99472 370384
rect 99152 370294 99222 370350
rect 99278 370294 99346 370350
rect 99402 370294 99472 370350
rect 99152 370226 99472 370294
rect 99152 370170 99222 370226
rect 99278 370170 99346 370226
rect 99402 370170 99472 370226
rect 99152 370102 99472 370170
rect 99152 370046 99222 370102
rect 99278 370046 99346 370102
rect 99402 370046 99472 370102
rect 99152 369978 99472 370046
rect 99152 369922 99222 369978
rect 99278 369922 99346 369978
rect 99402 369922 99472 369978
rect 99152 369888 99472 369922
rect 129872 370350 130192 370384
rect 129872 370294 129942 370350
rect 129998 370294 130066 370350
rect 130122 370294 130192 370350
rect 129872 370226 130192 370294
rect 129872 370170 129942 370226
rect 129998 370170 130066 370226
rect 130122 370170 130192 370226
rect 129872 370102 130192 370170
rect 129872 370046 129942 370102
rect 129998 370046 130066 370102
rect 130122 370046 130192 370102
rect 129872 369978 130192 370046
rect 129872 369922 129942 369978
rect 129998 369922 130066 369978
rect 130122 369922 130192 369978
rect 129872 369888 130192 369922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 4172 347508 4228 361172
rect 4172 347442 4228 347452
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect 5418 346350 6038 363922
rect 22352 364350 22672 364384
rect 22352 364294 22422 364350
rect 22478 364294 22546 364350
rect 22602 364294 22672 364350
rect 22352 364226 22672 364294
rect 22352 364170 22422 364226
rect 22478 364170 22546 364226
rect 22602 364170 22672 364226
rect 22352 364102 22672 364170
rect 22352 364046 22422 364102
rect 22478 364046 22546 364102
rect 22602 364046 22672 364102
rect 22352 363978 22672 364046
rect 22352 363922 22422 363978
rect 22478 363922 22546 363978
rect 22602 363922 22672 363978
rect 22352 363888 22672 363922
rect 53072 364350 53392 364384
rect 53072 364294 53142 364350
rect 53198 364294 53266 364350
rect 53322 364294 53392 364350
rect 53072 364226 53392 364294
rect 53072 364170 53142 364226
rect 53198 364170 53266 364226
rect 53322 364170 53392 364226
rect 53072 364102 53392 364170
rect 53072 364046 53142 364102
rect 53198 364046 53266 364102
rect 53322 364046 53392 364102
rect 53072 363978 53392 364046
rect 53072 363922 53142 363978
rect 53198 363922 53266 363978
rect 53322 363922 53392 363978
rect 53072 363888 53392 363922
rect 83792 364350 84112 364384
rect 83792 364294 83862 364350
rect 83918 364294 83986 364350
rect 84042 364294 84112 364350
rect 83792 364226 84112 364294
rect 83792 364170 83862 364226
rect 83918 364170 83986 364226
rect 84042 364170 84112 364226
rect 83792 364102 84112 364170
rect 83792 364046 83862 364102
rect 83918 364046 83986 364102
rect 84042 364046 84112 364102
rect 83792 363978 84112 364046
rect 83792 363922 83862 363978
rect 83918 363922 83986 363978
rect 84042 363922 84112 363978
rect 83792 363888 84112 363922
rect 114512 364350 114832 364384
rect 114512 364294 114582 364350
rect 114638 364294 114706 364350
rect 114762 364294 114832 364350
rect 114512 364226 114832 364294
rect 114512 364170 114582 364226
rect 114638 364170 114706 364226
rect 114762 364170 114832 364226
rect 114512 364102 114832 364170
rect 114512 364046 114582 364102
rect 114638 364046 114706 364102
rect 114762 364046 114832 364102
rect 114512 363978 114832 364046
rect 114512 363922 114582 363978
rect 114638 363922 114706 363978
rect 114762 363922 114832 363978
rect 114512 363888 114832 363922
rect 145232 364350 145552 364384
rect 145232 364294 145302 364350
rect 145358 364294 145426 364350
rect 145482 364294 145552 364350
rect 145232 364226 145552 364294
rect 145232 364170 145302 364226
rect 145358 364170 145426 364226
rect 145482 364170 145552 364226
rect 145232 364102 145552 364170
rect 145232 364046 145302 364102
rect 145358 364046 145426 364102
rect 145482 364046 145552 364102
rect 145232 363978 145552 364046
rect 145232 363922 145302 363978
rect 145358 363922 145426 363978
rect 145482 363922 145552 363978
rect 145232 363888 145552 363922
rect 37712 352350 38032 352384
rect 37712 352294 37782 352350
rect 37838 352294 37906 352350
rect 37962 352294 38032 352350
rect 37712 352226 38032 352294
rect 37712 352170 37782 352226
rect 37838 352170 37906 352226
rect 37962 352170 38032 352226
rect 37712 352102 38032 352170
rect 37712 352046 37782 352102
rect 37838 352046 37906 352102
rect 37962 352046 38032 352102
rect 37712 351978 38032 352046
rect 37712 351922 37782 351978
rect 37838 351922 37906 351978
rect 37962 351922 38032 351978
rect 37712 351888 38032 351922
rect 68432 352350 68752 352384
rect 68432 352294 68502 352350
rect 68558 352294 68626 352350
rect 68682 352294 68752 352350
rect 68432 352226 68752 352294
rect 68432 352170 68502 352226
rect 68558 352170 68626 352226
rect 68682 352170 68752 352226
rect 68432 352102 68752 352170
rect 68432 352046 68502 352102
rect 68558 352046 68626 352102
rect 68682 352046 68752 352102
rect 68432 351978 68752 352046
rect 68432 351922 68502 351978
rect 68558 351922 68626 351978
rect 68682 351922 68752 351978
rect 68432 351888 68752 351922
rect 99152 352350 99472 352384
rect 99152 352294 99222 352350
rect 99278 352294 99346 352350
rect 99402 352294 99472 352350
rect 99152 352226 99472 352294
rect 99152 352170 99222 352226
rect 99278 352170 99346 352226
rect 99402 352170 99472 352226
rect 99152 352102 99472 352170
rect 99152 352046 99222 352102
rect 99278 352046 99346 352102
rect 99402 352046 99472 352102
rect 99152 351978 99472 352046
rect 99152 351922 99222 351978
rect 99278 351922 99346 351978
rect 99402 351922 99472 351978
rect 99152 351888 99472 351922
rect 129872 352350 130192 352384
rect 129872 352294 129942 352350
rect 129998 352294 130066 352350
rect 130122 352294 130192 352350
rect 129872 352226 130192 352294
rect 129872 352170 129942 352226
rect 129998 352170 130066 352226
rect 130122 352170 130192 352226
rect 129872 352102 130192 352170
rect 129872 352046 129942 352102
rect 129998 352046 130066 352102
rect 130122 352046 130192 352102
rect 129872 351978 130192 352046
rect 129872 351922 129942 351978
rect 129998 351922 130066 351978
rect 130122 351922 130192 351978
rect 129872 351888 130192 351922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5418 328350 6038 345922
rect 22352 346350 22672 346384
rect 22352 346294 22422 346350
rect 22478 346294 22546 346350
rect 22602 346294 22672 346350
rect 22352 346226 22672 346294
rect 22352 346170 22422 346226
rect 22478 346170 22546 346226
rect 22602 346170 22672 346226
rect 22352 346102 22672 346170
rect 22352 346046 22422 346102
rect 22478 346046 22546 346102
rect 22602 346046 22672 346102
rect 22352 345978 22672 346046
rect 22352 345922 22422 345978
rect 22478 345922 22546 345978
rect 22602 345922 22672 345978
rect 22352 345888 22672 345922
rect 53072 346350 53392 346384
rect 53072 346294 53142 346350
rect 53198 346294 53266 346350
rect 53322 346294 53392 346350
rect 53072 346226 53392 346294
rect 53072 346170 53142 346226
rect 53198 346170 53266 346226
rect 53322 346170 53392 346226
rect 53072 346102 53392 346170
rect 53072 346046 53142 346102
rect 53198 346046 53266 346102
rect 53322 346046 53392 346102
rect 53072 345978 53392 346046
rect 53072 345922 53142 345978
rect 53198 345922 53266 345978
rect 53322 345922 53392 345978
rect 53072 345888 53392 345922
rect 83792 346350 84112 346384
rect 83792 346294 83862 346350
rect 83918 346294 83986 346350
rect 84042 346294 84112 346350
rect 83792 346226 84112 346294
rect 83792 346170 83862 346226
rect 83918 346170 83986 346226
rect 84042 346170 84112 346226
rect 83792 346102 84112 346170
rect 83792 346046 83862 346102
rect 83918 346046 83986 346102
rect 84042 346046 84112 346102
rect 83792 345978 84112 346046
rect 83792 345922 83862 345978
rect 83918 345922 83986 345978
rect 84042 345922 84112 345978
rect 83792 345888 84112 345922
rect 114512 346350 114832 346384
rect 114512 346294 114582 346350
rect 114638 346294 114706 346350
rect 114762 346294 114832 346350
rect 114512 346226 114832 346294
rect 114512 346170 114582 346226
rect 114638 346170 114706 346226
rect 114762 346170 114832 346226
rect 114512 346102 114832 346170
rect 114512 346046 114582 346102
rect 114638 346046 114706 346102
rect 114762 346046 114832 346102
rect 114512 345978 114832 346046
rect 114512 345922 114582 345978
rect 114638 345922 114706 345978
rect 114762 345922 114832 345978
rect 114512 345888 114832 345922
rect 145232 346350 145552 346384
rect 145232 346294 145302 346350
rect 145358 346294 145426 346350
rect 145482 346294 145552 346350
rect 145232 346226 145552 346294
rect 145232 346170 145302 346226
rect 145358 346170 145426 346226
rect 145482 346170 145552 346226
rect 145232 346102 145552 346170
rect 145232 346046 145302 346102
rect 145358 346046 145426 346102
rect 145482 346046 145552 346102
rect 145232 345978 145552 346046
rect 145232 345922 145302 345978
rect 145358 345922 145426 345978
rect 145482 345922 145552 345978
rect 145232 345888 145552 345922
rect 37712 334350 38032 334384
rect 37712 334294 37782 334350
rect 37838 334294 37906 334350
rect 37962 334294 38032 334350
rect 37712 334226 38032 334294
rect 37712 334170 37782 334226
rect 37838 334170 37906 334226
rect 37962 334170 38032 334226
rect 37712 334102 38032 334170
rect 37712 334046 37782 334102
rect 37838 334046 37906 334102
rect 37962 334046 38032 334102
rect 37712 333978 38032 334046
rect 37712 333922 37782 333978
rect 37838 333922 37906 333978
rect 37962 333922 38032 333978
rect 37712 333888 38032 333922
rect 68432 334350 68752 334384
rect 68432 334294 68502 334350
rect 68558 334294 68626 334350
rect 68682 334294 68752 334350
rect 68432 334226 68752 334294
rect 68432 334170 68502 334226
rect 68558 334170 68626 334226
rect 68682 334170 68752 334226
rect 68432 334102 68752 334170
rect 68432 334046 68502 334102
rect 68558 334046 68626 334102
rect 68682 334046 68752 334102
rect 68432 333978 68752 334046
rect 68432 333922 68502 333978
rect 68558 333922 68626 333978
rect 68682 333922 68752 333978
rect 68432 333888 68752 333922
rect 99152 334350 99472 334384
rect 99152 334294 99222 334350
rect 99278 334294 99346 334350
rect 99402 334294 99472 334350
rect 99152 334226 99472 334294
rect 99152 334170 99222 334226
rect 99278 334170 99346 334226
rect 99402 334170 99472 334226
rect 99152 334102 99472 334170
rect 99152 334046 99222 334102
rect 99278 334046 99346 334102
rect 99402 334046 99472 334102
rect 99152 333978 99472 334046
rect 99152 333922 99222 333978
rect 99278 333922 99346 333978
rect 99402 333922 99472 333978
rect 99152 333888 99472 333922
rect 129872 334350 130192 334384
rect 129872 334294 129942 334350
rect 129998 334294 130066 334350
rect 130122 334294 130192 334350
rect 129872 334226 130192 334294
rect 129872 334170 129942 334226
rect 129998 334170 130066 334226
rect 130122 334170 130192 334226
rect 129872 334102 130192 334170
rect 129872 334046 129942 334102
rect 129998 334046 130066 334102
rect 130122 334046 130192 334102
rect 129872 333978 130192 334046
rect 129872 333922 129942 333978
rect 129998 333922 130066 333978
rect 130122 333922 130192 333978
rect 129872 333888 130192 333922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect 3388 319060 3444 319070
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect 2492 276724 2548 276734
rect 2492 16324 2548 276668
rect 3388 36932 3444 319004
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 3388 36866 3444 36876
rect 3500 290836 3556 290846
rect 3500 23492 3556 290780
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 4172 262612 4228 262622
rect 4172 31948 4228 262556
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 3500 23426 3556 23436
rect 4060 31892 4228 31948
rect 4284 234388 4340 234398
rect 4060 21028 4116 31892
rect 4060 20962 4116 20972
rect 4172 26628 4228 26638
rect 4172 17578 4228 26572
rect 4284 19236 4340 234332
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 7532 333172 7588 333182
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 4284 19170 4340 19180
rect 4396 177940 4452 177950
rect 4396 17780 4452 177884
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 4508 149716 4564 149726
rect 4508 26628 4564 149660
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 4508 26562 4564 26572
rect 4620 135604 4676 135614
rect 4396 17714 4452 17724
rect 4508 26404 4564 26414
rect 4172 17522 4452 17578
rect 4172 16772 4228 16782
rect 4172 16678 4228 16716
rect 4172 16612 4228 16622
rect 4396 16548 4452 17522
rect 4396 16482 4452 16492
rect 4508 16436 4564 26348
rect 4620 18004 4676 135548
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 4732 65044 4788 65054
rect 4732 26404 4788 64988
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 4732 26338 4788 26348
rect 4844 50932 4900 50942
rect 4844 26218 4900 50876
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 4620 17938 4676 17948
rect 4732 26162 4900 26218
rect 4956 36820 5012 36830
rect 4732 17892 4788 26162
rect 4956 26038 5012 36764
rect 4844 25982 5012 26038
rect 4844 19348 4900 25982
rect 4844 19282 4900 19292
rect 4956 22708 5012 22718
rect 4956 18340 5012 22652
rect 4956 18274 5012 18284
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 4732 17826 4788 17836
rect 4508 16370 4564 16380
rect 2492 16258 2548 16268
rect 4172 14420 4228 14430
rect 4172 8820 4228 14364
rect 4172 8754 4228 8764
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 4350 6038 21922
rect 6188 192052 6244 192062
rect 6188 18452 6244 191996
rect 7532 20020 7588 333116
rect 22352 328350 22672 328384
rect 22352 328294 22422 328350
rect 22478 328294 22546 328350
rect 22602 328294 22672 328350
rect 22352 328226 22672 328294
rect 22352 328170 22422 328226
rect 22478 328170 22546 328226
rect 22602 328170 22672 328226
rect 22352 328102 22672 328170
rect 22352 328046 22422 328102
rect 22478 328046 22546 328102
rect 22602 328046 22672 328102
rect 22352 327978 22672 328046
rect 22352 327922 22422 327978
rect 22478 327922 22546 327978
rect 22602 327922 22672 327978
rect 22352 327888 22672 327922
rect 53072 328350 53392 328384
rect 53072 328294 53142 328350
rect 53198 328294 53266 328350
rect 53322 328294 53392 328350
rect 53072 328226 53392 328294
rect 53072 328170 53142 328226
rect 53198 328170 53266 328226
rect 53322 328170 53392 328226
rect 53072 328102 53392 328170
rect 53072 328046 53142 328102
rect 53198 328046 53266 328102
rect 53322 328046 53392 328102
rect 53072 327978 53392 328046
rect 53072 327922 53142 327978
rect 53198 327922 53266 327978
rect 53322 327922 53392 327978
rect 53072 327888 53392 327922
rect 83792 328350 84112 328384
rect 83792 328294 83862 328350
rect 83918 328294 83986 328350
rect 84042 328294 84112 328350
rect 83792 328226 84112 328294
rect 83792 328170 83862 328226
rect 83918 328170 83986 328226
rect 84042 328170 84112 328226
rect 83792 328102 84112 328170
rect 83792 328046 83862 328102
rect 83918 328046 83986 328102
rect 84042 328046 84112 328102
rect 83792 327978 84112 328046
rect 83792 327922 83862 327978
rect 83918 327922 83986 327978
rect 84042 327922 84112 327978
rect 83792 327888 84112 327922
rect 114512 328350 114832 328384
rect 114512 328294 114582 328350
rect 114638 328294 114706 328350
rect 114762 328294 114832 328350
rect 114512 328226 114832 328294
rect 114512 328170 114582 328226
rect 114638 328170 114706 328226
rect 114762 328170 114832 328226
rect 114512 328102 114832 328170
rect 114512 328046 114582 328102
rect 114638 328046 114706 328102
rect 114762 328046 114832 328102
rect 114512 327978 114832 328046
rect 114512 327922 114582 327978
rect 114638 327922 114706 327978
rect 114762 327922 114832 327978
rect 114512 327888 114832 327922
rect 145232 328350 145552 328384
rect 145232 328294 145302 328350
rect 145358 328294 145426 328350
rect 145482 328294 145552 328350
rect 145232 328226 145552 328294
rect 145232 328170 145302 328226
rect 145358 328170 145426 328226
rect 145482 328170 145552 328226
rect 145232 328102 145552 328170
rect 145232 328046 145302 328102
rect 145358 328046 145426 328102
rect 145482 328046 145552 328102
rect 145232 327978 145552 328046
rect 145232 327922 145302 327978
rect 145358 327922 145426 327978
rect 145482 327922 145552 327978
rect 145232 327888 145552 327922
rect 37712 316350 38032 316384
rect 37712 316294 37782 316350
rect 37838 316294 37906 316350
rect 37962 316294 38032 316350
rect 37712 316226 38032 316294
rect 37712 316170 37782 316226
rect 37838 316170 37906 316226
rect 37962 316170 38032 316226
rect 37712 316102 38032 316170
rect 37712 316046 37782 316102
rect 37838 316046 37906 316102
rect 37962 316046 38032 316102
rect 37712 315978 38032 316046
rect 37712 315922 37782 315978
rect 37838 315922 37906 315978
rect 37962 315922 38032 315978
rect 37712 315888 38032 315922
rect 68432 316350 68752 316384
rect 68432 316294 68502 316350
rect 68558 316294 68626 316350
rect 68682 316294 68752 316350
rect 68432 316226 68752 316294
rect 68432 316170 68502 316226
rect 68558 316170 68626 316226
rect 68682 316170 68752 316226
rect 68432 316102 68752 316170
rect 68432 316046 68502 316102
rect 68558 316046 68626 316102
rect 68682 316046 68752 316102
rect 68432 315978 68752 316046
rect 68432 315922 68502 315978
rect 68558 315922 68626 315978
rect 68682 315922 68752 315978
rect 68432 315888 68752 315922
rect 99152 316350 99472 316384
rect 99152 316294 99222 316350
rect 99278 316294 99346 316350
rect 99402 316294 99472 316350
rect 99152 316226 99472 316294
rect 99152 316170 99222 316226
rect 99278 316170 99346 316226
rect 99402 316170 99472 316226
rect 99152 316102 99472 316170
rect 99152 316046 99222 316102
rect 99278 316046 99346 316102
rect 99402 316046 99472 316102
rect 99152 315978 99472 316046
rect 99152 315922 99222 315978
rect 99278 315922 99346 315978
rect 99402 315922 99472 315978
rect 99152 315888 99472 315922
rect 129872 316350 130192 316384
rect 129872 316294 129942 316350
rect 129998 316294 130066 316350
rect 130122 316294 130192 316350
rect 129872 316226 130192 316294
rect 129872 316170 129942 316226
rect 129998 316170 130066 316226
rect 130122 316170 130192 316226
rect 129872 316102 130192 316170
rect 129872 316046 129942 316102
rect 129998 316046 130066 316102
rect 130122 316046 130192 316102
rect 129872 315978 130192 316046
rect 129872 315922 129942 315978
rect 129998 315922 130066 315978
rect 130122 315922 130192 315978
rect 129872 315888 130192 315922
rect 22352 310350 22672 310384
rect 22352 310294 22422 310350
rect 22478 310294 22546 310350
rect 22602 310294 22672 310350
rect 22352 310226 22672 310294
rect 22352 310170 22422 310226
rect 22478 310170 22546 310226
rect 22602 310170 22672 310226
rect 22352 310102 22672 310170
rect 22352 310046 22422 310102
rect 22478 310046 22546 310102
rect 22602 310046 22672 310102
rect 22352 309978 22672 310046
rect 22352 309922 22422 309978
rect 22478 309922 22546 309978
rect 22602 309922 22672 309978
rect 22352 309888 22672 309922
rect 53072 310350 53392 310384
rect 53072 310294 53142 310350
rect 53198 310294 53266 310350
rect 53322 310294 53392 310350
rect 53072 310226 53392 310294
rect 53072 310170 53142 310226
rect 53198 310170 53266 310226
rect 53322 310170 53392 310226
rect 53072 310102 53392 310170
rect 53072 310046 53142 310102
rect 53198 310046 53266 310102
rect 53322 310046 53392 310102
rect 53072 309978 53392 310046
rect 53072 309922 53142 309978
rect 53198 309922 53266 309978
rect 53322 309922 53392 309978
rect 53072 309888 53392 309922
rect 83792 310350 84112 310384
rect 83792 310294 83862 310350
rect 83918 310294 83986 310350
rect 84042 310294 84112 310350
rect 83792 310226 84112 310294
rect 83792 310170 83862 310226
rect 83918 310170 83986 310226
rect 84042 310170 84112 310226
rect 83792 310102 84112 310170
rect 83792 310046 83862 310102
rect 83918 310046 83986 310102
rect 84042 310046 84112 310102
rect 83792 309978 84112 310046
rect 83792 309922 83862 309978
rect 83918 309922 83986 309978
rect 84042 309922 84112 309978
rect 83792 309888 84112 309922
rect 114512 310350 114832 310384
rect 114512 310294 114582 310350
rect 114638 310294 114706 310350
rect 114762 310294 114832 310350
rect 114512 310226 114832 310294
rect 114512 310170 114582 310226
rect 114638 310170 114706 310226
rect 114762 310170 114832 310226
rect 114512 310102 114832 310170
rect 114512 310046 114582 310102
rect 114638 310046 114706 310102
rect 114762 310046 114832 310102
rect 114512 309978 114832 310046
rect 114512 309922 114582 309978
rect 114638 309922 114706 309978
rect 114762 309922 114832 309978
rect 114512 309888 114832 309922
rect 145232 310350 145552 310384
rect 145232 310294 145302 310350
rect 145358 310294 145426 310350
rect 145482 310294 145552 310350
rect 145232 310226 145552 310294
rect 145232 310170 145302 310226
rect 145358 310170 145426 310226
rect 145482 310170 145552 310226
rect 145232 310102 145552 310170
rect 145232 310046 145302 310102
rect 145358 310046 145426 310102
rect 145482 310046 145552 310102
rect 145232 309978 145552 310046
rect 145232 309922 145302 309978
rect 145358 309922 145426 309978
rect 145482 309922 145552 309978
rect 145232 309888 145552 309922
rect 9212 304948 9268 304958
rect 7756 220276 7812 220286
rect 7532 19954 7588 19964
rect 7644 107380 7700 107390
rect 6188 18386 6244 18396
rect 7644 16660 7700 107324
rect 7756 20132 7812 220220
rect 7756 20066 7812 20076
rect 7980 206164 8036 206174
rect 7980 19796 8036 206108
rect 8204 121492 8260 121502
rect 8204 19908 8260 121436
rect 8204 19842 8260 19852
rect 8988 93268 9044 93278
rect 7980 19730 8036 19740
rect 8988 18228 9044 93212
rect 9212 19684 9268 304892
rect 37712 298350 38032 298384
rect 37712 298294 37782 298350
rect 37838 298294 37906 298350
rect 37962 298294 38032 298350
rect 37712 298226 38032 298294
rect 37712 298170 37782 298226
rect 37838 298170 37906 298226
rect 37962 298170 38032 298226
rect 37712 298102 38032 298170
rect 37712 298046 37782 298102
rect 37838 298046 37906 298102
rect 37962 298046 38032 298102
rect 37712 297978 38032 298046
rect 37712 297922 37782 297978
rect 37838 297922 37906 297978
rect 37962 297922 38032 297978
rect 37712 297888 38032 297922
rect 68432 298350 68752 298384
rect 68432 298294 68502 298350
rect 68558 298294 68626 298350
rect 68682 298294 68752 298350
rect 68432 298226 68752 298294
rect 68432 298170 68502 298226
rect 68558 298170 68626 298226
rect 68682 298170 68752 298226
rect 68432 298102 68752 298170
rect 68432 298046 68502 298102
rect 68558 298046 68626 298102
rect 68682 298046 68752 298102
rect 68432 297978 68752 298046
rect 68432 297922 68502 297978
rect 68558 297922 68626 297978
rect 68682 297922 68752 297978
rect 68432 297888 68752 297922
rect 99152 298350 99472 298384
rect 99152 298294 99222 298350
rect 99278 298294 99346 298350
rect 99402 298294 99472 298350
rect 99152 298226 99472 298294
rect 99152 298170 99222 298226
rect 99278 298170 99346 298226
rect 99402 298170 99472 298226
rect 99152 298102 99472 298170
rect 99152 298046 99222 298102
rect 99278 298046 99346 298102
rect 99402 298046 99472 298102
rect 99152 297978 99472 298046
rect 99152 297922 99222 297978
rect 99278 297922 99346 297978
rect 99402 297922 99472 297978
rect 99152 297888 99472 297922
rect 129872 298350 130192 298384
rect 129872 298294 129942 298350
rect 129998 298294 130066 298350
rect 130122 298294 130192 298350
rect 129872 298226 130192 298294
rect 129872 298170 129942 298226
rect 129998 298170 130066 298226
rect 130122 298170 130192 298226
rect 129872 298102 130192 298170
rect 129872 298046 129942 298102
rect 129998 298046 130066 298102
rect 130122 298046 130192 298102
rect 129872 297978 130192 298046
rect 129872 297922 129942 297978
rect 129998 297922 130066 297978
rect 130122 297922 130192 297978
rect 129872 297888 130192 297922
rect 22352 292350 22672 292384
rect 22352 292294 22422 292350
rect 22478 292294 22546 292350
rect 22602 292294 22672 292350
rect 22352 292226 22672 292294
rect 22352 292170 22422 292226
rect 22478 292170 22546 292226
rect 22602 292170 22672 292226
rect 22352 292102 22672 292170
rect 22352 292046 22422 292102
rect 22478 292046 22546 292102
rect 22602 292046 22672 292102
rect 22352 291978 22672 292046
rect 22352 291922 22422 291978
rect 22478 291922 22546 291978
rect 22602 291922 22672 291978
rect 22352 291888 22672 291922
rect 53072 292350 53392 292384
rect 53072 292294 53142 292350
rect 53198 292294 53266 292350
rect 53322 292294 53392 292350
rect 53072 292226 53392 292294
rect 53072 292170 53142 292226
rect 53198 292170 53266 292226
rect 53322 292170 53392 292226
rect 53072 292102 53392 292170
rect 53072 292046 53142 292102
rect 53198 292046 53266 292102
rect 53322 292046 53392 292102
rect 53072 291978 53392 292046
rect 53072 291922 53142 291978
rect 53198 291922 53266 291978
rect 53322 291922 53392 291978
rect 53072 291888 53392 291922
rect 83792 292350 84112 292384
rect 83792 292294 83862 292350
rect 83918 292294 83986 292350
rect 84042 292294 84112 292350
rect 83792 292226 84112 292294
rect 83792 292170 83862 292226
rect 83918 292170 83986 292226
rect 84042 292170 84112 292226
rect 83792 292102 84112 292170
rect 83792 292046 83862 292102
rect 83918 292046 83986 292102
rect 84042 292046 84112 292102
rect 83792 291978 84112 292046
rect 83792 291922 83862 291978
rect 83918 291922 83986 291978
rect 84042 291922 84112 291978
rect 83792 291888 84112 291922
rect 114512 292350 114832 292384
rect 114512 292294 114582 292350
rect 114638 292294 114706 292350
rect 114762 292294 114832 292350
rect 114512 292226 114832 292294
rect 114512 292170 114582 292226
rect 114638 292170 114706 292226
rect 114762 292170 114832 292226
rect 114512 292102 114832 292170
rect 114512 292046 114582 292102
rect 114638 292046 114706 292102
rect 114762 292046 114832 292102
rect 114512 291978 114832 292046
rect 114512 291922 114582 291978
rect 114638 291922 114706 291978
rect 114762 291922 114832 291978
rect 114512 291888 114832 291922
rect 145232 292350 145552 292384
rect 145232 292294 145302 292350
rect 145358 292294 145426 292350
rect 145482 292294 145552 292350
rect 145232 292226 145552 292294
rect 145232 292170 145302 292226
rect 145358 292170 145426 292226
rect 145482 292170 145552 292226
rect 145232 292102 145552 292170
rect 145232 292046 145302 292102
rect 145358 292046 145426 292102
rect 145482 292046 145552 292102
rect 145232 291978 145552 292046
rect 145232 291922 145302 291978
rect 145358 291922 145426 291978
rect 145482 291922 145552 291978
rect 145232 291888 145552 291922
rect 37712 280350 38032 280384
rect 37712 280294 37782 280350
rect 37838 280294 37906 280350
rect 37962 280294 38032 280350
rect 37712 280226 38032 280294
rect 37712 280170 37782 280226
rect 37838 280170 37906 280226
rect 37962 280170 38032 280226
rect 37712 280102 38032 280170
rect 37712 280046 37782 280102
rect 37838 280046 37906 280102
rect 37962 280046 38032 280102
rect 37712 279978 38032 280046
rect 37712 279922 37782 279978
rect 37838 279922 37906 279978
rect 37962 279922 38032 279978
rect 37712 279888 38032 279922
rect 68432 280350 68752 280384
rect 68432 280294 68502 280350
rect 68558 280294 68626 280350
rect 68682 280294 68752 280350
rect 68432 280226 68752 280294
rect 68432 280170 68502 280226
rect 68558 280170 68626 280226
rect 68682 280170 68752 280226
rect 68432 280102 68752 280170
rect 68432 280046 68502 280102
rect 68558 280046 68626 280102
rect 68682 280046 68752 280102
rect 68432 279978 68752 280046
rect 68432 279922 68502 279978
rect 68558 279922 68626 279978
rect 68682 279922 68752 279978
rect 68432 279888 68752 279922
rect 99152 280350 99472 280384
rect 99152 280294 99222 280350
rect 99278 280294 99346 280350
rect 99402 280294 99472 280350
rect 99152 280226 99472 280294
rect 99152 280170 99222 280226
rect 99278 280170 99346 280226
rect 99402 280170 99472 280226
rect 99152 280102 99472 280170
rect 99152 280046 99222 280102
rect 99278 280046 99346 280102
rect 99402 280046 99472 280102
rect 99152 279978 99472 280046
rect 99152 279922 99222 279978
rect 99278 279922 99346 279978
rect 99402 279922 99472 279978
rect 99152 279888 99472 279922
rect 129872 280350 130192 280384
rect 129872 280294 129942 280350
rect 129998 280294 130066 280350
rect 130122 280294 130192 280350
rect 129872 280226 130192 280294
rect 129872 280170 129942 280226
rect 129998 280170 130066 280226
rect 130122 280170 130192 280226
rect 129872 280102 130192 280170
rect 129872 280046 129942 280102
rect 129998 280046 130066 280102
rect 130122 280046 130192 280102
rect 129872 279978 130192 280046
rect 129872 279922 129942 279978
rect 129998 279922 130066 279978
rect 130122 279922 130192 279978
rect 129872 279888 130192 279922
rect 22352 274350 22672 274384
rect 22352 274294 22422 274350
rect 22478 274294 22546 274350
rect 22602 274294 22672 274350
rect 22352 274226 22672 274294
rect 22352 274170 22422 274226
rect 22478 274170 22546 274226
rect 22602 274170 22672 274226
rect 22352 274102 22672 274170
rect 22352 274046 22422 274102
rect 22478 274046 22546 274102
rect 22602 274046 22672 274102
rect 22352 273978 22672 274046
rect 22352 273922 22422 273978
rect 22478 273922 22546 273978
rect 22602 273922 22672 273978
rect 22352 273888 22672 273922
rect 53072 274350 53392 274384
rect 53072 274294 53142 274350
rect 53198 274294 53266 274350
rect 53322 274294 53392 274350
rect 53072 274226 53392 274294
rect 53072 274170 53142 274226
rect 53198 274170 53266 274226
rect 53322 274170 53392 274226
rect 53072 274102 53392 274170
rect 53072 274046 53142 274102
rect 53198 274046 53266 274102
rect 53322 274046 53392 274102
rect 53072 273978 53392 274046
rect 53072 273922 53142 273978
rect 53198 273922 53266 273978
rect 53322 273922 53392 273978
rect 53072 273888 53392 273922
rect 83792 274350 84112 274384
rect 83792 274294 83862 274350
rect 83918 274294 83986 274350
rect 84042 274294 84112 274350
rect 83792 274226 84112 274294
rect 83792 274170 83862 274226
rect 83918 274170 83986 274226
rect 84042 274170 84112 274226
rect 83792 274102 84112 274170
rect 83792 274046 83862 274102
rect 83918 274046 83986 274102
rect 84042 274046 84112 274102
rect 83792 273978 84112 274046
rect 83792 273922 83862 273978
rect 83918 273922 83986 273978
rect 84042 273922 84112 273978
rect 83792 273888 84112 273922
rect 114512 274350 114832 274384
rect 114512 274294 114582 274350
rect 114638 274294 114706 274350
rect 114762 274294 114832 274350
rect 114512 274226 114832 274294
rect 114512 274170 114582 274226
rect 114638 274170 114706 274226
rect 114762 274170 114832 274226
rect 114512 274102 114832 274170
rect 114512 274046 114582 274102
rect 114638 274046 114706 274102
rect 114762 274046 114832 274102
rect 114512 273978 114832 274046
rect 114512 273922 114582 273978
rect 114638 273922 114706 273978
rect 114762 273922 114832 273978
rect 114512 273888 114832 273922
rect 145232 274350 145552 274384
rect 145232 274294 145302 274350
rect 145358 274294 145426 274350
rect 145482 274294 145552 274350
rect 145232 274226 145552 274294
rect 145232 274170 145302 274226
rect 145358 274170 145426 274226
rect 145482 274170 145552 274226
rect 145232 274102 145552 274170
rect 145232 274046 145302 274102
rect 145358 274046 145426 274102
rect 145482 274046 145552 274102
rect 145232 273978 145552 274046
rect 145232 273922 145302 273978
rect 145358 273922 145426 273978
rect 145482 273922 145552 273978
rect 145232 273888 145552 273922
rect 37712 262350 38032 262384
rect 37712 262294 37782 262350
rect 37838 262294 37906 262350
rect 37962 262294 38032 262350
rect 37712 262226 38032 262294
rect 37712 262170 37782 262226
rect 37838 262170 37906 262226
rect 37962 262170 38032 262226
rect 37712 262102 38032 262170
rect 37712 262046 37782 262102
rect 37838 262046 37906 262102
rect 37962 262046 38032 262102
rect 37712 261978 38032 262046
rect 37712 261922 37782 261978
rect 37838 261922 37906 261978
rect 37962 261922 38032 261978
rect 37712 261888 38032 261922
rect 68432 262350 68752 262384
rect 68432 262294 68502 262350
rect 68558 262294 68626 262350
rect 68682 262294 68752 262350
rect 68432 262226 68752 262294
rect 68432 262170 68502 262226
rect 68558 262170 68626 262226
rect 68682 262170 68752 262226
rect 68432 262102 68752 262170
rect 68432 262046 68502 262102
rect 68558 262046 68626 262102
rect 68682 262046 68752 262102
rect 68432 261978 68752 262046
rect 68432 261922 68502 261978
rect 68558 261922 68626 261978
rect 68682 261922 68752 261978
rect 68432 261888 68752 261922
rect 99152 262350 99472 262384
rect 99152 262294 99222 262350
rect 99278 262294 99346 262350
rect 99402 262294 99472 262350
rect 99152 262226 99472 262294
rect 99152 262170 99222 262226
rect 99278 262170 99346 262226
rect 99402 262170 99472 262226
rect 99152 262102 99472 262170
rect 99152 262046 99222 262102
rect 99278 262046 99346 262102
rect 99402 262046 99472 262102
rect 99152 261978 99472 262046
rect 99152 261922 99222 261978
rect 99278 261922 99346 261978
rect 99402 261922 99472 261978
rect 99152 261888 99472 261922
rect 129872 262350 130192 262384
rect 129872 262294 129942 262350
rect 129998 262294 130066 262350
rect 130122 262294 130192 262350
rect 129872 262226 130192 262294
rect 129872 262170 129942 262226
rect 129998 262170 130066 262226
rect 130122 262170 130192 262226
rect 129872 262102 130192 262170
rect 129872 262046 129942 262102
rect 129998 262046 130066 262102
rect 130122 262046 130192 262102
rect 129872 261978 130192 262046
rect 129872 261922 129942 261978
rect 129998 261922 130066 261978
rect 130122 261922 130192 261978
rect 129872 261888 130192 261922
rect 22352 256350 22672 256384
rect 22352 256294 22422 256350
rect 22478 256294 22546 256350
rect 22602 256294 22672 256350
rect 22352 256226 22672 256294
rect 22352 256170 22422 256226
rect 22478 256170 22546 256226
rect 22602 256170 22672 256226
rect 22352 256102 22672 256170
rect 22352 256046 22422 256102
rect 22478 256046 22546 256102
rect 22602 256046 22672 256102
rect 22352 255978 22672 256046
rect 22352 255922 22422 255978
rect 22478 255922 22546 255978
rect 22602 255922 22672 255978
rect 22352 255888 22672 255922
rect 53072 256350 53392 256384
rect 53072 256294 53142 256350
rect 53198 256294 53266 256350
rect 53322 256294 53392 256350
rect 53072 256226 53392 256294
rect 53072 256170 53142 256226
rect 53198 256170 53266 256226
rect 53322 256170 53392 256226
rect 53072 256102 53392 256170
rect 53072 256046 53142 256102
rect 53198 256046 53266 256102
rect 53322 256046 53392 256102
rect 53072 255978 53392 256046
rect 53072 255922 53142 255978
rect 53198 255922 53266 255978
rect 53322 255922 53392 255978
rect 53072 255888 53392 255922
rect 83792 256350 84112 256384
rect 83792 256294 83862 256350
rect 83918 256294 83986 256350
rect 84042 256294 84112 256350
rect 83792 256226 84112 256294
rect 83792 256170 83862 256226
rect 83918 256170 83986 256226
rect 84042 256170 84112 256226
rect 83792 256102 84112 256170
rect 83792 256046 83862 256102
rect 83918 256046 83986 256102
rect 84042 256046 84112 256102
rect 83792 255978 84112 256046
rect 83792 255922 83862 255978
rect 83918 255922 83986 255978
rect 84042 255922 84112 255978
rect 83792 255888 84112 255922
rect 114512 256350 114832 256384
rect 114512 256294 114582 256350
rect 114638 256294 114706 256350
rect 114762 256294 114832 256350
rect 114512 256226 114832 256294
rect 114512 256170 114582 256226
rect 114638 256170 114706 256226
rect 114762 256170 114832 256226
rect 114512 256102 114832 256170
rect 114512 256046 114582 256102
rect 114638 256046 114706 256102
rect 114762 256046 114832 256102
rect 114512 255978 114832 256046
rect 114512 255922 114582 255978
rect 114638 255922 114706 255978
rect 114762 255922 114832 255978
rect 114512 255888 114832 255922
rect 145232 256350 145552 256384
rect 145232 256294 145302 256350
rect 145358 256294 145426 256350
rect 145482 256294 145552 256350
rect 145232 256226 145552 256294
rect 145232 256170 145302 256226
rect 145358 256170 145426 256226
rect 145482 256170 145552 256226
rect 145232 256102 145552 256170
rect 145232 256046 145302 256102
rect 145358 256046 145426 256102
rect 145482 256046 145552 256102
rect 145232 255978 145552 256046
rect 145232 255922 145302 255978
rect 145358 255922 145426 255978
rect 145482 255922 145552 255978
rect 145232 255888 145552 255922
rect 9884 248500 9940 248510
rect 9212 19618 9268 19628
rect 9436 163828 9492 163838
rect 9436 19460 9492 163772
rect 9660 79156 9716 79166
rect 9660 19572 9716 79100
rect 9660 19506 9716 19516
rect 9436 19394 9492 19404
rect 8988 18162 9044 18172
rect 7644 16594 7700 16604
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 10350 9758 19026
rect 9884 18116 9940 248444
rect 37712 244350 38032 244384
rect 37712 244294 37782 244350
rect 37838 244294 37906 244350
rect 37962 244294 38032 244350
rect 37712 244226 38032 244294
rect 37712 244170 37782 244226
rect 37838 244170 37906 244226
rect 37962 244170 38032 244226
rect 37712 244102 38032 244170
rect 37712 244046 37782 244102
rect 37838 244046 37906 244102
rect 37962 244046 38032 244102
rect 37712 243978 38032 244046
rect 37712 243922 37782 243978
rect 37838 243922 37906 243978
rect 37962 243922 38032 243978
rect 37712 243888 38032 243922
rect 68432 244350 68752 244384
rect 68432 244294 68502 244350
rect 68558 244294 68626 244350
rect 68682 244294 68752 244350
rect 68432 244226 68752 244294
rect 68432 244170 68502 244226
rect 68558 244170 68626 244226
rect 68682 244170 68752 244226
rect 68432 244102 68752 244170
rect 68432 244046 68502 244102
rect 68558 244046 68626 244102
rect 68682 244046 68752 244102
rect 68432 243978 68752 244046
rect 68432 243922 68502 243978
rect 68558 243922 68626 243978
rect 68682 243922 68752 243978
rect 68432 243888 68752 243922
rect 99152 244350 99472 244384
rect 99152 244294 99222 244350
rect 99278 244294 99346 244350
rect 99402 244294 99472 244350
rect 99152 244226 99472 244294
rect 99152 244170 99222 244226
rect 99278 244170 99346 244226
rect 99402 244170 99472 244226
rect 99152 244102 99472 244170
rect 99152 244046 99222 244102
rect 99278 244046 99346 244102
rect 99402 244046 99472 244102
rect 99152 243978 99472 244046
rect 99152 243922 99222 243978
rect 99278 243922 99346 243978
rect 99402 243922 99472 243978
rect 99152 243888 99472 243922
rect 129872 244350 130192 244384
rect 129872 244294 129942 244350
rect 129998 244294 130066 244350
rect 130122 244294 130192 244350
rect 129872 244226 130192 244294
rect 129872 244170 129942 244226
rect 129998 244170 130066 244226
rect 130122 244170 130192 244226
rect 129872 244102 130192 244170
rect 129872 244046 129942 244102
rect 129998 244046 130066 244102
rect 130122 244046 130192 244102
rect 129872 243978 130192 244046
rect 129872 243922 129942 243978
rect 129998 243922 130066 243978
rect 130122 243922 130192 243978
rect 129872 243888 130192 243922
rect 22352 238350 22672 238384
rect 22352 238294 22422 238350
rect 22478 238294 22546 238350
rect 22602 238294 22672 238350
rect 22352 238226 22672 238294
rect 22352 238170 22422 238226
rect 22478 238170 22546 238226
rect 22602 238170 22672 238226
rect 22352 238102 22672 238170
rect 22352 238046 22422 238102
rect 22478 238046 22546 238102
rect 22602 238046 22672 238102
rect 22352 237978 22672 238046
rect 22352 237922 22422 237978
rect 22478 237922 22546 237978
rect 22602 237922 22672 237978
rect 22352 237888 22672 237922
rect 53072 238350 53392 238384
rect 53072 238294 53142 238350
rect 53198 238294 53266 238350
rect 53322 238294 53392 238350
rect 53072 238226 53392 238294
rect 53072 238170 53142 238226
rect 53198 238170 53266 238226
rect 53322 238170 53392 238226
rect 53072 238102 53392 238170
rect 53072 238046 53142 238102
rect 53198 238046 53266 238102
rect 53322 238046 53392 238102
rect 53072 237978 53392 238046
rect 53072 237922 53142 237978
rect 53198 237922 53266 237978
rect 53322 237922 53392 237978
rect 53072 237888 53392 237922
rect 83792 238350 84112 238384
rect 83792 238294 83862 238350
rect 83918 238294 83986 238350
rect 84042 238294 84112 238350
rect 83792 238226 84112 238294
rect 83792 238170 83862 238226
rect 83918 238170 83986 238226
rect 84042 238170 84112 238226
rect 83792 238102 84112 238170
rect 83792 238046 83862 238102
rect 83918 238046 83986 238102
rect 84042 238046 84112 238102
rect 83792 237978 84112 238046
rect 83792 237922 83862 237978
rect 83918 237922 83986 237978
rect 84042 237922 84112 237978
rect 83792 237888 84112 237922
rect 114512 238350 114832 238384
rect 114512 238294 114582 238350
rect 114638 238294 114706 238350
rect 114762 238294 114832 238350
rect 114512 238226 114832 238294
rect 114512 238170 114582 238226
rect 114638 238170 114706 238226
rect 114762 238170 114832 238226
rect 114512 238102 114832 238170
rect 114512 238046 114582 238102
rect 114638 238046 114706 238102
rect 114762 238046 114832 238102
rect 114512 237978 114832 238046
rect 114512 237922 114582 237978
rect 114638 237922 114706 237978
rect 114762 237922 114832 237978
rect 114512 237888 114832 237922
rect 145232 238350 145552 238384
rect 145232 238294 145302 238350
rect 145358 238294 145426 238350
rect 145482 238294 145552 238350
rect 145232 238226 145552 238294
rect 145232 238170 145302 238226
rect 145358 238170 145426 238226
rect 145482 238170 145552 238226
rect 145232 238102 145552 238170
rect 145232 238046 145302 238102
rect 145358 238046 145426 238102
rect 145482 238046 145552 238102
rect 145232 237978 145552 238046
rect 145232 237922 145302 237978
rect 145358 237922 145426 237978
rect 145482 237922 145552 237978
rect 145232 237888 145552 237922
rect 37712 226350 38032 226384
rect 37712 226294 37782 226350
rect 37838 226294 37906 226350
rect 37962 226294 38032 226350
rect 37712 226226 38032 226294
rect 37712 226170 37782 226226
rect 37838 226170 37906 226226
rect 37962 226170 38032 226226
rect 37712 226102 38032 226170
rect 37712 226046 37782 226102
rect 37838 226046 37906 226102
rect 37962 226046 38032 226102
rect 37712 225978 38032 226046
rect 37712 225922 37782 225978
rect 37838 225922 37906 225978
rect 37962 225922 38032 225978
rect 37712 225888 38032 225922
rect 68432 226350 68752 226384
rect 68432 226294 68502 226350
rect 68558 226294 68626 226350
rect 68682 226294 68752 226350
rect 68432 226226 68752 226294
rect 68432 226170 68502 226226
rect 68558 226170 68626 226226
rect 68682 226170 68752 226226
rect 68432 226102 68752 226170
rect 68432 226046 68502 226102
rect 68558 226046 68626 226102
rect 68682 226046 68752 226102
rect 68432 225978 68752 226046
rect 68432 225922 68502 225978
rect 68558 225922 68626 225978
rect 68682 225922 68752 225978
rect 68432 225888 68752 225922
rect 99152 226350 99472 226384
rect 99152 226294 99222 226350
rect 99278 226294 99346 226350
rect 99402 226294 99472 226350
rect 99152 226226 99472 226294
rect 99152 226170 99222 226226
rect 99278 226170 99346 226226
rect 99402 226170 99472 226226
rect 99152 226102 99472 226170
rect 99152 226046 99222 226102
rect 99278 226046 99346 226102
rect 99402 226046 99472 226102
rect 99152 225978 99472 226046
rect 99152 225922 99222 225978
rect 99278 225922 99346 225978
rect 99402 225922 99472 225978
rect 99152 225888 99472 225922
rect 129872 226350 130192 226384
rect 129872 226294 129942 226350
rect 129998 226294 130066 226350
rect 130122 226294 130192 226350
rect 129872 226226 130192 226294
rect 129872 226170 129942 226226
rect 129998 226170 130066 226226
rect 130122 226170 130192 226226
rect 129872 226102 130192 226170
rect 129872 226046 129942 226102
rect 129998 226046 130066 226102
rect 130122 226046 130192 226102
rect 129872 225978 130192 226046
rect 129872 225922 129942 225978
rect 129998 225922 130066 225978
rect 130122 225922 130192 225978
rect 129872 225888 130192 225922
rect 22352 220350 22672 220384
rect 22352 220294 22422 220350
rect 22478 220294 22546 220350
rect 22602 220294 22672 220350
rect 22352 220226 22672 220294
rect 22352 220170 22422 220226
rect 22478 220170 22546 220226
rect 22602 220170 22672 220226
rect 22352 220102 22672 220170
rect 22352 220046 22422 220102
rect 22478 220046 22546 220102
rect 22602 220046 22672 220102
rect 22352 219978 22672 220046
rect 22352 219922 22422 219978
rect 22478 219922 22546 219978
rect 22602 219922 22672 219978
rect 22352 219888 22672 219922
rect 53072 220350 53392 220384
rect 53072 220294 53142 220350
rect 53198 220294 53266 220350
rect 53322 220294 53392 220350
rect 53072 220226 53392 220294
rect 53072 220170 53142 220226
rect 53198 220170 53266 220226
rect 53322 220170 53392 220226
rect 53072 220102 53392 220170
rect 53072 220046 53142 220102
rect 53198 220046 53266 220102
rect 53322 220046 53392 220102
rect 53072 219978 53392 220046
rect 53072 219922 53142 219978
rect 53198 219922 53266 219978
rect 53322 219922 53392 219978
rect 53072 219888 53392 219922
rect 83792 220350 84112 220384
rect 83792 220294 83862 220350
rect 83918 220294 83986 220350
rect 84042 220294 84112 220350
rect 83792 220226 84112 220294
rect 83792 220170 83862 220226
rect 83918 220170 83986 220226
rect 84042 220170 84112 220226
rect 83792 220102 84112 220170
rect 83792 220046 83862 220102
rect 83918 220046 83986 220102
rect 84042 220046 84112 220102
rect 83792 219978 84112 220046
rect 83792 219922 83862 219978
rect 83918 219922 83986 219978
rect 84042 219922 84112 219978
rect 83792 219888 84112 219922
rect 114512 220350 114832 220384
rect 114512 220294 114582 220350
rect 114638 220294 114706 220350
rect 114762 220294 114832 220350
rect 114512 220226 114832 220294
rect 114512 220170 114582 220226
rect 114638 220170 114706 220226
rect 114762 220170 114832 220226
rect 114512 220102 114832 220170
rect 114512 220046 114582 220102
rect 114638 220046 114706 220102
rect 114762 220046 114832 220102
rect 114512 219978 114832 220046
rect 114512 219922 114582 219978
rect 114638 219922 114706 219978
rect 114762 219922 114832 219978
rect 114512 219888 114832 219922
rect 145232 220350 145552 220384
rect 145232 220294 145302 220350
rect 145358 220294 145426 220350
rect 145482 220294 145552 220350
rect 145232 220226 145552 220294
rect 145232 220170 145302 220226
rect 145358 220170 145426 220226
rect 145482 220170 145552 220226
rect 145232 220102 145552 220170
rect 145232 220046 145302 220102
rect 145358 220046 145426 220102
rect 145482 220046 145552 220102
rect 145232 219978 145552 220046
rect 145232 219922 145302 219978
rect 145358 219922 145426 219978
rect 145482 219922 145552 219978
rect 145232 219888 145552 219922
rect 37712 208350 38032 208384
rect 37712 208294 37782 208350
rect 37838 208294 37906 208350
rect 37962 208294 38032 208350
rect 37712 208226 38032 208294
rect 37712 208170 37782 208226
rect 37838 208170 37906 208226
rect 37962 208170 38032 208226
rect 37712 208102 38032 208170
rect 37712 208046 37782 208102
rect 37838 208046 37906 208102
rect 37962 208046 38032 208102
rect 37712 207978 38032 208046
rect 37712 207922 37782 207978
rect 37838 207922 37906 207978
rect 37962 207922 38032 207978
rect 37712 207888 38032 207922
rect 68432 208350 68752 208384
rect 68432 208294 68502 208350
rect 68558 208294 68626 208350
rect 68682 208294 68752 208350
rect 68432 208226 68752 208294
rect 68432 208170 68502 208226
rect 68558 208170 68626 208226
rect 68682 208170 68752 208226
rect 68432 208102 68752 208170
rect 68432 208046 68502 208102
rect 68558 208046 68626 208102
rect 68682 208046 68752 208102
rect 68432 207978 68752 208046
rect 68432 207922 68502 207978
rect 68558 207922 68626 207978
rect 68682 207922 68752 207978
rect 68432 207888 68752 207922
rect 99152 208350 99472 208384
rect 99152 208294 99222 208350
rect 99278 208294 99346 208350
rect 99402 208294 99472 208350
rect 99152 208226 99472 208294
rect 99152 208170 99222 208226
rect 99278 208170 99346 208226
rect 99402 208170 99472 208226
rect 99152 208102 99472 208170
rect 99152 208046 99222 208102
rect 99278 208046 99346 208102
rect 99402 208046 99472 208102
rect 99152 207978 99472 208046
rect 99152 207922 99222 207978
rect 99278 207922 99346 207978
rect 99402 207922 99472 207978
rect 99152 207888 99472 207922
rect 129872 208350 130192 208384
rect 129872 208294 129942 208350
rect 129998 208294 130066 208350
rect 130122 208294 130192 208350
rect 129872 208226 130192 208294
rect 129872 208170 129942 208226
rect 129998 208170 130066 208226
rect 130122 208170 130192 208226
rect 129872 208102 130192 208170
rect 129872 208046 129942 208102
rect 129998 208046 130066 208102
rect 130122 208046 130192 208102
rect 129872 207978 130192 208046
rect 129872 207922 129942 207978
rect 129998 207922 130066 207978
rect 130122 207922 130192 207978
rect 129872 207888 130192 207922
rect 22352 202350 22672 202384
rect 22352 202294 22422 202350
rect 22478 202294 22546 202350
rect 22602 202294 22672 202350
rect 22352 202226 22672 202294
rect 22352 202170 22422 202226
rect 22478 202170 22546 202226
rect 22602 202170 22672 202226
rect 22352 202102 22672 202170
rect 22352 202046 22422 202102
rect 22478 202046 22546 202102
rect 22602 202046 22672 202102
rect 22352 201978 22672 202046
rect 22352 201922 22422 201978
rect 22478 201922 22546 201978
rect 22602 201922 22672 201978
rect 22352 201888 22672 201922
rect 53072 202350 53392 202384
rect 53072 202294 53142 202350
rect 53198 202294 53266 202350
rect 53322 202294 53392 202350
rect 53072 202226 53392 202294
rect 53072 202170 53142 202226
rect 53198 202170 53266 202226
rect 53322 202170 53392 202226
rect 53072 202102 53392 202170
rect 53072 202046 53142 202102
rect 53198 202046 53266 202102
rect 53322 202046 53392 202102
rect 53072 201978 53392 202046
rect 53072 201922 53142 201978
rect 53198 201922 53266 201978
rect 53322 201922 53392 201978
rect 53072 201888 53392 201922
rect 83792 202350 84112 202384
rect 83792 202294 83862 202350
rect 83918 202294 83986 202350
rect 84042 202294 84112 202350
rect 83792 202226 84112 202294
rect 83792 202170 83862 202226
rect 83918 202170 83986 202226
rect 84042 202170 84112 202226
rect 83792 202102 84112 202170
rect 83792 202046 83862 202102
rect 83918 202046 83986 202102
rect 84042 202046 84112 202102
rect 83792 201978 84112 202046
rect 83792 201922 83862 201978
rect 83918 201922 83986 201978
rect 84042 201922 84112 201978
rect 83792 201888 84112 201922
rect 114512 202350 114832 202384
rect 114512 202294 114582 202350
rect 114638 202294 114706 202350
rect 114762 202294 114832 202350
rect 114512 202226 114832 202294
rect 114512 202170 114582 202226
rect 114638 202170 114706 202226
rect 114762 202170 114832 202226
rect 114512 202102 114832 202170
rect 114512 202046 114582 202102
rect 114638 202046 114706 202102
rect 114762 202046 114832 202102
rect 114512 201978 114832 202046
rect 114512 201922 114582 201978
rect 114638 201922 114706 201978
rect 114762 201922 114832 201978
rect 114512 201888 114832 201922
rect 145232 202350 145552 202384
rect 145232 202294 145302 202350
rect 145358 202294 145426 202350
rect 145482 202294 145552 202350
rect 145232 202226 145552 202294
rect 145232 202170 145302 202226
rect 145358 202170 145426 202226
rect 145482 202170 145552 202226
rect 145232 202102 145552 202170
rect 145232 202046 145302 202102
rect 145358 202046 145426 202102
rect 145482 202046 145552 202102
rect 145232 201978 145552 202046
rect 145232 201922 145302 201978
rect 145358 201922 145426 201978
rect 145482 201922 145552 201978
rect 145232 201888 145552 201922
rect 37712 190350 38032 190384
rect 37712 190294 37782 190350
rect 37838 190294 37906 190350
rect 37962 190294 38032 190350
rect 37712 190226 38032 190294
rect 37712 190170 37782 190226
rect 37838 190170 37906 190226
rect 37962 190170 38032 190226
rect 37712 190102 38032 190170
rect 37712 190046 37782 190102
rect 37838 190046 37906 190102
rect 37962 190046 38032 190102
rect 37712 189978 38032 190046
rect 37712 189922 37782 189978
rect 37838 189922 37906 189978
rect 37962 189922 38032 189978
rect 37712 189888 38032 189922
rect 68432 190350 68752 190384
rect 68432 190294 68502 190350
rect 68558 190294 68626 190350
rect 68682 190294 68752 190350
rect 68432 190226 68752 190294
rect 68432 190170 68502 190226
rect 68558 190170 68626 190226
rect 68682 190170 68752 190226
rect 68432 190102 68752 190170
rect 68432 190046 68502 190102
rect 68558 190046 68626 190102
rect 68682 190046 68752 190102
rect 68432 189978 68752 190046
rect 68432 189922 68502 189978
rect 68558 189922 68626 189978
rect 68682 189922 68752 189978
rect 68432 189888 68752 189922
rect 99152 190350 99472 190384
rect 99152 190294 99222 190350
rect 99278 190294 99346 190350
rect 99402 190294 99472 190350
rect 99152 190226 99472 190294
rect 99152 190170 99222 190226
rect 99278 190170 99346 190226
rect 99402 190170 99472 190226
rect 99152 190102 99472 190170
rect 99152 190046 99222 190102
rect 99278 190046 99346 190102
rect 99402 190046 99472 190102
rect 99152 189978 99472 190046
rect 99152 189922 99222 189978
rect 99278 189922 99346 189978
rect 99402 189922 99472 189978
rect 99152 189888 99472 189922
rect 129872 190350 130192 190384
rect 129872 190294 129942 190350
rect 129998 190294 130066 190350
rect 130122 190294 130192 190350
rect 129872 190226 130192 190294
rect 129872 190170 129942 190226
rect 129998 190170 130066 190226
rect 130122 190170 130192 190226
rect 129872 190102 130192 190170
rect 129872 190046 129942 190102
rect 129998 190046 130066 190102
rect 130122 190046 130192 190102
rect 129872 189978 130192 190046
rect 129872 189922 129942 189978
rect 129998 189922 130066 189978
rect 130122 189922 130192 189978
rect 129872 189888 130192 189922
rect 22352 184350 22672 184384
rect 22352 184294 22422 184350
rect 22478 184294 22546 184350
rect 22602 184294 22672 184350
rect 22352 184226 22672 184294
rect 22352 184170 22422 184226
rect 22478 184170 22546 184226
rect 22602 184170 22672 184226
rect 22352 184102 22672 184170
rect 22352 184046 22422 184102
rect 22478 184046 22546 184102
rect 22602 184046 22672 184102
rect 22352 183978 22672 184046
rect 22352 183922 22422 183978
rect 22478 183922 22546 183978
rect 22602 183922 22672 183978
rect 22352 183888 22672 183922
rect 53072 184350 53392 184384
rect 53072 184294 53142 184350
rect 53198 184294 53266 184350
rect 53322 184294 53392 184350
rect 53072 184226 53392 184294
rect 53072 184170 53142 184226
rect 53198 184170 53266 184226
rect 53322 184170 53392 184226
rect 53072 184102 53392 184170
rect 53072 184046 53142 184102
rect 53198 184046 53266 184102
rect 53322 184046 53392 184102
rect 53072 183978 53392 184046
rect 53072 183922 53142 183978
rect 53198 183922 53266 183978
rect 53322 183922 53392 183978
rect 53072 183888 53392 183922
rect 83792 184350 84112 184384
rect 83792 184294 83862 184350
rect 83918 184294 83986 184350
rect 84042 184294 84112 184350
rect 83792 184226 84112 184294
rect 83792 184170 83862 184226
rect 83918 184170 83986 184226
rect 84042 184170 84112 184226
rect 83792 184102 84112 184170
rect 83792 184046 83862 184102
rect 83918 184046 83986 184102
rect 84042 184046 84112 184102
rect 83792 183978 84112 184046
rect 83792 183922 83862 183978
rect 83918 183922 83986 183978
rect 84042 183922 84112 183978
rect 83792 183888 84112 183922
rect 114512 184350 114832 184384
rect 114512 184294 114582 184350
rect 114638 184294 114706 184350
rect 114762 184294 114832 184350
rect 114512 184226 114832 184294
rect 114512 184170 114582 184226
rect 114638 184170 114706 184226
rect 114762 184170 114832 184226
rect 114512 184102 114832 184170
rect 114512 184046 114582 184102
rect 114638 184046 114706 184102
rect 114762 184046 114832 184102
rect 114512 183978 114832 184046
rect 114512 183922 114582 183978
rect 114638 183922 114706 183978
rect 114762 183922 114832 183978
rect 114512 183888 114832 183922
rect 145232 184350 145552 184384
rect 145232 184294 145302 184350
rect 145358 184294 145426 184350
rect 145482 184294 145552 184350
rect 145232 184226 145552 184294
rect 145232 184170 145302 184226
rect 145358 184170 145426 184226
rect 145482 184170 145552 184226
rect 145232 184102 145552 184170
rect 145232 184046 145302 184102
rect 145358 184046 145426 184102
rect 145482 184046 145552 184102
rect 145232 183978 145552 184046
rect 145232 183922 145302 183978
rect 145358 183922 145426 183978
rect 145482 183922 145552 183978
rect 145232 183888 145552 183922
rect 37712 172350 38032 172384
rect 37712 172294 37782 172350
rect 37838 172294 37906 172350
rect 37962 172294 38032 172350
rect 37712 172226 38032 172294
rect 37712 172170 37782 172226
rect 37838 172170 37906 172226
rect 37962 172170 38032 172226
rect 37712 172102 38032 172170
rect 37712 172046 37782 172102
rect 37838 172046 37906 172102
rect 37962 172046 38032 172102
rect 37712 171978 38032 172046
rect 37712 171922 37782 171978
rect 37838 171922 37906 171978
rect 37962 171922 38032 171978
rect 37712 171888 38032 171922
rect 68432 172350 68752 172384
rect 68432 172294 68502 172350
rect 68558 172294 68626 172350
rect 68682 172294 68752 172350
rect 68432 172226 68752 172294
rect 68432 172170 68502 172226
rect 68558 172170 68626 172226
rect 68682 172170 68752 172226
rect 68432 172102 68752 172170
rect 68432 172046 68502 172102
rect 68558 172046 68626 172102
rect 68682 172046 68752 172102
rect 68432 171978 68752 172046
rect 68432 171922 68502 171978
rect 68558 171922 68626 171978
rect 68682 171922 68752 171978
rect 68432 171888 68752 171922
rect 99152 172350 99472 172384
rect 99152 172294 99222 172350
rect 99278 172294 99346 172350
rect 99402 172294 99472 172350
rect 99152 172226 99472 172294
rect 99152 172170 99222 172226
rect 99278 172170 99346 172226
rect 99402 172170 99472 172226
rect 99152 172102 99472 172170
rect 99152 172046 99222 172102
rect 99278 172046 99346 172102
rect 99402 172046 99472 172102
rect 99152 171978 99472 172046
rect 99152 171922 99222 171978
rect 99278 171922 99346 171978
rect 99402 171922 99472 171978
rect 99152 171888 99472 171922
rect 129872 172350 130192 172384
rect 129872 172294 129942 172350
rect 129998 172294 130066 172350
rect 130122 172294 130192 172350
rect 129872 172226 130192 172294
rect 129872 172170 129942 172226
rect 129998 172170 130066 172226
rect 130122 172170 130192 172226
rect 129872 172102 130192 172170
rect 129872 172046 129942 172102
rect 129998 172046 130066 172102
rect 130122 172046 130192 172102
rect 129872 171978 130192 172046
rect 129872 171922 129942 171978
rect 129998 171922 130066 171978
rect 130122 171922 130192 171978
rect 129872 171888 130192 171922
rect 22352 166350 22672 166384
rect 22352 166294 22422 166350
rect 22478 166294 22546 166350
rect 22602 166294 22672 166350
rect 22352 166226 22672 166294
rect 22352 166170 22422 166226
rect 22478 166170 22546 166226
rect 22602 166170 22672 166226
rect 22352 166102 22672 166170
rect 22352 166046 22422 166102
rect 22478 166046 22546 166102
rect 22602 166046 22672 166102
rect 22352 165978 22672 166046
rect 22352 165922 22422 165978
rect 22478 165922 22546 165978
rect 22602 165922 22672 165978
rect 22352 165888 22672 165922
rect 53072 166350 53392 166384
rect 53072 166294 53142 166350
rect 53198 166294 53266 166350
rect 53322 166294 53392 166350
rect 53072 166226 53392 166294
rect 53072 166170 53142 166226
rect 53198 166170 53266 166226
rect 53322 166170 53392 166226
rect 53072 166102 53392 166170
rect 53072 166046 53142 166102
rect 53198 166046 53266 166102
rect 53322 166046 53392 166102
rect 53072 165978 53392 166046
rect 53072 165922 53142 165978
rect 53198 165922 53266 165978
rect 53322 165922 53392 165978
rect 53072 165888 53392 165922
rect 83792 166350 84112 166384
rect 83792 166294 83862 166350
rect 83918 166294 83986 166350
rect 84042 166294 84112 166350
rect 83792 166226 84112 166294
rect 83792 166170 83862 166226
rect 83918 166170 83986 166226
rect 84042 166170 84112 166226
rect 83792 166102 84112 166170
rect 83792 166046 83862 166102
rect 83918 166046 83986 166102
rect 84042 166046 84112 166102
rect 83792 165978 84112 166046
rect 83792 165922 83862 165978
rect 83918 165922 83986 165978
rect 84042 165922 84112 165978
rect 83792 165888 84112 165922
rect 114512 166350 114832 166384
rect 114512 166294 114582 166350
rect 114638 166294 114706 166350
rect 114762 166294 114832 166350
rect 114512 166226 114832 166294
rect 114512 166170 114582 166226
rect 114638 166170 114706 166226
rect 114762 166170 114832 166226
rect 114512 166102 114832 166170
rect 114512 166046 114582 166102
rect 114638 166046 114706 166102
rect 114762 166046 114832 166102
rect 114512 165978 114832 166046
rect 114512 165922 114582 165978
rect 114638 165922 114706 165978
rect 114762 165922 114832 165978
rect 114512 165888 114832 165922
rect 145232 166350 145552 166384
rect 145232 166294 145302 166350
rect 145358 166294 145426 166350
rect 145482 166294 145552 166350
rect 145232 166226 145552 166294
rect 145232 166170 145302 166226
rect 145358 166170 145426 166226
rect 145482 166170 145552 166226
rect 145232 166102 145552 166170
rect 145232 166046 145302 166102
rect 145358 166046 145426 166102
rect 145482 166046 145552 166102
rect 145232 165978 145552 166046
rect 145232 165922 145302 165978
rect 145358 165922 145426 165978
rect 145482 165922 145552 165978
rect 145232 165888 145552 165922
rect 37712 154350 38032 154384
rect 37712 154294 37782 154350
rect 37838 154294 37906 154350
rect 37962 154294 38032 154350
rect 37712 154226 38032 154294
rect 37712 154170 37782 154226
rect 37838 154170 37906 154226
rect 37962 154170 38032 154226
rect 37712 154102 38032 154170
rect 37712 154046 37782 154102
rect 37838 154046 37906 154102
rect 37962 154046 38032 154102
rect 37712 153978 38032 154046
rect 37712 153922 37782 153978
rect 37838 153922 37906 153978
rect 37962 153922 38032 153978
rect 37712 153888 38032 153922
rect 68432 154350 68752 154384
rect 68432 154294 68502 154350
rect 68558 154294 68626 154350
rect 68682 154294 68752 154350
rect 68432 154226 68752 154294
rect 68432 154170 68502 154226
rect 68558 154170 68626 154226
rect 68682 154170 68752 154226
rect 68432 154102 68752 154170
rect 68432 154046 68502 154102
rect 68558 154046 68626 154102
rect 68682 154046 68752 154102
rect 68432 153978 68752 154046
rect 68432 153922 68502 153978
rect 68558 153922 68626 153978
rect 68682 153922 68752 153978
rect 68432 153888 68752 153922
rect 99152 154350 99472 154384
rect 99152 154294 99222 154350
rect 99278 154294 99346 154350
rect 99402 154294 99472 154350
rect 99152 154226 99472 154294
rect 99152 154170 99222 154226
rect 99278 154170 99346 154226
rect 99402 154170 99472 154226
rect 99152 154102 99472 154170
rect 99152 154046 99222 154102
rect 99278 154046 99346 154102
rect 99402 154046 99472 154102
rect 99152 153978 99472 154046
rect 99152 153922 99222 153978
rect 99278 153922 99346 153978
rect 99402 153922 99472 153978
rect 99152 153888 99472 153922
rect 129872 154350 130192 154384
rect 129872 154294 129942 154350
rect 129998 154294 130066 154350
rect 130122 154294 130192 154350
rect 129872 154226 130192 154294
rect 129872 154170 129942 154226
rect 129998 154170 130066 154226
rect 130122 154170 130192 154226
rect 129872 154102 130192 154170
rect 129872 154046 129942 154102
rect 129998 154046 130066 154102
rect 130122 154046 130192 154102
rect 129872 153978 130192 154046
rect 129872 153922 129942 153978
rect 129998 153922 130066 153978
rect 130122 153922 130192 153978
rect 129872 153888 130192 153922
rect 22352 148350 22672 148384
rect 22352 148294 22422 148350
rect 22478 148294 22546 148350
rect 22602 148294 22672 148350
rect 22352 148226 22672 148294
rect 22352 148170 22422 148226
rect 22478 148170 22546 148226
rect 22602 148170 22672 148226
rect 22352 148102 22672 148170
rect 22352 148046 22422 148102
rect 22478 148046 22546 148102
rect 22602 148046 22672 148102
rect 22352 147978 22672 148046
rect 22352 147922 22422 147978
rect 22478 147922 22546 147978
rect 22602 147922 22672 147978
rect 22352 147888 22672 147922
rect 53072 148350 53392 148384
rect 53072 148294 53142 148350
rect 53198 148294 53266 148350
rect 53322 148294 53392 148350
rect 53072 148226 53392 148294
rect 53072 148170 53142 148226
rect 53198 148170 53266 148226
rect 53322 148170 53392 148226
rect 53072 148102 53392 148170
rect 53072 148046 53142 148102
rect 53198 148046 53266 148102
rect 53322 148046 53392 148102
rect 53072 147978 53392 148046
rect 53072 147922 53142 147978
rect 53198 147922 53266 147978
rect 53322 147922 53392 147978
rect 53072 147888 53392 147922
rect 83792 148350 84112 148384
rect 83792 148294 83862 148350
rect 83918 148294 83986 148350
rect 84042 148294 84112 148350
rect 83792 148226 84112 148294
rect 83792 148170 83862 148226
rect 83918 148170 83986 148226
rect 84042 148170 84112 148226
rect 83792 148102 84112 148170
rect 83792 148046 83862 148102
rect 83918 148046 83986 148102
rect 84042 148046 84112 148102
rect 83792 147978 84112 148046
rect 83792 147922 83862 147978
rect 83918 147922 83986 147978
rect 84042 147922 84112 147978
rect 83792 147888 84112 147922
rect 114512 148350 114832 148384
rect 114512 148294 114582 148350
rect 114638 148294 114706 148350
rect 114762 148294 114832 148350
rect 114512 148226 114832 148294
rect 114512 148170 114582 148226
rect 114638 148170 114706 148226
rect 114762 148170 114832 148226
rect 114512 148102 114832 148170
rect 114512 148046 114582 148102
rect 114638 148046 114706 148102
rect 114762 148046 114832 148102
rect 114512 147978 114832 148046
rect 114512 147922 114582 147978
rect 114638 147922 114706 147978
rect 114762 147922 114832 147978
rect 114512 147888 114832 147922
rect 145232 148350 145552 148384
rect 145232 148294 145302 148350
rect 145358 148294 145426 148350
rect 145482 148294 145552 148350
rect 145232 148226 145552 148294
rect 145232 148170 145302 148226
rect 145358 148170 145426 148226
rect 145482 148170 145552 148226
rect 145232 148102 145552 148170
rect 145232 148046 145302 148102
rect 145358 148046 145426 148102
rect 145482 148046 145552 148102
rect 145232 147978 145552 148046
rect 145232 147922 145302 147978
rect 145358 147922 145426 147978
rect 145482 147922 145552 147978
rect 145232 147888 145552 147922
rect 37712 136350 38032 136384
rect 37712 136294 37782 136350
rect 37838 136294 37906 136350
rect 37962 136294 38032 136350
rect 37712 136226 38032 136294
rect 37712 136170 37782 136226
rect 37838 136170 37906 136226
rect 37962 136170 38032 136226
rect 37712 136102 38032 136170
rect 37712 136046 37782 136102
rect 37838 136046 37906 136102
rect 37962 136046 38032 136102
rect 37712 135978 38032 136046
rect 37712 135922 37782 135978
rect 37838 135922 37906 135978
rect 37962 135922 38032 135978
rect 37712 135888 38032 135922
rect 68432 136350 68752 136384
rect 68432 136294 68502 136350
rect 68558 136294 68626 136350
rect 68682 136294 68752 136350
rect 68432 136226 68752 136294
rect 68432 136170 68502 136226
rect 68558 136170 68626 136226
rect 68682 136170 68752 136226
rect 68432 136102 68752 136170
rect 68432 136046 68502 136102
rect 68558 136046 68626 136102
rect 68682 136046 68752 136102
rect 68432 135978 68752 136046
rect 68432 135922 68502 135978
rect 68558 135922 68626 135978
rect 68682 135922 68752 135978
rect 68432 135888 68752 135922
rect 99152 136350 99472 136384
rect 99152 136294 99222 136350
rect 99278 136294 99346 136350
rect 99402 136294 99472 136350
rect 99152 136226 99472 136294
rect 99152 136170 99222 136226
rect 99278 136170 99346 136226
rect 99402 136170 99472 136226
rect 99152 136102 99472 136170
rect 99152 136046 99222 136102
rect 99278 136046 99346 136102
rect 99402 136046 99472 136102
rect 99152 135978 99472 136046
rect 99152 135922 99222 135978
rect 99278 135922 99346 135978
rect 99402 135922 99472 135978
rect 99152 135888 99472 135922
rect 129872 136350 130192 136384
rect 129872 136294 129942 136350
rect 129998 136294 130066 136350
rect 130122 136294 130192 136350
rect 129872 136226 130192 136294
rect 129872 136170 129942 136226
rect 129998 136170 130066 136226
rect 130122 136170 130192 136226
rect 129872 136102 130192 136170
rect 129872 136046 129942 136102
rect 129998 136046 130066 136102
rect 130122 136046 130192 136102
rect 129872 135978 130192 136046
rect 129872 135922 129942 135978
rect 129998 135922 130066 135978
rect 130122 135922 130192 135978
rect 129872 135888 130192 135922
rect 22352 130350 22672 130384
rect 22352 130294 22422 130350
rect 22478 130294 22546 130350
rect 22602 130294 22672 130350
rect 22352 130226 22672 130294
rect 22352 130170 22422 130226
rect 22478 130170 22546 130226
rect 22602 130170 22672 130226
rect 22352 130102 22672 130170
rect 22352 130046 22422 130102
rect 22478 130046 22546 130102
rect 22602 130046 22672 130102
rect 22352 129978 22672 130046
rect 22352 129922 22422 129978
rect 22478 129922 22546 129978
rect 22602 129922 22672 129978
rect 22352 129888 22672 129922
rect 53072 130350 53392 130384
rect 53072 130294 53142 130350
rect 53198 130294 53266 130350
rect 53322 130294 53392 130350
rect 53072 130226 53392 130294
rect 53072 130170 53142 130226
rect 53198 130170 53266 130226
rect 53322 130170 53392 130226
rect 53072 130102 53392 130170
rect 53072 130046 53142 130102
rect 53198 130046 53266 130102
rect 53322 130046 53392 130102
rect 53072 129978 53392 130046
rect 53072 129922 53142 129978
rect 53198 129922 53266 129978
rect 53322 129922 53392 129978
rect 53072 129888 53392 129922
rect 83792 130350 84112 130384
rect 83792 130294 83862 130350
rect 83918 130294 83986 130350
rect 84042 130294 84112 130350
rect 83792 130226 84112 130294
rect 83792 130170 83862 130226
rect 83918 130170 83986 130226
rect 84042 130170 84112 130226
rect 83792 130102 84112 130170
rect 83792 130046 83862 130102
rect 83918 130046 83986 130102
rect 84042 130046 84112 130102
rect 83792 129978 84112 130046
rect 83792 129922 83862 129978
rect 83918 129922 83986 129978
rect 84042 129922 84112 129978
rect 83792 129888 84112 129922
rect 114512 130350 114832 130384
rect 114512 130294 114582 130350
rect 114638 130294 114706 130350
rect 114762 130294 114832 130350
rect 114512 130226 114832 130294
rect 114512 130170 114582 130226
rect 114638 130170 114706 130226
rect 114762 130170 114832 130226
rect 114512 130102 114832 130170
rect 114512 130046 114582 130102
rect 114638 130046 114706 130102
rect 114762 130046 114832 130102
rect 114512 129978 114832 130046
rect 114512 129922 114582 129978
rect 114638 129922 114706 129978
rect 114762 129922 114832 129978
rect 114512 129888 114832 129922
rect 145232 130350 145552 130384
rect 145232 130294 145302 130350
rect 145358 130294 145426 130350
rect 145482 130294 145552 130350
rect 145232 130226 145552 130294
rect 145232 130170 145302 130226
rect 145358 130170 145426 130226
rect 145482 130170 145552 130226
rect 145232 130102 145552 130170
rect 145232 130046 145302 130102
rect 145358 130046 145426 130102
rect 145482 130046 145552 130102
rect 145232 129978 145552 130046
rect 145232 129922 145302 129978
rect 145358 129922 145426 129978
rect 145482 129922 145552 129978
rect 145232 129888 145552 129922
rect 37712 118350 38032 118384
rect 37712 118294 37782 118350
rect 37838 118294 37906 118350
rect 37962 118294 38032 118350
rect 37712 118226 38032 118294
rect 37712 118170 37782 118226
rect 37838 118170 37906 118226
rect 37962 118170 38032 118226
rect 37712 118102 38032 118170
rect 37712 118046 37782 118102
rect 37838 118046 37906 118102
rect 37962 118046 38032 118102
rect 37712 117978 38032 118046
rect 37712 117922 37782 117978
rect 37838 117922 37906 117978
rect 37962 117922 38032 117978
rect 37712 117888 38032 117922
rect 68432 118350 68752 118384
rect 68432 118294 68502 118350
rect 68558 118294 68626 118350
rect 68682 118294 68752 118350
rect 68432 118226 68752 118294
rect 68432 118170 68502 118226
rect 68558 118170 68626 118226
rect 68682 118170 68752 118226
rect 68432 118102 68752 118170
rect 68432 118046 68502 118102
rect 68558 118046 68626 118102
rect 68682 118046 68752 118102
rect 68432 117978 68752 118046
rect 68432 117922 68502 117978
rect 68558 117922 68626 117978
rect 68682 117922 68752 117978
rect 68432 117888 68752 117922
rect 99152 118350 99472 118384
rect 99152 118294 99222 118350
rect 99278 118294 99346 118350
rect 99402 118294 99472 118350
rect 99152 118226 99472 118294
rect 99152 118170 99222 118226
rect 99278 118170 99346 118226
rect 99402 118170 99472 118226
rect 99152 118102 99472 118170
rect 99152 118046 99222 118102
rect 99278 118046 99346 118102
rect 99402 118046 99472 118102
rect 99152 117978 99472 118046
rect 99152 117922 99222 117978
rect 99278 117922 99346 117978
rect 99402 117922 99472 117978
rect 99152 117888 99472 117922
rect 129872 118350 130192 118384
rect 129872 118294 129942 118350
rect 129998 118294 130066 118350
rect 130122 118294 130192 118350
rect 129872 118226 130192 118294
rect 129872 118170 129942 118226
rect 129998 118170 130066 118226
rect 130122 118170 130192 118226
rect 129872 118102 130192 118170
rect 129872 118046 129942 118102
rect 129998 118046 130066 118102
rect 130122 118046 130192 118102
rect 129872 117978 130192 118046
rect 129872 117922 129942 117978
rect 129998 117922 130066 117978
rect 130122 117922 130192 117978
rect 129872 117888 130192 117922
rect 22352 112350 22672 112384
rect 22352 112294 22422 112350
rect 22478 112294 22546 112350
rect 22602 112294 22672 112350
rect 22352 112226 22672 112294
rect 22352 112170 22422 112226
rect 22478 112170 22546 112226
rect 22602 112170 22672 112226
rect 22352 112102 22672 112170
rect 22352 112046 22422 112102
rect 22478 112046 22546 112102
rect 22602 112046 22672 112102
rect 22352 111978 22672 112046
rect 22352 111922 22422 111978
rect 22478 111922 22546 111978
rect 22602 111922 22672 111978
rect 22352 111888 22672 111922
rect 53072 112350 53392 112384
rect 53072 112294 53142 112350
rect 53198 112294 53266 112350
rect 53322 112294 53392 112350
rect 53072 112226 53392 112294
rect 53072 112170 53142 112226
rect 53198 112170 53266 112226
rect 53322 112170 53392 112226
rect 53072 112102 53392 112170
rect 53072 112046 53142 112102
rect 53198 112046 53266 112102
rect 53322 112046 53392 112102
rect 53072 111978 53392 112046
rect 53072 111922 53142 111978
rect 53198 111922 53266 111978
rect 53322 111922 53392 111978
rect 53072 111888 53392 111922
rect 83792 112350 84112 112384
rect 83792 112294 83862 112350
rect 83918 112294 83986 112350
rect 84042 112294 84112 112350
rect 83792 112226 84112 112294
rect 83792 112170 83862 112226
rect 83918 112170 83986 112226
rect 84042 112170 84112 112226
rect 83792 112102 84112 112170
rect 83792 112046 83862 112102
rect 83918 112046 83986 112102
rect 84042 112046 84112 112102
rect 83792 111978 84112 112046
rect 83792 111922 83862 111978
rect 83918 111922 83986 111978
rect 84042 111922 84112 111978
rect 83792 111888 84112 111922
rect 114512 112350 114832 112384
rect 114512 112294 114582 112350
rect 114638 112294 114706 112350
rect 114762 112294 114832 112350
rect 114512 112226 114832 112294
rect 114512 112170 114582 112226
rect 114638 112170 114706 112226
rect 114762 112170 114832 112226
rect 114512 112102 114832 112170
rect 114512 112046 114582 112102
rect 114638 112046 114706 112102
rect 114762 112046 114832 112102
rect 114512 111978 114832 112046
rect 114512 111922 114582 111978
rect 114638 111922 114706 111978
rect 114762 111922 114832 111978
rect 114512 111888 114832 111922
rect 145232 112350 145552 112384
rect 145232 112294 145302 112350
rect 145358 112294 145426 112350
rect 145482 112294 145552 112350
rect 145232 112226 145552 112294
rect 145232 112170 145302 112226
rect 145358 112170 145426 112226
rect 145482 112170 145552 112226
rect 145232 112102 145552 112170
rect 145232 112046 145302 112102
rect 145358 112046 145426 112102
rect 145482 112046 145552 112102
rect 145232 111978 145552 112046
rect 145232 111922 145302 111978
rect 145358 111922 145426 111978
rect 145482 111922 145552 111978
rect 145232 111888 145552 111922
rect 37712 100350 38032 100384
rect 37712 100294 37782 100350
rect 37838 100294 37906 100350
rect 37962 100294 38032 100350
rect 37712 100226 38032 100294
rect 37712 100170 37782 100226
rect 37838 100170 37906 100226
rect 37962 100170 38032 100226
rect 37712 100102 38032 100170
rect 37712 100046 37782 100102
rect 37838 100046 37906 100102
rect 37962 100046 38032 100102
rect 37712 99978 38032 100046
rect 37712 99922 37782 99978
rect 37838 99922 37906 99978
rect 37962 99922 38032 99978
rect 37712 99888 38032 99922
rect 68432 100350 68752 100384
rect 68432 100294 68502 100350
rect 68558 100294 68626 100350
rect 68682 100294 68752 100350
rect 68432 100226 68752 100294
rect 68432 100170 68502 100226
rect 68558 100170 68626 100226
rect 68682 100170 68752 100226
rect 68432 100102 68752 100170
rect 68432 100046 68502 100102
rect 68558 100046 68626 100102
rect 68682 100046 68752 100102
rect 68432 99978 68752 100046
rect 68432 99922 68502 99978
rect 68558 99922 68626 99978
rect 68682 99922 68752 99978
rect 68432 99888 68752 99922
rect 99152 100350 99472 100384
rect 99152 100294 99222 100350
rect 99278 100294 99346 100350
rect 99402 100294 99472 100350
rect 99152 100226 99472 100294
rect 99152 100170 99222 100226
rect 99278 100170 99346 100226
rect 99402 100170 99472 100226
rect 99152 100102 99472 100170
rect 99152 100046 99222 100102
rect 99278 100046 99346 100102
rect 99402 100046 99472 100102
rect 99152 99978 99472 100046
rect 99152 99922 99222 99978
rect 99278 99922 99346 99978
rect 99402 99922 99472 99978
rect 99152 99888 99472 99922
rect 129872 100350 130192 100384
rect 129872 100294 129942 100350
rect 129998 100294 130066 100350
rect 130122 100294 130192 100350
rect 129872 100226 130192 100294
rect 129872 100170 129942 100226
rect 129998 100170 130066 100226
rect 130122 100170 130192 100226
rect 129872 100102 130192 100170
rect 129872 100046 129942 100102
rect 129998 100046 130066 100102
rect 130122 100046 130192 100102
rect 129872 99978 130192 100046
rect 129872 99922 129942 99978
rect 129998 99922 130066 99978
rect 130122 99922 130192 99978
rect 129872 99888 130192 99922
rect 22352 94350 22672 94384
rect 22352 94294 22422 94350
rect 22478 94294 22546 94350
rect 22602 94294 22672 94350
rect 22352 94226 22672 94294
rect 22352 94170 22422 94226
rect 22478 94170 22546 94226
rect 22602 94170 22672 94226
rect 22352 94102 22672 94170
rect 22352 94046 22422 94102
rect 22478 94046 22546 94102
rect 22602 94046 22672 94102
rect 22352 93978 22672 94046
rect 22352 93922 22422 93978
rect 22478 93922 22546 93978
rect 22602 93922 22672 93978
rect 22352 93888 22672 93922
rect 53072 94350 53392 94384
rect 53072 94294 53142 94350
rect 53198 94294 53266 94350
rect 53322 94294 53392 94350
rect 53072 94226 53392 94294
rect 53072 94170 53142 94226
rect 53198 94170 53266 94226
rect 53322 94170 53392 94226
rect 53072 94102 53392 94170
rect 53072 94046 53142 94102
rect 53198 94046 53266 94102
rect 53322 94046 53392 94102
rect 53072 93978 53392 94046
rect 53072 93922 53142 93978
rect 53198 93922 53266 93978
rect 53322 93922 53392 93978
rect 53072 93888 53392 93922
rect 83792 94350 84112 94384
rect 83792 94294 83862 94350
rect 83918 94294 83986 94350
rect 84042 94294 84112 94350
rect 83792 94226 84112 94294
rect 83792 94170 83862 94226
rect 83918 94170 83986 94226
rect 84042 94170 84112 94226
rect 83792 94102 84112 94170
rect 83792 94046 83862 94102
rect 83918 94046 83986 94102
rect 84042 94046 84112 94102
rect 83792 93978 84112 94046
rect 83792 93922 83862 93978
rect 83918 93922 83986 93978
rect 84042 93922 84112 93978
rect 83792 93888 84112 93922
rect 114512 94350 114832 94384
rect 114512 94294 114582 94350
rect 114638 94294 114706 94350
rect 114762 94294 114832 94350
rect 114512 94226 114832 94294
rect 114512 94170 114582 94226
rect 114638 94170 114706 94226
rect 114762 94170 114832 94226
rect 114512 94102 114832 94170
rect 114512 94046 114582 94102
rect 114638 94046 114706 94102
rect 114762 94046 114832 94102
rect 114512 93978 114832 94046
rect 114512 93922 114582 93978
rect 114638 93922 114706 93978
rect 114762 93922 114832 93978
rect 114512 93888 114832 93922
rect 145232 94350 145552 94384
rect 145232 94294 145302 94350
rect 145358 94294 145426 94350
rect 145482 94294 145552 94350
rect 145232 94226 145552 94294
rect 145232 94170 145302 94226
rect 145358 94170 145426 94226
rect 145482 94170 145552 94226
rect 145232 94102 145552 94170
rect 145232 94046 145302 94102
rect 145358 94046 145426 94102
rect 145482 94046 145552 94102
rect 145232 93978 145552 94046
rect 145232 93922 145302 93978
rect 145358 93922 145426 93978
rect 145482 93922 145552 93978
rect 145232 93888 145552 93922
rect 37712 82350 38032 82384
rect 37712 82294 37782 82350
rect 37838 82294 37906 82350
rect 37962 82294 38032 82350
rect 37712 82226 38032 82294
rect 37712 82170 37782 82226
rect 37838 82170 37906 82226
rect 37962 82170 38032 82226
rect 37712 82102 38032 82170
rect 37712 82046 37782 82102
rect 37838 82046 37906 82102
rect 37962 82046 38032 82102
rect 37712 81978 38032 82046
rect 37712 81922 37782 81978
rect 37838 81922 37906 81978
rect 37962 81922 38032 81978
rect 37712 81888 38032 81922
rect 68432 82350 68752 82384
rect 68432 82294 68502 82350
rect 68558 82294 68626 82350
rect 68682 82294 68752 82350
rect 68432 82226 68752 82294
rect 68432 82170 68502 82226
rect 68558 82170 68626 82226
rect 68682 82170 68752 82226
rect 68432 82102 68752 82170
rect 68432 82046 68502 82102
rect 68558 82046 68626 82102
rect 68682 82046 68752 82102
rect 68432 81978 68752 82046
rect 68432 81922 68502 81978
rect 68558 81922 68626 81978
rect 68682 81922 68752 81978
rect 68432 81888 68752 81922
rect 99152 82350 99472 82384
rect 99152 82294 99222 82350
rect 99278 82294 99346 82350
rect 99402 82294 99472 82350
rect 99152 82226 99472 82294
rect 99152 82170 99222 82226
rect 99278 82170 99346 82226
rect 99402 82170 99472 82226
rect 99152 82102 99472 82170
rect 99152 82046 99222 82102
rect 99278 82046 99346 82102
rect 99402 82046 99472 82102
rect 99152 81978 99472 82046
rect 99152 81922 99222 81978
rect 99278 81922 99346 81978
rect 99402 81922 99472 81978
rect 99152 81888 99472 81922
rect 129872 82350 130192 82384
rect 129872 82294 129942 82350
rect 129998 82294 130066 82350
rect 130122 82294 130192 82350
rect 129872 82226 130192 82294
rect 129872 82170 129942 82226
rect 129998 82170 130066 82226
rect 130122 82170 130192 82226
rect 129872 82102 130192 82170
rect 129872 82046 129942 82102
rect 129998 82046 130066 82102
rect 130122 82046 130192 82102
rect 129872 81978 130192 82046
rect 129872 81922 129942 81978
rect 129998 81922 130066 81978
rect 130122 81922 130192 81978
rect 129872 81888 130192 81922
rect 22352 76350 22672 76384
rect 22352 76294 22422 76350
rect 22478 76294 22546 76350
rect 22602 76294 22672 76350
rect 22352 76226 22672 76294
rect 22352 76170 22422 76226
rect 22478 76170 22546 76226
rect 22602 76170 22672 76226
rect 22352 76102 22672 76170
rect 22352 76046 22422 76102
rect 22478 76046 22546 76102
rect 22602 76046 22672 76102
rect 22352 75978 22672 76046
rect 22352 75922 22422 75978
rect 22478 75922 22546 75978
rect 22602 75922 22672 75978
rect 22352 75888 22672 75922
rect 53072 76350 53392 76384
rect 53072 76294 53142 76350
rect 53198 76294 53266 76350
rect 53322 76294 53392 76350
rect 53072 76226 53392 76294
rect 53072 76170 53142 76226
rect 53198 76170 53266 76226
rect 53322 76170 53392 76226
rect 53072 76102 53392 76170
rect 53072 76046 53142 76102
rect 53198 76046 53266 76102
rect 53322 76046 53392 76102
rect 53072 75978 53392 76046
rect 53072 75922 53142 75978
rect 53198 75922 53266 75978
rect 53322 75922 53392 75978
rect 53072 75888 53392 75922
rect 83792 76350 84112 76384
rect 83792 76294 83862 76350
rect 83918 76294 83986 76350
rect 84042 76294 84112 76350
rect 83792 76226 84112 76294
rect 83792 76170 83862 76226
rect 83918 76170 83986 76226
rect 84042 76170 84112 76226
rect 83792 76102 84112 76170
rect 83792 76046 83862 76102
rect 83918 76046 83986 76102
rect 84042 76046 84112 76102
rect 83792 75978 84112 76046
rect 83792 75922 83862 75978
rect 83918 75922 83986 75978
rect 84042 75922 84112 75978
rect 83792 75888 84112 75922
rect 114512 76350 114832 76384
rect 114512 76294 114582 76350
rect 114638 76294 114706 76350
rect 114762 76294 114832 76350
rect 114512 76226 114832 76294
rect 114512 76170 114582 76226
rect 114638 76170 114706 76226
rect 114762 76170 114832 76226
rect 114512 76102 114832 76170
rect 114512 76046 114582 76102
rect 114638 76046 114706 76102
rect 114762 76046 114832 76102
rect 114512 75978 114832 76046
rect 114512 75922 114582 75978
rect 114638 75922 114706 75978
rect 114762 75922 114832 75978
rect 114512 75888 114832 75922
rect 145232 76350 145552 76384
rect 145232 76294 145302 76350
rect 145358 76294 145426 76350
rect 145482 76294 145552 76350
rect 145232 76226 145552 76294
rect 145232 76170 145302 76226
rect 145358 76170 145426 76226
rect 145482 76170 145552 76226
rect 145232 76102 145552 76170
rect 145232 76046 145302 76102
rect 145358 76046 145426 76102
rect 145482 76046 145552 76102
rect 145232 75978 145552 76046
rect 145232 75922 145302 75978
rect 145358 75922 145426 75978
rect 145482 75922 145552 75978
rect 145232 75888 145552 75922
rect 37712 64350 38032 64384
rect 37712 64294 37782 64350
rect 37838 64294 37906 64350
rect 37962 64294 38032 64350
rect 37712 64226 38032 64294
rect 37712 64170 37782 64226
rect 37838 64170 37906 64226
rect 37962 64170 38032 64226
rect 37712 64102 38032 64170
rect 37712 64046 37782 64102
rect 37838 64046 37906 64102
rect 37962 64046 38032 64102
rect 37712 63978 38032 64046
rect 37712 63922 37782 63978
rect 37838 63922 37906 63978
rect 37962 63922 38032 63978
rect 37712 63888 38032 63922
rect 68432 64350 68752 64384
rect 68432 64294 68502 64350
rect 68558 64294 68626 64350
rect 68682 64294 68752 64350
rect 68432 64226 68752 64294
rect 68432 64170 68502 64226
rect 68558 64170 68626 64226
rect 68682 64170 68752 64226
rect 68432 64102 68752 64170
rect 68432 64046 68502 64102
rect 68558 64046 68626 64102
rect 68682 64046 68752 64102
rect 68432 63978 68752 64046
rect 68432 63922 68502 63978
rect 68558 63922 68626 63978
rect 68682 63922 68752 63978
rect 68432 63888 68752 63922
rect 99152 64350 99472 64384
rect 99152 64294 99222 64350
rect 99278 64294 99346 64350
rect 99402 64294 99472 64350
rect 99152 64226 99472 64294
rect 99152 64170 99222 64226
rect 99278 64170 99346 64226
rect 99402 64170 99472 64226
rect 99152 64102 99472 64170
rect 99152 64046 99222 64102
rect 99278 64046 99346 64102
rect 99402 64046 99472 64102
rect 99152 63978 99472 64046
rect 99152 63922 99222 63978
rect 99278 63922 99346 63978
rect 99402 63922 99472 63978
rect 99152 63888 99472 63922
rect 129872 64350 130192 64384
rect 129872 64294 129942 64350
rect 129998 64294 130066 64350
rect 130122 64294 130192 64350
rect 129872 64226 130192 64294
rect 129872 64170 129942 64226
rect 129998 64170 130066 64226
rect 130122 64170 130192 64226
rect 129872 64102 130192 64170
rect 129872 64046 129942 64102
rect 129998 64046 130066 64102
rect 130122 64046 130192 64102
rect 129872 63978 130192 64046
rect 129872 63922 129942 63978
rect 129998 63922 130066 63978
rect 130122 63922 130192 63978
rect 129872 63888 130192 63922
rect 22352 58350 22672 58384
rect 22352 58294 22422 58350
rect 22478 58294 22546 58350
rect 22602 58294 22672 58350
rect 22352 58226 22672 58294
rect 22352 58170 22422 58226
rect 22478 58170 22546 58226
rect 22602 58170 22672 58226
rect 22352 58102 22672 58170
rect 22352 58046 22422 58102
rect 22478 58046 22546 58102
rect 22602 58046 22672 58102
rect 22352 57978 22672 58046
rect 22352 57922 22422 57978
rect 22478 57922 22546 57978
rect 22602 57922 22672 57978
rect 22352 57888 22672 57922
rect 53072 58350 53392 58384
rect 53072 58294 53142 58350
rect 53198 58294 53266 58350
rect 53322 58294 53392 58350
rect 53072 58226 53392 58294
rect 53072 58170 53142 58226
rect 53198 58170 53266 58226
rect 53322 58170 53392 58226
rect 53072 58102 53392 58170
rect 53072 58046 53142 58102
rect 53198 58046 53266 58102
rect 53322 58046 53392 58102
rect 53072 57978 53392 58046
rect 53072 57922 53142 57978
rect 53198 57922 53266 57978
rect 53322 57922 53392 57978
rect 53072 57888 53392 57922
rect 83792 58350 84112 58384
rect 83792 58294 83862 58350
rect 83918 58294 83986 58350
rect 84042 58294 84112 58350
rect 83792 58226 84112 58294
rect 83792 58170 83862 58226
rect 83918 58170 83986 58226
rect 84042 58170 84112 58226
rect 83792 58102 84112 58170
rect 83792 58046 83862 58102
rect 83918 58046 83986 58102
rect 84042 58046 84112 58102
rect 83792 57978 84112 58046
rect 83792 57922 83862 57978
rect 83918 57922 83986 57978
rect 84042 57922 84112 57978
rect 83792 57888 84112 57922
rect 114512 58350 114832 58384
rect 114512 58294 114582 58350
rect 114638 58294 114706 58350
rect 114762 58294 114832 58350
rect 114512 58226 114832 58294
rect 114512 58170 114582 58226
rect 114638 58170 114706 58226
rect 114762 58170 114832 58226
rect 114512 58102 114832 58170
rect 114512 58046 114582 58102
rect 114638 58046 114706 58102
rect 114762 58046 114832 58102
rect 114512 57978 114832 58046
rect 114512 57922 114582 57978
rect 114638 57922 114706 57978
rect 114762 57922 114832 57978
rect 114512 57888 114832 57922
rect 145232 58350 145552 58384
rect 145232 58294 145302 58350
rect 145358 58294 145426 58350
rect 145482 58294 145552 58350
rect 145232 58226 145552 58294
rect 145232 58170 145302 58226
rect 145358 58170 145426 58226
rect 145482 58170 145552 58226
rect 145232 58102 145552 58170
rect 145232 58046 145302 58102
rect 145358 58046 145426 58102
rect 145482 58046 145552 58102
rect 145232 57978 145552 58046
rect 145232 57922 145302 57978
rect 145358 57922 145426 57978
rect 145482 57922 145552 57978
rect 145232 57888 145552 57922
rect 37712 46350 38032 46384
rect 37712 46294 37782 46350
rect 37838 46294 37906 46350
rect 37962 46294 38032 46350
rect 37712 46226 38032 46294
rect 37712 46170 37782 46226
rect 37838 46170 37906 46226
rect 37962 46170 38032 46226
rect 37712 46102 38032 46170
rect 37712 46046 37782 46102
rect 37838 46046 37906 46102
rect 37962 46046 38032 46102
rect 37712 45978 38032 46046
rect 37712 45922 37782 45978
rect 37838 45922 37906 45978
rect 37962 45922 38032 45978
rect 37712 45888 38032 45922
rect 68432 46350 68752 46384
rect 68432 46294 68502 46350
rect 68558 46294 68626 46350
rect 68682 46294 68752 46350
rect 68432 46226 68752 46294
rect 68432 46170 68502 46226
rect 68558 46170 68626 46226
rect 68682 46170 68752 46226
rect 68432 46102 68752 46170
rect 68432 46046 68502 46102
rect 68558 46046 68626 46102
rect 68682 46046 68752 46102
rect 68432 45978 68752 46046
rect 68432 45922 68502 45978
rect 68558 45922 68626 45978
rect 68682 45922 68752 45978
rect 68432 45888 68752 45922
rect 99152 46350 99472 46384
rect 99152 46294 99222 46350
rect 99278 46294 99346 46350
rect 99402 46294 99472 46350
rect 99152 46226 99472 46294
rect 99152 46170 99222 46226
rect 99278 46170 99346 46226
rect 99402 46170 99472 46226
rect 99152 46102 99472 46170
rect 99152 46046 99222 46102
rect 99278 46046 99346 46102
rect 99402 46046 99472 46102
rect 99152 45978 99472 46046
rect 99152 45922 99222 45978
rect 99278 45922 99346 45978
rect 99402 45922 99472 45978
rect 99152 45888 99472 45922
rect 129872 46350 130192 46384
rect 129872 46294 129942 46350
rect 129998 46294 130066 46350
rect 130122 46294 130192 46350
rect 129872 46226 130192 46294
rect 129872 46170 129942 46226
rect 129998 46170 130066 46226
rect 130122 46170 130192 46226
rect 129872 46102 130192 46170
rect 129872 46046 129942 46102
rect 129998 46046 130066 46102
rect 130122 46046 130192 46102
rect 129872 45978 130192 46046
rect 129872 45922 129942 45978
rect 129998 45922 130066 45978
rect 130122 45922 130192 45978
rect 129872 45888 130192 45922
rect 150332 43652 150388 371420
rect 150556 371364 150612 371374
rect 150556 44548 150612 371308
rect 150780 47236 150836 372204
rect 150892 353668 150948 353678
rect 150892 254212 150948 353612
rect 150892 254146 150948 254156
rect 151004 341908 151060 341918
rect 151004 182532 151060 341852
rect 151004 182466 151060 182476
rect 151116 325780 151172 325790
rect 151116 112644 151172 325724
rect 151116 112578 151172 112588
rect 152012 53620 152068 394268
rect 442652 394324 442708 394334
rect 162092 394212 162148 394222
rect 152012 53554 152068 53564
rect 152124 384020 152180 384030
rect 152124 51716 152180 383964
rect 159018 382350 159638 393242
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 152124 51650 152180 51660
rect 152236 375508 152292 375518
rect 152236 47908 152292 375452
rect 153804 374836 153860 374846
rect 153692 372820 153748 372830
rect 153692 347396 153748 372764
rect 153804 358148 153860 374780
rect 157164 371476 157220 371486
rect 155036 369460 155092 369470
rect 153804 358082 153860 358092
rect 153916 364756 153972 364766
rect 153692 347330 153748 347340
rect 152348 340340 152404 340350
rect 152348 229124 152404 340284
rect 153804 326452 153860 326462
rect 152348 229058 152404 229068
rect 153692 323764 153748 323774
rect 152908 112644 152964 112654
rect 152908 96516 152964 112588
rect 152908 96450 152964 96460
rect 153692 85764 153748 323708
rect 153804 100100 153860 326396
rect 153916 304388 153972 364700
rect 154364 362852 154420 362862
rect 154364 354564 154420 362796
rect 154364 354498 154420 354508
rect 154476 357924 154532 357934
rect 154476 350980 154532 357868
rect 154476 350914 154532 350924
rect 154364 348628 154420 348638
rect 154252 343252 154308 343262
rect 154140 337876 154196 337886
rect 153916 304322 153972 304332
rect 154028 332500 154084 332510
rect 153804 100034 153860 100044
rect 153916 265524 153972 265534
rect 153692 85698 153748 85708
rect 153804 96628 153860 96638
rect 153804 78596 153860 96572
rect 153804 78530 153860 78540
rect 152236 47842 152292 47852
rect 153692 75348 153748 75358
rect 150780 47170 150836 47180
rect 150556 44482 150612 44492
rect 150332 43586 150388 43596
rect 152012 41860 152068 41870
rect 22352 40350 22672 40384
rect 22352 40294 22422 40350
rect 22478 40294 22546 40350
rect 22602 40294 22672 40350
rect 22352 40226 22672 40294
rect 22352 40170 22422 40226
rect 22478 40170 22546 40226
rect 22602 40170 22672 40226
rect 22352 40102 22672 40170
rect 22352 40046 22422 40102
rect 22478 40046 22546 40102
rect 22602 40046 22672 40102
rect 22352 39978 22672 40046
rect 22352 39922 22422 39978
rect 22478 39922 22546 39978
rect 22602 39922 22672 39978
rect 22352 39888 22672 39922
rect 53072 40350 53392 40384
rect 53072 40294 53142 40350
rect 53198 40294 53266 40350
rect 53322 40294 53392 40350
rect 53072 40226 53392 40294
rect 53072 40170 53142 40226
rect 53198 40170 53266 40226
rect 53322 40170 53392 40226
rect 53072 40102 53392 40170
rect 53072 40046 53142 40102
rect 53198 40046 53266 40102
rect 53322 40046 53392 40102
rect 53072 39978 53392 40046
rect 53072 39922 53142 39978
rect 53198 39922 53266 39978
rect 53322 39922 53392 39978
rect 53072 39888 53392 39922
rect 83792 40350 84112 40384
rect 83792 40294 83862 40350
rect 83918 40294 83986 40350
rect 84042 40294 84112 40350
rect 83792 40226 84112 40294
rect 83792 40170 83862 40226
rect 83918 40170 83986 40226
rect 84042 40170 84112 40226
rect 83792 40102 84112 40170
rect 83792 40046 83862 40102
rect 83918 40046 83986 40102
rect 84042 40046 84112 40102
rect 83792 39978 84112 40046
rect 83792 39922 83862 39978
rect 83918 39922 83986 39978
rect 84042 39922 84112 39978
rect 83792 39888 84112 39922
rect 114512 40350 114832 40384
rect 114512 40294 114582 40350
rect 114638 40294 114706 40350
rect 114762 40294 114832 40350
rect 114512 40226 114832 40294
rect 114512 40170 114582 40226
rect 114638 40170 114706 40226
rect 114762 40170 114832 40226
rect 114512 40102 114832 40170
rect 114512 40046 114582 40102
rect 114638 40046 114706 40102
rect 114762 40046 114832 40102
rect 114512 39978 114832 40046
rect 114512 39922 114582 39978
rect 114638 39922 114706 39978
rect 114762 39922 114832 39978
rect 114512 39888 114832 39922
rect 145232 40350 145552 40384
rect 145232 40294 145302 40350
rect 145358 40294 145426 40350
rect 145482 40294 145552 40350
rect 145232 40226 145552 40294
rect 145232 40170 145302 40226
rect 145358 40170 145426 40226
rect 145482 40170 145552 40226
rect 145232 40102 145552 40170
rect 145232 40046 145302 40102
rect 145358 40046 145426 40102
rect 145482 40046 145552 40102
rect 145232 39978 145552 40046
rect 145232 39922 145302 39978
rect 145358 39922 145426 39978
rect 145482 39922 145552 39978
rect 145232 39888 145552 39922
rect 150332 36484 150388 36494
rect 37712 28350 38032 28384
rect 37712 28294 37782 28350
rect 37838 28294 37906 28350
rect 37962 28294 38032 28350
rect 37712 28226 38032 28294
rect 37712 28170 37782 28226
rect 37838 28170 37906 28226
rect 37962 28170 38032 28226
rect 37712 28102 38032 28170
rect 37712 28046 37782 28102
rect 37838 28046 37906 28102
rect 37962 28046 38032 28102
rect 37712 27978 38032 28046
rect 37712 27922 37782 27978
rect 37838 27922 37906 27978
rect 37962 27922 38032 27978
rect 37712 27888 38032 27922
rect 68432 28350 68752 28384
rect 68432 28294 68502 28350
rect 68558 28294 68626 28350
rect 68682 28294 68752 28350
rect 68432 28226 68752 28294
rect 68432 28170 68502 28226
rect 68558 28170 68626 28226
rect 68682 28170 68752 28226
rect 68432 28102 68752 28170
rect 68432 28046 68502 28102
rect 68558 28046 68626 28102
rect 68682 28046 68752 28102
rect 68432 27978 68752 28046
rect 68432 27922 68502 27978
rect 68558 27922 68626 27978
rect 68682 27922 68752 27978
rect 68432 27888 68752 27922
rect 99152 28350 99472 28384
rect 99152 28294 99222 28350
rect 99278 28294 99346 28350
rect 99402 28294 99472 28350
rect 99152 28226 99472 28294
rect 99152 28170 99222 28226
rect 99278 28170 99346 28226
rect 99402 28170 99472 28226
rect 99152 28102 99472 28170
rect 99152 28046 99222 28102
rect 99278 28046 99346 28102
rect 99402 28046 99472 28102
rect 99152 27978 99472 28046
rect 99152 27922 99222 27978
rect 99278 27922 99346 27978
rect 99402 27922 99472 27978
rect 99152 27888 99472 27922
rect 129872 28350 130192 28384
rect 129872 28294 129942 28350
rect 129998 28294 130066 28350
rect 130122 28294 130192 28350
rect 129872 28226 130192 28294
rect 129872 28170 129942 28226
rect 129998 28170 130066 28226
rect 130122 28170 130192 28226
rect 129872 28102 130192 28170
rect 129872 28046 129942 28102
rect 129998 28046 130066 28102
rect 130122 28046 130192 28102
rect 129872 27978 130192 28046
rect 129872 27922 129942 27978
rect 129998 27922 130066 27978
rect 130122 27922 130192 27978
rect 129872 27888 130192 27922
rect 149772 22148 149828 22158
rect 9884 18050 9940 18060
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 23436 13618 23492 13628
rect 17276 9298 17332 9308
rect 11564 5878 11620 5888
rect 11564 3444 11620 5822
rect 17276 4228 17332 9242
rect 23436 4340 23492 13562
rect 23436 4274 23492 4284
rect 26796 6058 26852 6068
rect 17276 4162 17332 4172
rect 11564 3378 11620 3388
rect 13356 3444 13412 3454
rect 13356 3358 13412 3388
rect 26796 3444 26852 6002
rect 26796 3378 26852 3388
rect 36138 4350 36758 19026
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 13356 3292 13412 3302
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 10350 40478 19026
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 44492 11818 44548 11828
rect 44492 7588 44548 11762
rect 44492 7522 44548 7532
rect 55356 7678 55412 7688
rect 41804 7498 41860 7508
rect 41804 3780 41860 7442
rect 55356 3892 55412 7622
rect 55356 3826 55412 3836
rect 66858 4350 67478 19026
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 41804 3714 41860 3724
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 10350 71198 19026
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 4350 98198 19026
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 10350 101918 19026
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 4350 128918 19026
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 10350 132638 19026
rect 149772 14420 149828 22092
rect 150332 19236 150388 36428
rect 150332 19170 150388 19180
rect 150444 25732 150500 25742
rect 150444 16436 150500 25676
rect 152012 16678 152068 41804
rect 153692 35588 153748 75292
rect 153916 64260 153972 265468
rect 154028 132356 154084 332444
rect 154140 161028 154196 337820
rect 154252 189700 154308 343196
rect 154364 218372 154420 348572
rect 155036 329476 155092 369404
rect 155596 368788 155652 368798
rect 155372 368116 155428 368126
rect 155036 329410 155092 329420
rect 155148 366772 155204 366782
rect 155148 315140 155204 366716
rect 155372 322308 155428 368060
rect 155596 325892 155652 368732
rect 156828 367444 156884 367454
rect 156156 354004 156212 354014
rect 156044 343924 156100 343934
rect 155932 341236 155988 341246
rect 155820 338548 155876 338558
rect 155596 325826 155652 325836
rect 155708 330148 155764 330158
rect 155372 322242 155428 322252
rect 155148 315074 155204 315084
rect 155484 320068 155540 320078
rect 155372 315028 155428 315038
rect 154476 304948 154532 304958
rect 154476 261380 154532 304892
rect 154476 261314 154532 261324
rect 154364 218306 154420 218316
rect 154252 189634 154308 189644
rect 154140 160962 154196 160972
rect 154364 160468 154420 160478
rect 154028 132290 154084 132300
rect 154140 158004 154196 158014
rect 153916 64194 153972 64204
rect 154028 74788 154084 74798
rect 154028 53508 154084 74732
rect 154140 57092 154196 157948
rect 154364 146692 154420 160412
rect 154364 146626 154420 146636
rect 154252 132468 154308 132478
rect 154252 128772 154308 132412
rect 154252 128706 154308 128716
rect 154476 123508 154532 123518
rect 154476 118020 154532 123452
rect 154476 117954 154532 117964
rect 154476 91588 154532 91598
rect 154476 89348 154532 91532
rect 154476 89282 154532 89292
rect 154252 84868 154308 84878
rect 154252 71428 154308 84812
rect 154252 71362 154308 71372
rect 154140 57026 154196 57036
rect 154028 53442 154084 53452
rect 155372 49924 155428 314972
rect 155484 135940 155540 320012
rect 155484 135874 155540 135884
rect 155596 315140 155652 315150
rect 155372 49858 155428 49868
rect 155484 89908 155540 89918
rect 155484 39172 155540 89852
rect 155596 75012 155652 315084
rect 155708 150276 155764 330092
rect 155820 164612 155876 338492
rect 155932 178948 155988 341180
rect 156044 193284 156100 343868
rect 156156 247044 156212 353948
rect 156828 318724 156884 367388
rect 157052 367108 157108 367118
rect 156828 318658 156884 318668
rect 156940 360388 156996 360398
rect 156940 307972 156996 360332
rect 157052 333060 157108 367052
rect 157164 340228 157220 371420
rect 157836 366100 157892 366110
rect 157164 340162 157220 340172
rect 157724 358708 157780 358718
rect 157612 339220 157668 339230
rect 157500 336532 157556 336542
rect 157052 332994 157108 333004
rect 157388 333844 157444 333854
rect 157276 331156 157332 331166
rect 157164 325332 157220 325342
rect 156940 307906 156996 307916
rect 157052 318500 157108 318510
rect 156156 246978 156212 246988
rect 156044 193218 156100 193228
rect 155932 178882 155988 178892
rect 155820 164546 155876 164556
rect 155708 150210 155764 150220
rect 156044 163828 156100 163838
rect 155596 74946 155652 74956
rect 156044 42756 156100 163772
rect 157052 92932 157108 318444
rect 157164 110852 157220 325276
rect 157276 125188 157332 331100
rect 157388 139524 157444 333788
rect 157500 153860 157556 336476
rect 157612 168196 157668 339164
rect 157724 272132 157780 358652
rect 157836 311556 157892 366044
rect 159018 364350 159638 381922
rect 160748 374164 160804 374174
rect 160524 373492 160580 373502
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 157836 311490 157892 311500
rect 158508 356020 158564 356030
rect 157724 272066 157780 272076
rect 158508 257796 158564 355964
rect 158508 257730 158564 257740
rect 158620 353332 158676 353342
rect 158620 243460 158676 353276
rect 159018 346350 159638 363922
rect 160412 370804 160468 370814
rect 159018 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 159638 346350
rect 159018 346226 159638 346294
rect 159018 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 159638 346226
rect 159018 346102 159638 346170
rect 159018 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 159638 346102
rect 159018 345978 159638 346046
rect 159018 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 159638 345978
rect 158844 331828 158900 331838
rect 158620 243394 158676 243404
rect 158732 322420 158788 322430
rect 157612 168130 157668 168140
rect 157500 153794 157556 153804
rect 157388 139458 157444 139468
rect 157276 125122 157332 125132
rect 157500 125188 157556 125198
rect 157164 110786 157220 110796
rect 157052 92866 157108 92876
rect 157500 46340 157556 125132
rect 158732 96628 158788 322364
rect 158844 132468 158900 331772
rect 158844 132402 158900 132412
rect 159018 328350 159638 345922
rect 159018 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 159638 328350
rect 159018 328226 159638 328294
rect 159018 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 159638 328226
rect 159018 328102 159638 328170
rect 159018 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 159638 328102
rect 159018 327978 159638 328046
rect 159018 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 159638 327978
rect 159018 310350 159638 327922
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 159018 292350 159638 309922
rect 160300 362180 160356 362190
rect 160300 300804 160356 362124
rect 160412 336644 160468 370748
rect 160524 357924 160580 373436
rect 160748 362852 160804 374108
rect 160748 362786 160804 362796
rect 160524 357858 160580 357868
rect 161196 361396 161252 361406
rect 161084 345268 161140 345278
rect 160412 336578 160468 336588
rect 160860 339892 160916 339902
rect 160748 334516 160804 334526
rect 160636 329140 160692 329150
rect 160300 300738 160356 300748
rect 160412 323092 160468 323102
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 159018 274350 159638 291922
rect 159018 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 159638 274350
rect 159018 274226 159638 274294
rect 159018 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 159638 274226
rect 159018 274102 159638 274170
rect 159018 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 159638 274102
rect 159018 273978 159638 274046
rect 159018 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 159638 273978
rect 159018 256350 159638 273922
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 159018 202350 159638 219922
rect 159018 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 159638 202350
rect 159018 202226 159638 202294
rect 159018 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 159638 202226
rect 159018 202102 159638 202170
rect 159018 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 159638 202102
rect 159018 201978 159638 202046
rect 159018 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 159638 201978
rect 159018 184350 159638 201922
rect 159018 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 159638 184350
rect 159018 184226 159638 184294
rect 159018 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 159638 184226
rect 159018 184102 159638 184170
rect 159018 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 159638 184102
rect 159018 183978 159638 184046
rect 159018 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 159638 183978
rect 159018 166350 159638 183922
rect 159018 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 159638 166350
rect 159018 166226 159638 166294
rect 159018 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 159638 166226
rect 159018 166102 159638 166170
rect 159018 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 159638 166102
rect 159018 165978 159638 166046
rect 159018 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 159638 165978
rect 159018 148350 159638 165922
rect 159018 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 159638 148350
rect 159018 148226 159638 148294
rect 159018 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 159638 148226
rect 159018 148102 159638 148170
rect 159018 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 159638 148102
rect 159018 147978 159638 148046
rect 159018 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 159638 147978
rect 158732 96562 158788 96572
rect 159018 130350 159638 147922
rect 159018 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 159638 130350
rect 159018 130226 159638 130294
rect 159018 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 159638 130226
rect 159018 130102 159638 130170
rect 159018 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 159638 130102
rect 159018 129978 159638 130046
rect 159018 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 159638 129978
rect 159018 112350 159638 129922
rect 159018 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 159638 112350
rect 159018 112226 159638 112294
rect 159018 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 159638 112226
rect 159018 112102 159638 112170
rect 159018 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 159638 112102
rect 159018 111978 159638 112046
rect 159018 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 159638 111978
rect 157500 46274 157556 46284
rect 159018 94350 159638 111922
rect 159018 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 159638 94350
rect 159018 94226 159638 94294
rect 159018 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 159638 94226
rect 159018 94102 159638 94170
rect 159018 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 159638 94102
rect 159018 93978 159638 94046
rect 159018 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 159638 93978
rect 159018 76350 159638 93922
rect 160412 82180 160468 323036
rect 160412 82114 160468 82124
rect 160524 303268 160580 303278
rect 159018 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 159638 76350
rect 159018 76226 159638 76294
rect 159018 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 159638 76226
rect 159018 76102 159638 76170
rect 159018 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 159638 76102
rect 159018 75978 159638 76046
rect 159018 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 159638 75978
rect 159018 58350 159638 75922
rect 160524 60676 160580 303212
rect 160636 114436 160692 329084
rect 160748 143108 160804 334460
rect 160860 171780 160916 339836
rect 160860 171714 160916 171724
rect 160972 318388 161028 318398
rect 160972 158004 161028 318332
rect 161084 200452 161140 345212
rect 161196 286468 161252 361340
rect 161196 286402 161252 286412
rect 161980 319732 162036 319742
rect 161980 265524 162036 319676
rect 161980 265458 162036 265468
rect 161084 200386 161140 200396
rect 160972 157938 161028 157948
rect 160748 143042 160804 143052
rect 160636 114370 160692 114380
rect 160524 60610 160580 60620
rect 159018 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 159638 58350
rect 159018 58226 159638 58294
rect 159018 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 159638 58226
rect 159018 58102 159638 58170
rect 159018 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 159638 58102
rect 159018 57978 159638 58046
rect 159018 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 159638 57978
rect 156044 42690 156100 42700
rect 155484 39106 155540 39116
rect 159018 40350 159638 57922
rect 162092 49028 162148 394156
rect 437612 394212 437668 394222
rect 162316 394100 162372 394110
rect 162204 390740 162260 390750
rect 162204 50820 162260 390684
rect 162316 56196 162372 394044
rect 427532 394100 427588 394110
rect 166012 393988 166068 393998
rect 162738 388350 163358 393242
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 165900 390628 165956 390638
rect 165788 383908 165844 383918
rect 163996 377300 164052 377310
rect 163884 373828 163940 373838
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162738 352350 163358 369922
rect 162738 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163358 352350
rect 162738 352226 163358 352294
rect 162738 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163358 352226
rect 162738 352102 163358 352170
rect 162738 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163358 352102
rect 162738 351978 163358 352046
rect 162738 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163358 351978
rect 162540 351092 162596 351102
rect 162428 327124 162484 327134
rect 162428 103684 162484 327068
rect 162540 232708 162596 351036
rect 162540 232642 162596 232652
rect 162738 334350 163358 351922
rect 162738 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 163358 334350
rect 162738 334226 163358 334294
rect 162738 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 163358 334226
rect 162738 334102 163358 334170
rect 162738 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 163358 334102
rect 162738 333978 163358 334046
rect 162738 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 163358 333978
rect 162738 316350 163358 333922
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 162738 298350 163358 315922
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 162738 280350 163358 297922
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 162738 262350 163358 279922
rect 162738 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 163358 262350
rect 162738 262226 163358 262294
rect 162738 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 163358 262226
rect 162738 262102 163358 262170
rect 162738 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 163358 262102
rect 162738 261978 163358 262046
rect 162738 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 163358 261978
rect 162738 244350 163358 261922
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162428 103618 162484 103628
rect 162738 226350 163358 243922
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 162738 208350 163358 225922
rect 162738 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163358 208350
rect 162738 208226 163358 208294
rect 162738 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163358 208226
rect 162738 208102 163358 208170
rect 162738 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163358 208102
rect 162738 207978 163358 208046
rect 162738 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163358 207978
rect 162738 190350 163358 207922
rect 162738 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 163358 190350
rect 162738 190226 163358 190294
rect 162738 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 163358 190226
rect 162738 190102 163358 190170
rect 162738 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 163358 190102
rect 162738 189978 163358 190046
rect 162738 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 163358 189978
rect 162738 172350 163358 189922
rect 162738 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 163358 172350
rect 162738 172226 163358 172294
rect 162738 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 163358 172226
rect 162738 172102 163358 172170
rect 162738 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 163358 172102
rect 162738 171978 163358 172046
rect 162738 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 163358 171978
rect 162738 154350 163358 171922
rect 162738 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 163358 154350
rect 162738 154226 163358 154294
rect 162738 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 163358 154226
rect 162738 154102 163358 154170
rect 162738 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 163358 154102
rect 162738 153978 163358 154046
rect 162738 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 163358 153978
rect 162738 136350 163358 153922
rect 162738 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 163358 136350
rect 162738 136226 163358 136294
rect 162738 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 163358 136226
rect 162738 136102 163358 136170
rect 162738 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 163358 136102
rect 162738 135978 163358 136046
rect 162738 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 163358 135978
rect 162738 118350 163358 135922
rect 162738 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 163358 118350
rect 162738 118226 163358 118294
rect 162738 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 163358 118226
rect 162738 118102 163358 118170
rect 162738 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 163358 118102
rect 162738 117978 163358 118046
rect 162738 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 163358 117978
rect 162316 56130 162372 56140
rect 162738 100350 163358 117922
rect 162738 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 163358 100350
rect 162738 100226 163358 100294
rect 162738 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 163358 100226
rect 162738 100102 163358 100170
rect 162738 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 163358 100102
rect 162738 99978 163358 100046
rect 162738 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 163358 99978
rect 162738 82350 163358 99922
rect 162738 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 163358 82350
rect 162738 82226 163358 82294
rect 162738 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 163358 82226
rect 162738 82102 163358 82170
rect 162738 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 163358 82102
rect 162738 81978 163358 82046
rect 162738 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 163358 81978
rect 162738 64350 163358 81922
rect 162738 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 163358 64350
rect 162738 64226 163358 64294
rect 162738 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 163358 64226
rect 162738 64102 163358 64170
rect 162738 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 163358 64102
rect 162738 63978 163358 64046
rect 162738 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 163358 63978
rect 162204 50754 162260 50764
rect 162092 48962 162148 48972
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 153692 35522 153748 35532
rect 155372 38276 155428 38286
rect 152236 32900 152292 32910
rect 152012 16612 152068 16622
rect 152124 31108 152180 31118
rect 152124 16548 152180 31052
rect 152236 17780 152292 32844
rect 153692 30212 153748 30222
rect 152348 23940 152404 23950
rect 152348 19348 152404 23884
rect 152348 19282 152404 19292
rect 153692 18004 153748 30156
rect 153692 17938 153748 17948
rect 153916 24836 153972 24846
rect 153916 17892 153972 24780
rect 155372 21028 155428 38220
rect 155372 20962 155428 20972
rect 159018 22350 159638 39922
rect 162738 46350 163358 63922
rect 163772 372148 163828 372158
rect 163772 49924 163828 372092
rect 163884 55300 163940 373772
rect 163996 57988 164052 377244
rect 165452 375508 165508 375518
rect 165452 361732 165508 375452
rect 165452 361666 165508 361676
rect 165676 347956 165732 347966
rect 165564 340564 165620 340574
rect 164220 334404 164276 334414
rect 164108 329252 164164 329262
rect 164108 186116 164164 329196
rect 164220 297220 164276 334348
rect 164220 297154 164276 297164
rect 165452 320404 165508 320414
rect 164108 186050 164164 186060
rect 163996 57922 164052 57932
rect 164556 74004 164612 74014
rect 163884 55234 163940 55244
rect 163772 49858 163828 49868
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 163660 47908 163716 47918
rect 163660 45444 163716 47852
rect 164556 46340 164612 73948
rect 165452 67956 165508 320348
rect 165564 175364 165620 340508
rect 165676 214788 165732 347900
rect 165676 214722 165732 214732
rect 165564 175298 165620 175308
rect 165452 67890 165508 67900
rect 165788 52612 165844 383852
rect 165900 55468 165956 390572
rect 166012 67228 166068 393932
rect 169708 389620 169764 389630
rect 168812 372148 168868 372158
rect 167468 362068 167524 362078
rect 166124 359380 166180 359390
rect 166124 275716 166180 359324
rect 167356 335188 167412 335198
rect 167244 330484 167300 330494
rect 166124 275650 166180 275660
rect 167132 317716 167188 317726
rect 167132 74788 167188 317660
rect 167244 121604 167300 330428
rect 167356 160468 167412 335132
rect 167468 290052 167524 362012
rect 167468 289986 167524 289996
rect 167580 355124 167636 355134
rect 167580 282884 167636 355068
rect 168812 343812 168868 372092
rect 169260 360052 169316 360062
rect 169148 349972 169204 349982
rect 168812 343746 168868 343756
rect 169036 349300 169092 349310
rect 168924 329812 168980 329822
rect 168812 317044 168868 317054
rect 167580 282818 167636 282828
rect 167692 289044 167748 289054
rect 167692 264964 167748 288988
rect 167692 264898 167748 264908
rect 167356 160402 167412 160412
rect 167244 121538 167300 121548
rect 168812 75348 168868 316988
rect 168924 123508 168980 329756
rect 169036 221956 169092 349244
rect 169148 225540 169204 349916
rect 169260 279300 169316 359996
rect 169372 356692 169428 356702
rect 169372 304948 169428 356636
rect 169372 304882 169428 304892
rect 169260 279234 169316 279244
rect 169148 225474 169204 225484
rect 169036 221890 169092 221900
rect 168924 123442 168980 123452
rect 168812 75282 168868 75292
rect 169596 76468 169652 76478
rect 167132 74722 167188 74732
rect 166012 67172 166292 67228
rect 165900 55412 166068 55468
rect 166012 54404 166068 55412
rect 166012 54338 166068 54348
rect 165788 52546 165844 52556
rect 166236 48132 166292 67172
rect 166236 48066 166292 48076
rect 164556 46274 164612 46284
rect 163660 45378 163716 45388
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 153916 17826 153972 17836
rect 152236 17714 152292 17724
rect 152124 16482 152180 16492
rect 150444 16370 150500 16380
rect 149772 14354 149828 14364
rect 134428 11998 134484 12008
rect 134428 11284 134484 11942
rect 134428 11218 134484 11228
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 4350 159638 21922
rect 159740 23044 159796 23054
rect 159740 18340 159796 22988
rect 159740 18274 159796 18284
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 10350 163358 27922
rect 163548 34692 163604 34702
rect 163548 19796 163604 34636
rect 163548 19730 163604 19740
rect 163772 33796 163828 33806
rect 163772 18452 163828 33740
rect 163884 32004 163940 32014
rect 163884 19460 163940 31948
rect 164108 29316 164164 29326
rect 163884 19394 163940 19404
rect 163996 28420 164052 28430
rect 163772 18386 163828 18396
rect 163996 16660 164052 28364
rect 164108 19908 164164 29260
rect 164108 19842 164164 19852
rect 164220 27524 164276 27534
rect 164220 18228 164276 27468
rect 164332 26628 164388 26638
rect 164332 19572 164388 26572
rect 164332 19506 164388 19516
rect 164220 18162 164276 18172
rect 164556 18564 164612 18574
rect 163996 16594 164052 16604
rect 164556 16324 164612 18508
rect 164556 16258 164612 16268
rect 169596 13438 169652 76412
rect 169708 74004 169764 389564
rect 425852 378868 425908 378878
rect 424172 377188 424228 377198
rect 420924 374836 420980 374846
rect 417564 373492 417620 373502
rect 193808 370350 194128 370384
rect 193808 370294 193878 370350
rect 193934 370294 194002 370350
rect 194058 370294 194128 370350
rect 193808 370226 194128 370294
rect 193808 370170 193878 370226
rect 193934 370170 194002 370226
rect 194058 370170 194128 370226
rect 169820 370132 169876 370142
rect 169820 367108 169876 370076
rect 193808 370102 194128 370170
rect 193808 370046 193878 370102
rect 193934 370046 194002 370102
rect 194058 370046 194128 370102
rect 193808 369978 194128 370046
rect 193808 369922 193878 369978
rect 193934 369922 194002 369978
rect 194058 369922 194128 369978
rect 193808 369888 194128 369922
rect 224528 370350 224848 370384
rect 224528 370294 224598 370350
rect 224654 370294 224722 370350
rect 224778 370294 224848 370350
rect 224528 370226 224848 370294
rect 224528 370170 224598 370226
rect 224654 370170 224722 370226
rect 224778 370170 224848 370226
rect 224528 370102 224848 370170
rect 224528 370046 224598 370102
rect 224654 370046 224722 370102
rect 224778 370046 224848 370102
rect 224528 369978 224848 370046
rect 224528 369922 224598 369978
rect 224654 369922 224722 369978
rect 224778 369922 224848 369978
rect 224528 369888 224848 369922
rect 255248 370350 255568 370384
rect 255248 370294 255318 370350
rect 255374 370294 255442 370350
rect 255498 370294 255568 370350
rect 255248 370226 255568 370294
rect 255248 370170 255318 370226
rect 255374 370170 255442 370226
rect 255498 370170 255568 370226
rect 255248 370102 255568 370170
rect 255248 370046 255318 370102
rect 255374 370046 255442 370102
rect 255498 370046 255568 370102
rect 255248 369978 255568 370046
rect 255248 369922 255318 369978
rect 255374 369922 255442 369978
rect 255498 369922 255568 369978
rect 255248 369888 255568 369922
rect 285968 370350 286288 370384
rect 285968 370294 286038 370350
rect 286094 370294 286162 370350
rect 286218 370294 286288 370350
rect 285968 370226 286288 370294
rect 285968 370170 286038 370226
rect 286094 370170 286162 370226
rect 286218 370170 286288 370226
rect 285968 370102 286288 370170
rect 285968 370046 286038 370102
rect 286094 370046 286162 370102
rect 286218 370046 286288 370102
rect 285968 369978 286288 370046
rect 285968 369922 286038 369978
rect 286094 369922 286162 369978
rect 286218 369922 286288 369978
rect 285968 369888 286288 369922
rect 316688 370350 317008 370384
rect 316688 370294 316758 370350
rect 316814 370294 316882 370350
rect 316938 370294 317008 370350
rect 316688 370226 317008 370294
rect 316688 370170 316758 370226
rect 316814 370170 316882 370226
rect 316938 370170 317008 370226
rect 316688 370102 317008 370170
rect 316688 370046 316758 370102
rect 316814 370046 316882 370102
rect 316938 370046 317008 370102
rect 316688 369978 317008 370046
rect 316688 369922 316758 369978
rect 316814 369922 316882 369978
rect 316938 369922 317008 369978
rect 316688 369888 317008 369922
rect 347408 370350 347728 370384
rect 347408 370294 347478 370350
rect 347534 370294 347602 370350
rect 347658 370294 347728 370350
rect 347408 370226 347728 370294
rect 347408 370170 347478 370226
rect 347534 370170 347602 370226
rect 347658 370170 347728 370226
rect 347408 370102 347728 370170
rect 347408 370046 347478 370102
rect 347534 370046 347602 370102
rect 347658 370046 347728 370102
rect 347408 369978 347728 370046
rect 347408 369922 347478 369978
rect 347534 369922 347602 369978
rect 347658 369922 347728 369978
rect 347408 369888 347728 369922
rect 378128 370350 378448 370384
rect 378128 370294 378198 370350
rect 378254 370294 378322 370350
rect 378378 370294 378448 370350
rect 378128 370226 378448 370294
rect 378128 370170 378198 370226
rect 378254 370170 378322 370226
rect 378378 370170 378448 370226
rect 378128 370102 378448 370170
rect 378128 370046 378198 370102
rect 378254 370046 378322 370102
rect 378378 370046 378448 370102
rect 378128 369978 378448 370046
rect 378128 369922 378198 369978
rect 378254 369922 378322 369978
rect 378378 369922 378448 369978
rect 378128 369888 378448 369922
rect 408848 370350 409168 370384
rect 408848 370294 408918 370350
rect 408974 370294 409042 370350
rect 409098 370294 409168 370350
rect 408848 370226 409168 370294
rect 408848 370170 408918 370226
rect 408974 370170 409042 370226
rect 409098 370170 409168 370226
rect 408848 370102 409168 370170
rect 408848 370046 408918 370102
rect 408974 370046 409042 370102
rect 409098 370046 409168 370102
rect 408848 369978 409168 370046
rect 408848 369922 408918 369978
rect 408974 369922 409042 369978
rect 409098 369922 409168 369978
rect 408848 369888 409168 369922
rect 169820 367042 169876 367052
rect 170828 365428 170884 365438
rect 169820 364084 169876 364094
rect 169820 362180 169876 364028
rect 169820 362114 169876 362124
rect 170492 363412 170548 363422
rect 170268 360724 170324 360734
rect 169820 355348 169876 355358
rect 169820 353668 169876 355292
rect 170268 355124 170324 360668
rect 170268 355058 170324 355068
rect 169820 353602 169876 353612
rect 169820 335860 169876 335870
rect 169820 330148 169876 335804
rect 170492 334404 170548 363356
rect 170828 360388 170884 365372
rect 416108 364756 416164 364766
rect 178448 364350 178768 364384
rect 178448 364294 178518 364350
rect 178574 364294 178642 364350
rect 178698 364294 178768 364350
rect 178448 364226 178768 364294
rect 178448 364170 178518 364226
rect 178574 364170 178642 364226
rect 178698 364170 178768 364226
rect 178448 364102 178768 364170
rect 178448 364046 178518 364102
rect 178574 364046 178642 364102
rect 178698 364046 178768 364102
rect 178448 363978 178768 364046
rect 178448 363922 178518 363978
rect 178574 363922 178642 363978
rect 178698 363922 178768 363978
rect 178448 363888 178768 363922
rect 209168 364350 209488 364384
rect 209168 364294 209238 364350
rect 209294 364294 209362 364350
rect 209418 364294 209488 364350
rect 209168 364226 209488 364294
rect 209168 364170 209238 364226
rect 209294 364170 209362 364226
rect 209418 364170 209488 364226
rect 209168 364102 209488 364170
rect 209168 364046 209238 364102
rect 209294 364046 209362 364102
rect 209418 364046 209488 364102
rect 209168 363978 209488 364046
rect 209168 363922 209238 363978
rect 209294 363922 209362 363978
rect 209418 363922 209488 363978
rect 209168 363888 209488 363922
rect 239888 364350 240208 364384
rect 239888 364294 239958 364350
rect 240014 364294 240082 364350
rect 240138 364294 240208 364350
rect 239888 364226 240208 364294
rect 239888 364170 239958 364226
rect 240014 364170 240082 364226
rect 240138 364170 240208 364226
rect 239888 364102 240208 364170
rect 239888 364046 239958 364102
rect 240014 364046 240082 364102
rect 240138 364046 240208 364102
rect 239888 363978 240208 364046
rect 239888 363922 239958 363978
rect 240014 363922 240082 363978
rect 240138 363922 240208 363978
rect 239888 363888 240208 363922
rect 270608 364350 270928 364384
rect 270608 364294 270678 364350
rect 270734 364294 270802 364350
rect 270858 364294 270928 364350
rect 270608 364226 270928 364294
rect 270608 364170 270678 364226
rect 270734 364170 270802 364226
rect 270858 364170 270928 364226
rect 270608 364102 270928 364170
rect 270608 364046 270678 364102
rect 270734 364046 270802 364102
rect 270858 364046 270928 364102
rect 270608 363978 270928 364046
rect 270608 363922 270678 363978
rect 270734 363922 270802 363978
rect 270858 363922 270928 363978
rect 270608 363888 270928 363922
rect 301328 364350 301648 364384
rect 301328 364294 301398 364350
rect 301454 364294 301522 364350
rect 301578 364294 301648 364350
rect 301328 364226 301648 364294
rect 301328 364170 301398 364226
rect 301454 364170 301522 364226
rect 301578 364170 301648 364226
rect 301328 364102 301648 364170
rect 301328 364046 301398 364102
rect 301454 364046 301522 364102
rect 301578 364046 301648 364102
rect 301328 363978 301648 364046
rect 301328 363922 301398 363978
rect 301454 363922 301522 363978
rect 301578 363922 301648 363978
rect 301328 363888 301648 363922
rect 332048 364350 332368 364384
rect 332048 364294 332118 364350
rect 332174 364294 332242 364350
rect 332298 364294 332368 364350
rect 332048 364226 332368 364294
rect 332048 364170 332118 364226
rect 332174 364170 332242 364226
rect 332298 364170 332368 364226
rect 332048 364102 332368 364170
rect 332048 364046 332118 364102
rect 332174 364046 332242 364102
rect 332298 364046 332368 364102
rect 332048 363978 332368 364046
rect 332048 363922 332118 363978
rect 332174 363922 332242 363978
rect 332298 363922 332368 363978
rect 332048 363888 332368 363922
rect 362768 364350 363088 364384
rect 362768 364294 362838 364350
rect 362894 364294 362962 364350
rect 363018 364294 363088 364350
rect 362768 364226 363088 364294
rect 362768 364170 362838 364226
rect 362894 364170 362962 364226
rect 363018 364170 363088 364226
rect 362768 364102 363088 364170
rect 362768 364046 362838 364102
rect 362894 364046 362962 364102
rect 363018 364046 363088 364102
rect 362768 363978 363088 364046
rect 362768 363922 362838 363978
rect 362894 363922 362962 363978
rect 363018 363922 363088 363978
rect 362768 363888 363088 363922
rect 393488 364350 393808 364384
rect 393488 364294 393558 364350
rect 393614 364294 393682 364350
rect 393738 364294 393808 364350
rect 393488 364226 393808 364294
rect 393488 364170 393558 364226
rect 393614 364170 393682 364226
rect 393738 364170 393808 364226
rect 393488 364102 393808 364170
rect 393488 364046 393558 364102
rect 393614 364046 393682 364102
rect 393738 364046 393808 364102
rect 393488 363978 393808 364046
rect 393488 363922 393558 363978
rect 393614 363922 393682 363978
rect 393738 363922 393808 363978
rect 393488 363888 393808 363922
rect 170828 360322 170884 360332
rect 172620 362740 172676 362750
rect 171052 357364 171108 357374
rect 170828 351988 170884 351998
rect 170492 334338 170548 334348
rect 170604 345940 170660 345950
rect 169820 330082 169876 330092
rect 170492 333172 170548 333182
rect 169820 328468 169876 328478
rect 169820 325332 169876 328412
rect 169820 325266 169876 325276
rect 169820 325108 169876 325118
rect 169820 318500 169876 325052
rect 169820 318434 169876 318444
rect 169932 321748 169988 321758
rect 169820 316372 169876 316382
rect 169820 315028 169876 316316
rect 169932 315140 169988 321692
rect 170492 320068 170548 333116
rect 170492 320002 170548 320012
rect 169932 315074 169988 315084
rect 169820 314962 169876 314972
rect 170492 314356 170548 314366
rect 170492 89908 170548 314300
rect 170604 204036 170660 345884
rect 170716 342580 170772 342590
rect 170716 329252 170772 342524
rect 170716 329186 170772 329196
rect 170604 203970 170660 203980
rect 170716 315700 170772 315710
rect 170716 125188 170772 315644
rect 170828 236292 170884 351932
rect 170940 350644 170996 350654
rect 170940 340340 170996 350588
rect 170940 340274 170996 340284
rect 170828 236226 170884 236236
rect 170940 315028 170996 315038
rect 170940 163828 170996 314972
rect 171052 289044 171108 357308
rect 172508 354676 172564 354686
rect 171276 352660 171332 352670
rect 171276 349468 171332 352604
rect 171276 349412 171444 349468
rect 171164 319060 171220 319070
rect 171164 303268 171220 319004
rect 171164 303202 171220 303212
rect 171052 288978 171108 288988
rect 171388 239876 171444 349412
rect 172396 344596 172452 344606
rect 172284 324436 172340 324446
rect 171388 239810 171444 239820
rect 172172 321076 172228 321086
rect 170940 163762 170996 163772
rect 170716 125122 170772 125132
rect 170492 89842 170548 89852
rect 172172 84868 172228 321020
rect 172284 91588 172340 324380
rect 172396 196868 172452 344540
rect 172508 250628 172564 354620
rect 172620 293636 172676 362684
rect 173180 357588 173236 357598
rect 172620 293570 172676 293580
rect 173068 327348 173124 327358
rect 172508 250562 172564 250572
rect 172396 196802 172452 196812
rect 173068 107268 173124 327292
rect 173180 268548 173236 357532
rect 415772 354004 415828 354014
rect 193808 352350 194128 352384
rect 193808 352294 193878 352350
rect 193934 352294 194002 352350
rect 194058 352294 194128 352350
rect 193808 352226 194128 352294
rect 193808 352170 193878 352226
rect 193934 352170 194002 352226
rect 194058 352170 194128 352226
rect 193808 352102 194128 352170
rect 193808 352046 193878 352102
rect 193934 352046 194002 352102
rect 194058 352046 194128 352102
rect 193808 351978 194128 352046
rect 193808 351922 193878 351978
rect 193934 351922 194002 351978
rect 194058 351922 194128 351978
rect 193808 351888 194128 351922
rect 224528 352350 224848 352384
rect 224528 352294 224598 352350
rect 224654 352294 224722 352350
rect 224778 352294 224848 352350
rect 224528 352226 224848 352294
rect 224528 352170 224598 352226
rect 224654 352170 224722 352226
rect 224778 352170 224848 352226
rect 224528 352102 224848 352170
rect 224528 352046 224598 352102
rect 224654 352046 224722 352102
rect 224778 352046 224848 352102
rect 224528 351978 224848 352046
rect 224528 351922 224598 351978
rect 224654 351922 224722 351978
rect 224778 351922 224848 351978
rect 224528 351888 224848 351922
rect 255248 352350 255568 352384
rect 255248 352294 255318 352350
rect 255374 352294 255442 352350
rect 255498 352294 255568 352350
rect 255248 352226 255568 352294
rect 255248 352170 255318 352226
rect 255374 352170 255442 352226
rect 255498 352170 255568 352226
rect 255248 352102 255568 352170
rect 255248 352046 255318 352102
rect 255374 352046 255442 352102
rect 255498 352046 255568 352102
rect 255248 351978 255568 352046
rect 255248 351922 255318 351978
rect 255374 351922 255442 351978
rect 255498 351922 255568 351978
rect 255248 351888 255568 351922
rect 285968 352350 286288 352384
rect 285968 352294 286038 352350
rect 286094 352294 286162 352350
rect 286218 352294 286288 352350
rect 285968 352226 286288 352294
rect 285968 352170 286038 352226
rect 286094 352170 286162 352226
rect 286218 352170 286288 352226
rect 285968 352102 286288 352170
rect 285968 352046 286038 352102
rect 286094 352046 286162 352102
rect 286218 352046 286288 352102
rect 285968 351978 286288 352046
rect 285968 351922 286038 351978
rect 286094 351922 286162 351978
rect 286218 351922 286288 351978
rect 285968 351888 286288 351922
rect 316688 352350 317008 352384
rect 316688 352294 316758 352350
rect 316814 352294 316882 352350
rect 316938 352294 317008 352350
rect 316688 352226 317008 352294
rect 316688 352170 316758 352226
rect 316814 352170 316882 352226
rect 316938 352170 317008 352226
rect 316688 352102 317008 352170
rect 316688 352046 316758 352102
rect 316814 352046 316882 352102
rect 316938 352046 317008 352102
rect 316688 351978 317008 352046
rect 316688 351922 316758 351978
rect 316814 351922 316882 351978
rect 316938 351922 317008 351978
rect 316688 351888 317008 351922
rect 347408 352350 347728 352384
rect 347408 352294 347478 352350
rect 347534 352294 347602 352350
rect 347658 352294 347728 352350
rect 347408 352226 347728 352294
rect 347408 352170 347478 352226
rect 347534 352170 347602 352226
rect 347658 352170 347728 352226
rect 347408 352102 347728 352170
rect 347408 352046 347478 352102
rect 347534 352046 347602 352102
rect 347658 352046 347728 352102
rect 347408 351978 347728 352046
rect 347408 351922 347478 351978
rect 347534 351922 347602 351978
rect 347658 351922 347728 351978
rect 347408 351888 347728 351922
rect 378128 352350 378448 352384
rect 378128 352294 378198 352350
rect 378254 352294 378322 352350
rect 378378 352294 378448 352350
rect 378128 352226 378448 352294
rect 378128 352170 378198 352226
rect 378254 352170 378322 352226
rect 378378 352170 378448 352226
rect 378128 352102 378448 352170
rect 378128 352046 378198 352102
rect 378254 352046 378322 352102
rect 378378 352046 378448 352102
rect 378128 351978 378448 352046
rect 378128 351922 378198 351978
rect 378254 351922 378322 351978
rect 378378 351922 378448 351978
rect 378128 351888 378448 351922
rect 408848 352350 409168 352384
rect 408848 352294 408918 352350
rect 408974 352294 409042 352350
rect 409098 352294 409168 352350
rect 408848 352226 409168 352294
rect 408848 352170 408918 352226
rect 408974 352170 409042 352226
rect 409098 352170 409168 352226
rect 408848 352102 409168 352170
rect 408848 352046 408918 352102
rect 408974 352046 409042 352102
rect 409098 352046 409168 352102
rect 408848 351978 409168 352046
rect 408848 351922 408918 351978
rect 408974 351922 409042 351978
rect 409098 351922 409168 351978
rect 408848 351888 409168 351922
rect 173180 268482 173236 268492
rect 173740 347284 173796 347294
rect 173740 211204 173796 347228
rect 174076 346612 174132 346622
rect 174076 337708 174132 346556
rect 178448 346350 178768 346384
rect 178448 346294 178518 346350
rect 178574 346294 178642 346350
rect 178698 346294 178768 346350
rect 178448 346226 178768 346294
rect 178448 346170 178518 346226
rect 178574 346170 178642 346226
rect 178698 346170 178768 346226
rect 178448 346102 178768 346170
rect 178448 346046 178518 346102
rect 178574 346046 178642 346102
rect 178698 346046 178768 346102
rect 178448 345978 178768 346046
rect 178448 345922 178518 345978
rect 178574 345922 178642 345978
rect 178698 345922 178768 345978
rect 178448 345888 178768 345922
rect 209168 346350 209488 346384
rect 209168 346294 209238 346350
rect 209294 346294 209362 346350
rect 209418 346294 209488 346350
rect 209168 346226 209488 346294
rect 209168 346170 209238 346226
rect 209294 346170 209362 346226
rect 209418 346170 209488 346226
rect 209168 346102 209488 346170
rect 209168 346046 209238 346102
rect 209294 346046 209362 346102
rect 209418 346046 209488 346102
rect 209168 345978 209488 346046
rect 209168 345922 209238 345978
rect 209294 345922 209362 345978
rect 209418 345922 209488 345978
rect 209168 345888 209488 345922
rect 239888 346350 240208 346384
rect 239888 346294 239958 346350
rect 240014 346294 240082 346350
rect 240138 346294 240208 346350
rect 239888 346226 240208 346294
rect 239888 346170 239958 346226
rect 240014 346170 240082 346226
rect 240138 346170 240208 346226
rect 239888 346102 240208 346170
rect 239888 346046 239958 346102
rect 240014 346046 240082 346102
rect 240138 346046 240208 346102
rect 239888 345978 240208 346046
rect 239888 345922 239958 345978
rect 240014 345922 240082 345978
rect 240138 345922 240208 345978
rect 239888 345888 240208 345922
rect 270608 346350 270928 346384
rect 270608 346294 270678 346350
rect 270734 346294 270802 346350
rect 270858 346294 270928 346350
rect 270608 346226 270928 346294
rect 270608 346170 270678 346226
rect 270734 346170 270802 346226
rect 270858 346170 270928 346226
rect 270608 346102 270928 346170
rect 270608 346046 270678 346102
rect 270734 346046 270802 346102
rect 270858 346046 270928 346102
rect 270608 345978 270928 346046
rect 270608 345922 270678 345978
rect 270734 345922 270802 345978
rect 270858 345922 270928 345978
rect 270608 345888 270928 345922
rect 301328 346350 301648 346384
rect 301328 346294 301398 346350
rect 301454 346294 301522 346350
rect 301578 346294 301648 346350
rect 301328 346226 301648 346294
rect 301328 346170 301398 346226
rect 301454 346170 301522 346226
rect 301578 346170 301648 346226
rect 301328 346102 301648 346170
rect 301328 346046 301398 346102
rect 301454 346046 301522 346102
rect 301578 346046 301648 346102
rect 301328 345978 301648 346046
rect 301328 345922 301398 345978
rect 301454 345922 301522 345978
rect 301578 345922 301648 345978
rect 301328 345888 301648 345922
rect 332048 346350 332368 346384
rect 332048 346294 332118 346350
rect 332174 346294 332242 346350
rect 332298 346294 332368 346350
rect 332048 346226 332368 346294
rect 332048 346170 332118 346226
rect 332174 346170 332242 346226
rect 332298 346170 332368 346226
rect 332048 346102 332368 346170
rect 332048 346046 332118 346102
rect 332174 346046 332242 346102
rect 332298 346046 332368 346102
rect 332048 345978 332368 346046
rect 332048 345922 332118 345978
rect 332174 345922 332242 345978
rect 332298 345922 332368 345978
rect 332048 345888 332368 345922
rect 362768 346350 363088 346384
rect 362768 346294 362838 346350
rect 362894 346294 362962 346350
rect 363018 346294 363088 346350
rect 362768 346226 363088 346294
rect 362768 346170 362838 346226
rect 362894 346170 362962 346226
rect 363018 346170 363088 346226
rect 362768 346102 363088 346170
rect 362768 346046 362838 346102
rect 362894 346046 362962 346102
rect 363018 346046 363088 346102
rect 362768 345978 363088 346046
rect 362768 345922 362838 345978
rect 362894 345922 362962 345978
rect 363018 345922 363088 345978
rect 362768 345888 363088 345922
rect 393488 346350 393808 346384
rect 393488 346294 393558 346350
rect 393614 346294 393682 346350
rect 393738 346294 393808 346350
rect 393488 346226 393808 346294
rect 393488 346170 393558 346226
rect 393614 346170 393682 346226
rect 393738 346170 393808 346226
rect 393488 346102 393808 346170
rect 393488 346046 393558 346102
rect 393614 346046 393682 346102
rect 393738 346046 393808 346102
rect 393488 345978 393808 346046
rect 393488 345922 393558 345978
rect 393614 345922 393682 345978
rect 393738 345922 393808 345978
rect 393488 345888 393808 345922
rect 173964 337652 174132 337708
rect 414092 337764 414148 337774
rect 173740 211138 173796 211148
rect 173852 304138 173908 304148
rect 173068 107202 173124 107212
rect 172284 91522 172340 91532
rect 172172 84802 172228 84812
rect 173852 79044 173908 304082
rect 173964 207620 174020 337652
rect 173964 207554 174020 207564
rect 174076 337204 174132 337214
rect 174076 157444 174132 337148
rect 193808 334350 194128 334384
rect 193808 334294 193878 334350
rect 193934 334294 194002 334350
rect 194058 334294 194128 334350
rect 193808 334226 194128 334294
rect 193808 334170 193878 334226
rect 193934 334170 194002 334226
rect 194058 334170 194128 334226
rect 193808 334102 194128 334170
rect 193808 334046 193878 334102
rect 193934 334046 194002 334102
rect 194058 334046 194128 334102
rect 193808 333978 194128 334046
rect 193808 333922 193878 333978
rect 193934 333922 194002 333978
rect 194058 333922 194128 333978
rect 193808 333888 194128 333922
rect 224528 334350 224848 334384
rect 224528 334294 224598 334350
rect 224654 334294 224722 334350
rect 224778 334294 224848 334350
rect 224528 334226 224848 334294
rect 224528 334170 224598 334226
rect 224654 334170 224722 334226
rect 224778 334170 224848 334226
rect 224528 334102 224848 334170
rect 224528 334046 224598 334102
rect 224654 334046 224722 334102
rect 224778 334046 224848 334102
rect 224528 333978 224848 334046
rect 224528 333922 224598 333978
rect 224654 333922 224722 333978
rect 224778 333922 224848 333978
rect 224528 333888 224848 333922
rect 255248 334350 255568 334384
rect 255248 334294 255318 334350
rect 255374 334294 255442 334350
rect 255498 334294 255568 334350
rect 255248 334226 255568 334294
rect 255248 334170 255318 334226
rect 255374 334170 255442 334226
rect 255498 334170 255568 334226
rect 255248 334102 255568 334170
rect 255248 334046 255318 334102
rect 255374 334046 255442 334102
rect 255498 334046 255568 334102
rect 255248 333978 255568 334046
rect 255248 333922 255318 333978
rect 255374 333922 255442 333978
rect 255498 333922 255568 333978
rect 255248 333888 255568 333922
rect 285968 334350 286288 334384
rect 285968 334294 286038 334350
rect 286094 334294 286162 334350
rect 286218 334294 286288 334350
rect 285968 334226 286288 334294
rect 285968 334170 286038 334226
rect 286094 334170 286162 334226
rect 286218 334170 286288 334226
rect 285968 334102 286288 334170
rect 285968 334046 286038 334102
rect 286094 334046 286162 334102
rect 286218 334046 286288 334102
rect 285968 333978 286288 334046
rect 285968 333922 286038 333978
rect 286094 333922 286162 333978
rect 286218 333922 286288 333978
rect 285968 333888 286288 333922
rect 316688 334350 317008 334384
rect 316688 334294 316758 334350
rect 316814 334294 316882 334350
rect 316938 334294 317008 334350
rect 316688 334226 317008 334294
rect 316688 334170 316758 334226
rect 316814 334170 316882 334226
rect 316938 334170 317008 334226
rect 316688 334102 317008 334170
rect 316688 334046 316758 334102
rect 316814 334046 316882 334102
rect 316938 334046 317008 334102
rect 316688 333978 317008 334046
rect 316688 333922 316758 333978
rect 316814 333922 316882 333978
rect 316938 333922 317008 333978
rect 316688 333888 317008 333922
rect 347408 334350 347728 334384
rect 347408 334294 347478 334350
rect 347534 334294 347602 334350
rect 347658 334294 347728 334350
rect 347408 334226 347728 334294
rect 347408 334170 347478 334226
rect 347534 334170 347602 334226
rect 347658 334170 347728 334226
rect 347408 334102 347728 334170
rect 347408 334046 347478 334102
rect 347534 334046 347602 334102
rect 347658 334046 347728 334102
rect 347408 333978 347728 334046
rect 347408 333922 347478 333978
rect 347534 333922 347602 333978
rect 347658 333922 347728 333978
rect 347408 333888 347728 333922
rect 378128 334350 378448 334384
rect 378128 334294 378198 334350
rect 378254 334294 378322 334350
rect 378378 334294 378448 334350
rect 378128 334226 378448 334294
rect 378128 334170 378198 334226
rect 378254 334170 378322 334226
rect 378378 334170 378448 334226
rect 378128 334102 378448 334170
rect 378128 334046 378198 334102
rect 378254 334046 378322 334102
rect 378378 334046 378448 334102
rect 378128 333978 378448 334046
rect 378128 333922 378198 333978
rect 378254 333922 378322 333978
rect 378378 333922 378448 333978
rect 378128 333888 378448 333922
rect 408848 334350 409168 334384
rect 408848 334294 408918 334350
rect 408974 334294 409042 334350
rect 409098 334294 409168 334350
rect 408848 334226 409168 334294
rect 408848 334170 408918 334226
rect 408974 334170 409042 334226
rect 409098 334170 409168 334226
rect 408848 334102 409168 334170
rect 408848 334046 408918 334102
rect 408974 334046 409042 334102
rect 409098 334046 409168 334102
rect 408848 333978 409168 334046
rect 408848 333922 408918 333978
rect 408974 333922 409042 333978
rect 409098 333922 409168 333978
rect 408848 333888 409168 333922
rect 178448 328350 178768 328384
rect 178448 328294 178518 328350
rect 178574 328294 178642 328350
rect 178698 328294 178768 328350
rect 178448 328226 178768 328294
rect 178448 328170 178518 328226
rect 178574 328170 178642 328226
rect 178698 328170 178768 328226
rect 178448 328102 178768 328170
rect 178448 328046 178518 328102
rect 178574 328046 178642 328102
rect 178698 328046 178768 328102
rect 178448 327978 178768 328046
rect 178448 327922 178518 327978
rect 178574 327922 178642 327978
rect 178698 327922 178768 327978
rect 178448 327888 178768 327922
rect 209168 328350 209488 328384
rect 209168 328294 209238 328350
rect 209294 328294 209362 328350
rect 209418 328294 209488 328350
rect 209168 328226 209488 328294
rect 209168 328170 209238 328226
rect 209294 328170 209362 328226
rect 209418 328170 209488 328226
rect 209168 328102 209488 328170
rect 209168 328046 209238 328102
rect 209294 328046 209362 328102
rect 209418 328046 209488 328102
rect 209168 327978 209488 328046
rect 209168 327922 209238 327978
rect 209294 327922 209362 327978
rect 209418 327922 209488 327978
rect 209168 327888 209488 327922
rect 239888 328350 240208 328384
rect 239888 328294 239958 328350
rect 240014 328294 240082 328350
rect 240138 328294 240208 328350
rect 239888 328226 240208 328294
rect 239888 328170 239958 328226
rect 240014 328170 240082 328226
rect 240138 328170 240208 328226
rect 239888 328102 240208 328170
rect 239888 328046 239958 328102
rect 240014 328046 240082 328102
rect 240138 328046 240208 328102
rect 239888 327978 240208 328046
rect 239888 327922 239958 327978
rect 240014 327922 240082 327978
rect 240138 327922 240208 327978
rect 239888 327888 240208 327922
rect 270608 328350 270928 328384
rect 270608 328294 270678 328350
rect 270734 328294 270802 328350
rect 270858 328294 270928 328350
rect 270608 328226 270928 328294
rect 270608 328170 270678 328226
rect 270734 328170 270802 328226
rect 270858 328170 270928 328226
rect 270608 328102 270928 328170
rect 270608 328046 270678 328102
rect 270734 328046 270802 328102
rect 270858 328046 270928 328102
rect 270608 327978 270928 328046
rect 270608 327922 270678 327978
rect 270734 327922 270802 327978
rect 270858 327922 270928 327978
rect 270608 327888 270928 327922
rect 301328 328350 301648 328384
rect 301328 328294 301398 328350
rect 301454 328294 301522 328350
rect 301578 328294 301648 328350
rect 301328 328226 301648 328294
rect 301328 328170 301398 328226
rect 301454 328170 301522 328226
rect 301578 328170 301648 328226
rect 301328 328102 301648 328170
rect 301328 328046 301398 328102
rect 301454 328046 301522 328102
rect 301578 328046 301648 328102
rect 301328 327978 301648 328046
rect 301328 327922 301398 327978
rect 301454 327922 301522 327978
rect 301578 327922 301648 327978
rect 301328 327888 301648 327922
rect 332048 328350 332368 328384
rect 332048 328294 332118 328350
rect 332174 328294 332242 328350
rect 332298 328294 332368 328350
rect 332048 328226 332368 328294
rect 332048 328170 332118 328226
rect 332174 328170 332242 328226
rect 332298 328170 332368 328226
rect 332048 328102 332368 328170
rect 332048 328046 332118 328102
rect 332174 328046 332242 328102
rect 332298 328046 332368 328102
rect 332048 327978 332368 328046
rect 332048 327922 332118 327978
rect 332174 327922 332242 327978
rect 332298 327922 332368 327978
rect 332048 327888 332368 327922
rect 362768 328350 363088 328384
rect 362768 328294 362838 328350
rect 362894 328294 362962 328350
rect 363018 328294 363088 328350
rect 362768 328226 363088 328294
rect 362768 328170 362838 328226
rect 362894 328170 362962 328226
rect 363018 328170 363088 328226
rect 362768 328102 363088 328170
rect 362768 328046 362838 328102
rect 362894 328046 362962 328102
rect 363018 328046 363088 328102
rect 362768 327978 363088 328046
rect 362768 327922 362838 327978
rect 362894 327922 362962 327978
rect 363018 327922 363088 327978
rect 362768 327888 363088 327922
rect 393488 328350 393808 328384
rect 393488 328294 393558 328350
rect 393614 328294 393682 328350
rect 393738 328294 393808 328350
rect 393488 328226 393808 328294
rect 393488 328170 393558 328226
rect 393614 328170 393682 328226
rect 393738 328170 393808 328226
rect 393488 328102 393808 328170
rect 393488 328046 393558 328102
rect 393614 328046 393682 328102
rect 393738 328046 393808 328102
rect 393488 327978 393808 328046
rect 393488 327922 393558 327978
rect 393614 327922 393682 327978
rect 393738 327922 393808 327978
rect 393488 327888 393808 327922
rect 193808 316350 194128 316384
rect 193808 316294 193878 316350
rect 193934 316294 194002 316350
rect 194058 316294 194128 316350
rect 193808 316226 194128 316294
rect 193808 316170 193878 316226
rect 193934 316170 194002 316226
rect 194058 316170 194128 316226
rect 193808 316102 194128 316170
rect 193808 316046 193878 316102
rect 193934 316046 194002 316102
rect 194058 316046 194128 316102
rect 193808 315978 194128 316046
rect 193808 315922 193878 315978
rect 193934 315922 194002 315978
rect 194058 315922 194128 315978
rect 193808 315888 194128 315922
rect 224528 316350 224848 316384
rect 224528 316294 224598 316350
rect 224654 316294 224722 316350
rect 224778 316294 224848 316350
rect 224528 316226 224848 316294
rect 224528 316170 224598 316226
rect 224654 316170 224722 316226
rect 224778 316170 224848 316226
rect 224528 316102 224848 316170
rect 224528 316046 224598 316102
rect 224654 316046 224722 316102
rect 224778 316046 224848 316102
rect 224528 315978 224848 316046
rect 224528 315922 224598 315978
rect 224654 315922 224722 315978
rect 224778 315922 224848 315978
rect 224528 315888 224848 315922
rect 255248 316350 255568 316384
rect 255248 316294 255318 316350
rect 255374 316294 255442 316350
rect 255498 316294 255568 316350
rect 255248 316226 255568 316294
rect 255248 316170 255318 316226
rect 255374 316170 255442 316226
rect 255498 316170 255568 316226
rect 255248 316102 255568 316170
rect 255248 316046 255318 316102
rect 255374 316046 255442 316102
rect 255498 316046 255568 316102
rect 255248 315978 255568 316046
rect 255248 315922 255318 315978
rect 255374 315922 255442 315978
rect 255498 315922 255568 315978
rect 255248 315888 255568 315922
rect 285968 316350 286288 316384
rect 285968 316294 286038 316350
rect 286094 316294 286162 316350
rect 286218 316294 286288 316350
rect 285968 316226 286288 316294
rect 285968 316170 286038 316226
rect 286094 316170 286162 316226
rect 286218 316170 286288 316226
rect 285968 316102 286288 316170
rect 285968 316046 286038 316102
rect 286094 316046 286162 316102
rect 286218 316046 286288 316102
rect 285968 315978 286288 316046
rect 285968 315922 286038 315978
rect 286094 315922 286162 315978
rect 286218 315922 286288 315978
rect 285968 315888 286288 315922
rect 316688 316350 317008 316384
rect 316688 316294 316758 316350
rect 316814 316294 316882 316350
rect 316938 316294 317008 316350
rect 316688 316226 317008 316294
rect 316688 316170 316758 316226
rect 316814 316170 316882 316226
rect 316938 316170 317008 316226
rect 316688 316102 317008 316170
rect 316688 316046 316758 316102
rect 316814 316046 316882 316102
rect 316938 316046 317008 316102
rect 316688 315978 317008 316046
rect 316688 315922 316758 315978
rect 316814 315922 316882 315978
rect 316938 315922 317008 315978
rect 316688 315888 317008 315922
rect 347408 316350 347728 316384
rect 347408 316294 347478 316350
rect 347534 316294 347602 316350
rect 347658 316294 347728 316350
rect 347408 316226 347728 316294
rect 347408 316170 347478 316226
rect 347534 316170 347602 316226
rect 347658 316170 347728 316226
rect 347408 316102 347728 316170
rect 347408 316046 347478 316102
rect 347534 316046 347602 316102
rect 347658 316046 347728 316102
rect 347408 315978 347728 316046
rect 347408 315922 347478 315978
rect 347534 315922 347602 315978
rect 347658 315922 347728 315978
rect 347408 315888 347728 315922
rect 378128 316350 378448 316384
rect 378128 316294 378198 316350
rect 378254 316294 378322 316350
rect 378378 316294 378448 316350
rect 378128 316226 378448 316294
rect 378128 316170 378198 316226
rect 378254 316170 378322 316226
rect 378378 316170 378448 316226
rect 378128 316102 378448 316170
rect 378128 316046 378198 316102
rect 378254 316046 378322 316102
rect 378378 316046 378448 316102
rect 378128 315978 378448 316046
rect 378128 315922 378198 315978
rect 378254 315922 378322 315978
rect 378378 315922 378448 315978
rect 378128 315888 378448 315922
rect 408848 316350 409168 316384
rect 408848 316294 408918 316350
rect 408974 316294 409042 316350
rect 409098 316294 409168 316350
rect 408848 316226 409168 316294
rect 408848 316170 408918 316226
rect 408974 316170 409042 316226
rect 409098 316170 409168 316226
rect 408848 316102 409168 316170
rect 408848 316046 408918 316102
rect 408974 316046 409042 316102
rect 409098 316046 409168 316102
rect 408848 315978 409168 316046
rect 408848 315922 408918 315978
rect 408974 315922 409042 315978
rect 409098 315922 409168 315978
rect 408848 315888 409168 315922
rect 272188 305732 272244 305742
rect 191772 304500 191828 304510
rect 191772 303156 191828 304444
rect 272188 304138 272244 305676
rect 272188 304072 272244 304082
rect 273980 305284 274036 305294
rect 191772 303090 191828 303100
rect 228732 301618 228788 301628
rect 218428 301258 218484 301268
rect 218428 300804 218484 301202
rect 218428 300738 218484 300748
rect 228732 300804 228788 301562
rect 228732 300738 228788 300748
rect 229180 301438 229236 301448
rect 229180 300804 229236 301382
rect 260540 301078 260596 301088
rect 229180 300738 229236 300748
rect 242172 300898 242228 300908
rect 242172 300804 242228 300842
rect 242172 300738 242228 300748
rect 260540 300804 260596 301022
rect 260540 300738 260596 300748
rect 237692 300178 237748 300188
rect 217980 299998 218036 300008
rect 217980 299460 218036 299942
rect 223356 299818 223412 299828
rect 223356 299572 223412 299762
rect 223356 299506 223412 299516
rect 237692 299572 237748 300122
rect 237692 299506 237748 299516
rect 217980 299394 218036 299404
rect 255612 298340 255668 298350
rect 255612 296996 255668 298284
rect 255612 296930 255668 296940
rect 260092 298340 260148 298350
rect 260092 296884 260148 298284
rect 260092 296818 260148 296828
rect 178448 292350 178768 292384
rect 178448 292294 178518 292350
rect 178574 292294 178642 292350
rect 178698 292294 178768 292350
rect 178448 292226 178768 292294
rect 178448 292170 178518 292226
rect 178574 292170 178642 292226
rect 178698 292170 178768 292226
rect 178448 292102 178768 292170
rect 178448 292046 178518 292102
rect 178574 292046 178642 292102
rect 178698 292046 178768 292102
rect 178448 291978 178768 292046
rect 178448 291922 178518 291978
rect 178574 291922 178642 291978
rect 178698 291922 178768 291978
rect 178448 291888 178768 291922
rect 209168 292350 209488 292384
rect 209168 292294 209238 292350
rect 209294 292294 209362 292350
rect 209418 292294 209488 292350
rect 209168 292226 209488 292294
rect 209168 292170 209238 292226
rect 209294 292170 209362 292226
rect 209418 292170 209488 292226
rect 209168 292102 209488 292170
rect 209168 292046 209238 292102
rect 209294 292046 209362 292102
rect 209418 292046 209488 292102
rect 209168 291978 209488 292046
rect 209168 291922 209238 291978
rect 209294 291922 209362 291978
rect 209418 291922 209488 291978
rect 209168 291888 209488 291922
rect 239888 292350 240208 292384
rect 239888 292294 239958 292350
rect 240014 292294 240082 292350
rect 240138 292294 240208 292350
rect 239888 292226 240208 292294
rect 239888 292170 239958 292226
rect 240014 292170 240082 292226
rect 240138 292170 240208 292226
rect 239888 292102 240208 292170
rect 239888 292046 239958 292102
rect 240014 292046 240082 292102
rect 240138 292046 240208 292102
rect 239888 291978 240208 292046
rect 239888 291922 239958 291978
rect 240014 291922 240082 291978
rect 240138 291922 240208 291978
rect 239888 291888 240208 291922
rect 270608 292350 270928 292384
rect 270608 292294 270678 292350
rect 270734 292294 270802 292350
rect 270858 292294 270928 292350
rect 270608 292226 270928 292294
rect 270608 292170 270678 292226
rect 270734 292170 270802 292226
rect 270858 292170 270928 292226
rect 270608 292102 270928 292170
rect 270608 292046 270678 292102
rect 270734 292046 270802 292102
rect 270858 292046 270928 292102
rect 270608 291978 270928 292046
rect 270608 291922 270678 291978
rect 270734 291922 270802 291978
rect 270858 291922 270928 291978
rect 270608 291888 270928 291922
rect 273980 290668 274036 305228
rect 273868 290612 274036 290668
rect 281898 292350 282518 306466
rect 281898 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 282518 292350
rect 281898 292226 282518 292294
rect 281898 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 282518 292226
rect 281898 292102 282518 292170
rect 281898 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 282518 292102
rect 281898 291978 282518 292046
rect 281898 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 282518 291978
rect 193808 280350 194128 280384
rect 193808 280294 193878 280350
rect 193934 280294 194002 280350
rect 194058 280294 194128 280350
rect 193808 280226 194128 280294
rect 193808 280170 193878 280226
rect 193934 280170 194002 280226
rect 194058 280170 194128 280226
rect 193808 280102 194128 280170
rect 193808 280046 193878 280102
rect 193934 280046 194002 280102
rect 194058 280046 194128 280102
rect 193808 279978 194128 280046
rect 193808 279922 193878 279978
rect 193934 279922 194002 279978
rect 194058 279922 194128 279978
rect 193808 279888 194128 279922
rect 224528 280350 224848 280384
rect 224528 280294 224598 280350
rect 224654 280294 224722 280350
rect 224778 280294 224848 280350
rect 224528 280226 224848 280294
rect 224528 280170 224598 280226
rect 224654 280170 224722 280226
rect 224778 280170 224848 280226
rect 224528 280102 224848 280170
rect 224528 280046 224598 280102
rect 224654 280046 224722 280102
rect 224778 280046 224848 280102
rect 224528 279978 224848 280046
rect 224528 279922 224598 279978
rect 224654 279922 224722 279978
rect 224778 279922 224848 279978
rect 224528 279888 224848 279922
rect 255248 280350 255568 280384
rect 255248 280294 255318 280350
rect 255374 280294 255442 280350
rect 255498 280294 255568 280350
rect 255248 280226 255568 280294
rect 255248 280170 255318 280226
rect 255374 280170 255442 280226
rect 255498 280170 255568 280226
rect 255248 280102 255568 280170
rect 255248 280046 255318 280102
rect 255374 280046 255442 280102
rect 255498 280046 255568 280102
rect 255248 279978 255568 280046
rect 255248 279922 255318 279978
rect 255374 279922 255442 279978
rect 255498 279922 255568 279978
rect 255248 279888 255568 279922
rect 178448 274350 178768 274384
rect 178448 274294 178518 274350
rect 178574 274294 178642 274350
rect 178698 274294 178768 274350
rect 178448 274226 178768 274294
rect 178448 274170 178518 274226
rect 178574 274170 178642 274226
rect 178698 274170 178768 274226
rect 178448 274102 178768 274170
rect 178448 274046 178518 274102
rect 178574 274046 178642 274102
rect 178698 274046 178768 274102
rect 178448 273978 178768 274046
rect 178448 273922 178518 273978
rect 178574 273922 178642 273978
rect 178698 273922 178768 273978
rect 178448 273888 178768 273922
rect 209168 274350 209488 274384
rect 209168 274294 209238 274350
rect 209294 274294 209362 274350
rect 209418 274294 209488 274350
rect 209168 274226 209488 274294
rect 209168 274170 209238 274226
rect 209294 274170 209362 274226
rect 209418 274170 209488 274226
rect 209168 274102 209488 274170
rect 209168 274046 209238 274102
rect 209294 274046 209362 274102
rect 209418 274046 209488 274102
rect 209168 273978 209488 274046
rect 209168 273922 209238 273978
rect 209294 273922 209362 273978
rect 209418 273922 209488 273978
rect 209168 273888 209488 273922
rect 239888 274350 240208 274384
rect 239888 274294 239958 274350
rect 240014 274294 240082 274350
rect 240138 274294 240208 274350
rect 239888 274226 240208 274294
rect 239888 274170 239958 274226
rect 240014 274170 240082 274226
rect 240138 274170 240208 274226
rect 239888 274102 240208 274170
rect 239888 274046 239958 274102
rect 240014 274046 240082 274102
rect 240138 274046 240208 274102
rect 239888 273978 240208 274046
rect 239888 273922 239958 273978
rect 240014 273922 240082 273978
rect 240138 273922 240208 273978
rect 239888 273888 240208 273922
rect 270608 274350 270928 274384
rect 270608 274294 270678 274350
rect 270734 274294 270802 274350
rect 270858 274294 270928 274350
rect 270608 274226 270928 274294
rect 270608 274170 270678 274226
rect 270734 274170 270802 274226
rect 270858 274170 270928 274226
rect 270608 274102 270928 274170
rect 270608 274046 270678 274102
rect 270734 274046 270802 274102
rect 270858 274046 270928 274102
rect 270608 273978 270928 274046
rect 270608 273922 270678 273978
rect 270734 273922 270802 273978
rect 270858 273922 270928 273978
rect 270608 273888 270928 273922
rect 193808 262350 194128 262384
rect 193808 262294 193878 262350
rect 193934 262294 194002 262350
rect 194058 262294 194128 262350
rect 193808 262226 194128 262294
rect 193808 262170 193878 262226
rect 193934 262170 194002 262226
rect 194058 262170 194128 262226
rect 193808 262102 194128 262170
rect 193808 262046 193878 262102
rect 193934 262046 194002 262102
rect 194058 262046 194128 262102
rect 193808 261978 194128 262046
rect 193808 261922 193878 261978
rect 193934 261922 194002 261978
rect 194058 261922 194128 261978
rect 193808 261888 194128 261922
rect 224528 262350 224848 262384
rect 224528 262294 224598 262350
rect 224654 262294 224722 262350
rect 224778 262294 224848 262350
rect 224528 262226 224848 262294
rect 224528 262170 224598 262226
rect 224654 262170 224722 262226
rect 224778 262170 224848 262226
rect 224528 262102 224848 262170
rect 224528 262046 224598 262102
rect 224654 262046 224722 262102
rect 224778 262046 224848 262102
rect 224528 261978 224848 262046
rect 224528 261922 224598 261978
rect 224654 261922 224722 261978
rect 224778 261922 224848 261978
rect 224528 261888 224848 261922
rect 255248 262350 255568 262384
rect 255248 262294 255318 262350
rect 255374 262294 255442 262350
rect 255498 262294 255568 262350
rect 255248 262226 255568 262294
rect 255248 262170 255318 262226
rect 255374 262170 255442 262226
rect 255498 262170 255568 262226
rect 255248 262102 255568 262170
rect 255248 262046 255318 262102
rect 255374 262046 255442 262102
rect 255498 262046 255568 262102
rect 255248 261978 255568 262046
rect 255248 261922 255318 261978
rect 255374 261922 255442 261978
rect 255498 261922 255568 261978
rect 255248 261888 255568 261922
rect 178448 256350 178768 256384
rect 178448 256294 178518 256350
rect 178574 256294 178642 256350
rect 178698 256294 178768 256350
rect 178448 256226 178768 256294
rect 178448 256170 178518 256226
rect 178574 256170 178642 256226
rect 178698 256170 178768 256226
rect 178448 256102 178768 256170
rect 178448 256046 178518 256102
rect 178574 256046 178642 256102
rect 178698 256046 178768 256102
rect 178448 255978 178768 256046
rect 178448 255922 178518 255978
rect 178574 255922 178642 255978
rect 178698 255922 178768 255978
rect 178448 255888 178768 255922
rect 209168 256350 209488 256384
rect 209168 256294 209238 256350
rect 209294 256294 209362 256350
rect 209418 256294 209488 256350
rect 209168 256226 209488 256294
rect 209168 256170 209238 256226
rect 209294 256170 209362 256226
rect 209418 256170 209488 256226
rect 209168 256102 209488 256170
rect 209168 256046 209238 256102
rect 209294 256046 209362 256102
rect 209418 256046 209488 256102
rect 209168 255978 209488 256046
rect 209168 255922 209238 255978
rect 209294 255922 209362 255978
rect 209418 255922 209488 255978
rect 209168 255888 209488 255922
rect 239888 256350 240208 256384
rect 239888 256294 239958 256350
rect 240014 256294 240082 256350
rect 240138 256294 240208 256350
rect 239888 256226 240208 256294
rect 239888 256170 239958 256226
rect 240014 256170 240082 256226
rect 240138 256170 240208 256226
rect 239888 256102 240208 256170
rect 239888 256046 239958 256102
rect 240014 256046 240082 256102
rect 240138 256046 240208 256102
rect 239888 255978 240208 256046
rect 239888 255922 239958 255978
rect 240014 255922 240082 255978
rect 240138 255922 240208 255978
rect 239888 255888 240208 255922
rect 270608 256350 270928 256384
rect 270608 256294 270678 256350
rect 270734 256294 270802 256350
rect 270858 256294 270928 256350
rect 270608 256226 270928 256294
rect 270608 256170 270678 256226
rect 270734 256170 270802 256226
rect 270858 256170 270928 256226
rect 270608 256102 270928 256170
rect 270608 256046 270678 256102
rect 270734 256046 270802 256102
rect 270858 256046 270928 256102
rect 270608 255978 270928 256046
rect 270608 255922 270678 255978
rect 270734 255922 270802 255978
rect 270858 255922 270928 255978
rect 270608 255888 270928 255922
rect 193808 244350 194128 244384
rect 193808 244294 193878 244350
rect 193934 244294 194002 244350
rect 194058 244294 194128 244350
rect 193808 244226 194128 244294
rect 193808 244170 193878 244226
rect 193934 244170 194002 244226
rect 194058 244170 194128 244226
rect 193808 244102 194128 244170
rect 193808 244046 193878 244102
rect 193934 244046 194002 244102
rect 194058 244046 194128 244102
rect 193808 243978 194128 244046
rect 193808 243922 193878 243978
rect 193934 243922 194002 243978
rect 194058 243922 194128 243978
rect 193808 243888 194128 243922
rect 224528 244350 224848 244384
rect 224528 244294 224598 244350
rect 224654 244294 224722 244350
rect 224778 244294 224848 244350
rect 224528 244226 224848 244294
rect 224528 244170 224598 244226
rect 224654 244170 224722 244226
rect 224778 244170 224848 244226
rect 224528 244102 224848 244170
rect 224528 244046 224598 244102
rect 224654 244046 224722 244102
rect 224778 244046 224848 244102
rect 224528 243978 224848 244046
rect 224528 243922 224598 243978
rect 224654 243922 224722 243978
rect 224778 243922 224848 243978
rect 224528 243888 224848 243922
rect 255248 244350 255568 244384
rect 255248 244294 255318 244350
rect 255374 244294 255442 244350
rect 255498 244294 255568 244350
rect 255248 244226 255568 244294
rect 255248 244170 255318 244226
rect 255374 244170 255442 244226
rect 255498 244170 255568 244226
rect 255248 244102 255568 244170
rect 255248 244046 255318 244102
rect 255374 244046 255442 244102
rect 255498 244046 255568 244102
rect 255248 243978 255568 244046
rect 255248 243922 255318 243978
rect 255374 243922 255442 243978
rect 255498 243922 255568 243978
rect 255248 243888 255568 243922
rect 178448 238350 178768 238384
rect 178448 238294 178518 238350
rect 178574 238294 178642 238350
rect 178698 238294 178768 238350
rect 178448 238226 178768 238294
rect 178448 238170 178518 238226
rect 178574 238170 178642 238226
rect 178698 238170 178768 238226
rect 178448 238102 178768 238170
rect 178448 238046 178518 238102
rect 178574 238046 178642 238102
rect 178698 238046 178768 238102
rect 178448 237978 178768 238046
rect 178448 237922 178518 237978
rect 178574 237922 178642 237978
rect 178698 237922 178768 237978
rect 178448 237888 178768 237922
rect 209168 238350 209488 238384
rect 209168 238294 209238 238350
rect 209294 238294 209362 238350
rect 209418 238294 209488 238350
rect 209168 238226 209488 238294
rect 209168 238170 209238 238226
rect 209294 238170 209362 238226
rect 209418 238170 209488 238226
rect 209168 238102 209488 238170
rect 209168 238046 209238 238102
rect 209294 238046 209362 238102
rect 209418 238046 209488 238102
rect 209168 237978 209488 238046
rect 209168 237922 209238 237978
rect 209294 237922 209362 237978
rect 209418 237922 209488 237978
rect 209168 237888 209488 237922
rect 239888 238350 240208 238384
rect 239888 238294 239958 238350
rect 240014 238294 240082 238350
rect 240138 238294 240208 238350
rect 239888 238226 240208 238294
rect 239888 238170 239958 238226
rect 240014 238170 240082 238226
rect 240138 238170 240208 238226
rect 239888 238102 240208 238170
rect 239888 238046 239958 238102
rect 240014 238046 240082 238102
rect 240138 238046 240208 238102
rect 239888 237978 240208 238046
rect 239888 237922 239958 237978
rect 240014 237922 240082 237978
rect 240138 237922 240208 237978
rect 239888 237888 240208 237922
rect 270608 238350 270928 238384
rect 270608 238294 270678 238350
rect 270734 238294 270802 238350
rect 270858 238294 270928 238350
rect 270608 238226 270928 238294
rect 270608 238170 270678 238226
rect 270734 238170 270802 238226
rect 270858 238170 270928 238226
rect 270608 238102 270928 238170
rect 270608 238046 270678 238102
rect 270734 238046 270802 238102
rect 270858 238046 270928 238102
rect 270608 237978 270928 238046
rect 270608 237922 270678 237978
rect 270734 237922 270802 237978
rect 270858 237922 270928 237978
rect 270608 237888 270928 237922
rect 272972 236852 273028 236862
rect 193808 226350 194128 226384
rect 193808 226294 193878 226350
rect 193934 226294 194002 226350
rect 194058 226294 194128 226350
rect 193808 226226 194128 226294
rect 193808 226170 193878 226226
rect 193934 226170 194002 226226
rect 194058 226170 194128 226226
rect 193808 226102 194128 226170
rect 193808 226046 193878 226102
rect 193934 226046 194002 226102
rect 194058 226046 194128 226102
rect 193808 225978 194128 226046
rect 193808 225922 193878 225978
rect 193934 225922 194002 225978
rect 194058 225922 194128 225978
rect 193808 225888 194128 225922
rect 224528 226350 224848 226384
rect 224528 226294 224598 226350
rect 224654 226294 224722 226350
rect 224778 226294 224848 226350
rect 224528 226226 224848 226294
rect 224528 226170 224598 226226
rect 224654 226170 224722 226226
rect 224778 226170 224848 226226
rect 224528 226102 224848 226170
rect 224528 226046 224598 226102
rect 224654 226046 224722 226102
rect 224778 226046 224848 226102
rect 224528 225978 224848 226046
rect 224528 225922 224598 225978
rect 224654 225922 224722 225978
rect 224778 225922 224848 225978
rect 224528 225888 224848 225922
rect 255248 226350 255568 226384
rect 255248 226294 255318 226350
rect 255374 226294 255442 226350
rect 255498 226294 255568 226350
rect 255248 226226 255568 226294
rect 255248 226170 255318 226226
rect 255374 226170 255442 226226
rect 255498 226170 255568 226226
rect 255248 226102 255568 226170
rect 255248 226046 255318 226102
rect 255374 226046 255442 226102
rect 255498 226046 255568 226102
rect 255248 225978 255568 226046
rect 255248 225922 255318 225978
rect 255374 225922 255442 225978
rect 255498 225922 255568 225978
rect 255248 225888 255568 225922
rect 178448 220350 178768 220384
rect 178448 220294 178518 220350
rect 178574 220294 178642 220350
rect 178698 220294 178768 220350
rect 178448 220226 178768 220294
rect 178448 220170 178518 220226
rect 178574 220170 178642 220226
rect 178698 220170 178768 220226
rect 178448 220102 178768 220170
rect 178448 220046 178518 220102
rect 178574 220046 178642 220102
rect 178698 220046 178768 220102
rect 178448 219978 178768 220046
rect 178448 219922 178518 219978
rect 178574 219922 178642 219978
rect 178698 219922 178768 219978
rect 178448 219888 178768 219922
rect 209168 220350 209488 220384
rect 209168 220294 209238 220350
rect 209294 220294 209362 220350
rect 209418 220294 209488 220350
rect 209168 220226 209488 220294
rect 209168 220170 209238 220226
rect 209294 220170 209362 220226
rect 209418 220170 209488 220226
rect 209168 220102 209488 220170
rect 209168 220046 209238 220102
rect 209294 220046 209362 220102
rect 209418 220046 209488 220102
rect 209168 219978 209488 220046
rect 209168 219922 209238 219978
rect 209294 219922 209362 219978
rect 209418 219922 209488 219978
rect 209168 219888 209488 219922
rect 239888 220350 240208 220384
rect 239888 220294 239958 220350
rect 240014 220294 240082 220350
rect 240138 220294 240208 220350
rect 239888 220226 240208 220294
rect 239888 220170 239958 220226
rect 240014 220170 240082 220226
rect 240138 220170 240208 220226
rect 239888 220102 240208 220170
rect 239888 220046 239958 220102
rect 240014 220046 240082 220102
rect 240138 220046 240208 220102
rect 239888 219978 240208 220046
rect 239888 219922 239958 219978
rect 240014 219922 240082 219978
rect 240138 219922 240208 219978
rect 239888 219888 240208 219922
rect 270608 220350 270928 220384
rect 270608 220294 270678 220350
rect 270734 220294 270802 220350
rect 270858 220294 270928 220350
rect 270608 220226 270928 220294
rect 270608 220170 270678 220226
rect 270734 220170 270802 220226
rect 270858 220170 270928 220226
rect 270608 220102 270928 220170
rect 270608 220046 270678 220102
rect 270734 220046 270802 220102
rect 270858 220046 270928 220102
rect 270608 219978 270928 220046
rect 270608 219922 270678 219978
rect 270734 219922 270802 219978
rect 270858 219922 270928 219978
rect 270608 219888 270928 219922
rect 193808 208350 194128 208384
rect 193808 208294 193878 208350
rect 193934 208294 194002 208350
rect 194058 208294 194128 208350
rect 193808 208226 194128 208294
rect 193808 208170 193878 208226
rect 193934 208170 194002 208226
rect 194058 208170 194128 208226
rect 193808 208102 194128 208170
rect 193808 208046 193878 208102
rect 193934 208046 194002 208102
rect 194058 208046 194128 208102
rect 193808 207978 194128 208046
rect 193808 207922 193878 207978
rect 193934 207922 194002 207978
rect 194058 207922 194128 207978
rect 193808 207888 194128 207922
rect 224528 208350 224848 208384
rect 224528 208294 224598 208350
rect 224654 208294 224722 208350
rect 224778 208294 224848 208350
rect 224528 208226 224848 208294
rect 224528 208170 224598 208226
rect 224654 208170 224722 208226
rect 224778 208170 224848 208226
rect 224528 208102 224848 208170
rect 224528 208046 224598 208102
rect 224654 208046 224722 208102
rect 224778 208046 224848 208102
rect 224528 207978 224848 208046
rect 224528 207922 224598 207978
rect 224654 207922 224722 207978
rect 224778 207922 224848 207978
rect 224528 207888 224848 207922
rect 255248 208350 255568 208384
rect 255248 208294 255318 208350
rect 255374 208294 255442 208350
rect 255498 208294 255568 208350
rect 255248 208226 255568 208294
rect 255248 208170 255318 208226
rect 255374 208170 255442 208226
rect 255498 208170 255568 208226
rect 255248 208102 255568 208170
rect 255248 208046 255318 208102
rect 255374 208046 255442 208102
rect 255498 208046 255568 208102
rect 255248 207978 255568 208046
rect 255248 207922 255318 207978
rect 255374 207922 255442 207978
rect 255498 207922 255568 207978
rect 255248 207888 255568 207922
rect 178448 202350 178768 202384
rect 178448 202294 178518 202350
rect 178574 202294 178642 202350
rect 178698 202294 178768 202350
rect 178448 202226 178768 202294
rect 178448 202170 178518 202226
rect 178574 202170 178642 202226
rect 178698 202170 178768 202226
rect 178448 202102 178768 202170
rect 178448 202046 178518 202102
rect 178574 202046 178642 202102
rect 178698 202046 178768 202102
rect 178448 201978 178768 202046
rect 178448 201922 178518 201978
rect 178574 201922 178642 201978
rect 178698 201922 178768 201978
rect 178448 201888 178768 201922
rect 209168 202350 209488 202384
rect 209168 202294 209238 202350
rect 209294 202294 209362 202350
rect 209418 202294 209488 202350
rect 209168 202226 209488 202294
rect 209168 202170 209238 202226
rect 209294 202170 209362 202226
rect 209418 202170 209488 202226
rect 209168 202102 209488 202170
rect 209168 202046 209238 202102
rect 209294 202046 209362 202102
rect 209418 202046 209488 202102
rect 209168 201978 209488 202046
rect 209168 201922 209238 201978
rect 209294 201922 209362 201978
rect 209418 201922 209488 201978
rect 209168 201888 209488 201922
rect 239888 202350 240208 202384
rect 239888 202294 239958 202350
rect 240014 202294 240082 202350
rect 240138 202294 240208 202350
rect 239888 202226 240208 202294
rect 239888 202170 239958 202226
rect 240014 202170 240082 202226
rect 240138 202170 240208 202226
rect 239888 202102 240208 202170
rect 239888 202046 239958 202102
rect 240014 202046 240082 202102
rect 240138 202046 240208 202102
rect 239888 201978 240208 202046
rect 239888 201922 239958 201978
rect 240014 201922 240082 201978
rect 240138 201922 240208 201978
rect 239888 201888 240208 201922
rect 270608 202350 270928 202384
rect 270608 202294 270678 202350
rect 270734 202294 270802 202350
rect 270858 202294 270928 202350
rect 270608 202226 270928 202294
rect 270608 202170 270678 202226
rect 270734 202170 270802 202226
rect 270858 202170 270928 202226
rect 270608 202102 270928 202170
rect 270608 202046 270678 202102
rect 270734 202046 270802 202102
rect 270858 202046 270928 202102
rect 270608 201978 270928 202046
rect 270608 201922 270678 201978
rect 270734 201922 270802 201978
rect 270858 201922 270928 201978
rect 270608 201888 270928 201922
rect 193808 190350 194128 190384
rect 193808 190294 193878 190350
rect 193934 190294 194002 190350
rect 194058 190294 194128 190350
rect 193808 190226 194128 190294
rect 193808 190170 193878 190226
rect 193934 190170 194002 190226
rect 194058 190170 194128 190226
rect 193808 190102 194128 190170
rect 193808 190046 193878 190102
rect 193934 190046 194002 190102
rect 194058 190046 194128 190102
rect 193808 189978 194128 190046
rect 193808 189922 193878 189978
rect 193934 189922 194002 189978
rect 194058 189922 194128 189978
rect 193808 189888 194128 189922
rect 224528 190350 224848 190384
rect 224528 190294 224598 190350
rect 224654 190294 224722 190350
rect 224778 190294 224848 190350
rect 224528 190226 224848 190294
rect 224528 190170 224598 190226
rect 224654 190170 224722 190226
rect 224778 190170 224848 190226
rect 224528 190102 224848 190170
rect 224528 190046 224598 190102
rect 224654 190046 224722 190102
rect 224778 190046 224848 190102
rect 224528 189978 224848 190046
rect 224528 189922 224598 189978
rect 224654 189922 224722 189978
rect 224778 189922 224848 189978
rect 224528 189888 224848 189922
rect 255248 190350 255568 190384
rect 255248 190294 255318 190350
rect 255374 190294 255442 190350
rect 255498 190294 255568 190350
rect 255248 190226 255568 190294
rect 255248 190170 255318 190226
rect 255374 190170 255442 190226
rect 255498 190170 255568 190226
rect 255248 190102 255568 190170
rect 255248 190046 255318 190102
rect 255374 190046 255442 190102
rect 255498 190046 255568 190102
rect 255248 189978 255568 190046
rect 255248 189922 255318 189978
rect 255374 189922 255442 189978
rect 255498 189922 255568 189978
rect 255248 189888 255568 189922
rect 178448 184350 178768 184384
rect 178448 184294 178518 184350
rect 178574 184294 178642 184350
rect 178698 184294 178768 184350
rect 178448 184226 178768 184294
rect 178448 184170 178518 184226
rect 178574 184170 178642 184226
rect 178698 184170 178768 184226
rect 178448 184102 178768 184170
rect 178448 184046 178518 184102
rect 178574 184046 178642 184102
rect 178698 184046 178768 184102
rect 178448 183978 178768 184046
rect 178448 183922 178518 183978
rect 178574 183922 178642 183978
rect 178698 183922 178768 183978
rect 178448 183888 178768 183922
rect 209168 184350 209488 184384
rect 209168 184294 209238 184350
rect 209294 184294 209362 184350
rect 209418 184294 209488 184350
rect 209168 184226 209488 184294
rect 209168 184170 209238 184226
rect 209294 184170 209362 184226
rect 209418 184170 209488 184226
rect 209168 184102 209488 184170
rect 209168 184046 209238 184102
rect 209294 184046 209362 184102
rect 209418 184046 209488 184102
rect 209168 183978 209488 184046
rect 209168 183922 209238 183978
rect 209294 183922 209362 183978
rect 209418 183922 209488 183978
rect 209168 183888 209488 183922
rect 239888 184350 240208 184384
rect 239888 184294 239958 184350
rect 240014 184294 240082 184350
rect 240138 184294 240208 184350
rect 239888 184226 240208 184294
rect 239888 184170 239958 184226
rect 240014 184170 240082 184226
rect 240138 184170 240208 184226
rect 239888 184102 240208 184170
rect 239888 184046 239958 184102
rect 240014 184046 240082 184102
rect 240138 184046 240208 184102
rect 239888 183978 240208 184046
rect 239888 183922 239958 183978
rect 240014 183922 240082 183978
rect 240138 183922 240208 183978
rect 239888 183888 240208 183922
rect 270608 184350 270928 184384
rect 270608 184294 270678 184350
rect 270734 184294 270802 184350
rect 270858 184294 270928 184350
rect 270608 184226 270928 184294
rect 270608 184170 270678 184226
rect 270734 184170 270802 184226
rect 270858 184170 270928 184226
rect 270608 184102 270928 184170
rect 270608 184046 270678 184102
rect 270734 184046 270802 184102
rect 270858 184046 270928 184102
rect 270608 183978 270928 184046
rect 270608 183922 270678 183978
rect 270734 183922 270802 183978
rect 270858 183922 270928 183978
rect 270608 183888 270928 183922
rect 193808 172350 194128 172384
rect 193808 172294 193878 172350
rect 193934 172294 194002 172350
rect 194058 172294 194128 172350
rect 193808 172226 194128 172294
rect 193808 172170 193878 172226
rect 193934 172170 194002 172226
rect 194058 172170 194128 172226
rect 193808 172102 194128 172170
rect 193808 172046 193878 172102
rect 193934 172046 194002 172102
rect 194058 172046 194128 172102
rect 193808 171978 194128 172046
rect 193808 171922 193878 171978
rect 193934 171922 194002 171978
rect 194058 171922 194128 171978
rect 193808 171888 194128 171922
rect 224528 172350 224848 172384
rect 224528 172294 224598 172350
rect 224654 172294 224722 172350
rect 224778 172294 224848 172350
rect 224528 172226 224848 172294
rect 224528 172170 224598 172226
rect 224654 172170 224722 172226
rect 224778 172170 224848 172226
rect 224528 172102 224848 172170
rect 224528 172046 224598 172102
rect 224654 172046 224722 172102
rect 224778 172046 224848 172102
rect 224528 171978 224848 172046
rect 224528 171922 224598 171978
rect 224654 171922 224722 171978
rect 224778 171922 224848 171978
rect 224528 171888 224848 171922
rect 255248 172350 255568 172384
rect 255248 172294 255318 172350
rect 255374 172294 255442 172350
rect 255498 172294 255568 172350
rect 255248 172226 255568 172294
rect 255248 172170 255318 172226
rect 255374 172170 255442 172226
rect 255498 172170 255568 172226
rect 255248 172102 255568 172170
rect 255248 172046 255318 172102
rect 255374 172046 255442 172102
rect 255498 172046 255568 172102
rect 255248 171978 255568 172046
rect 255248 171922 255318 171978
rect 255374 171922 255442 171978
rect 255498 171922 255568 171978
rect 255248 171888 255568 171922
rect 178448 166350 178768 166384
rect 178448 166294 178518 166350
rect 178574 166294 178642 166350
rect 178698 166294 178768 166350
rect 178448 166226 178768 166294
rect 178448 166170 178518 166226
rect 178574 166170 178642 166226
rect 178698 166170 178768 166226
rect 178448 166102 178768 166170
rect 178448 166046 178518 166102
rect 178574 166046 178642 166102
rect 178698 166046 178768 166102
rect 178448 165978 178768 166046
rect 178448 165922 178518 165978
rect 178574 165922 178642 165978
rect 178698 165922 178768 165978
rect 178448 165888 178768 165922
rect 209168 166350 209488 166384
rect 209168 166294 209238 166350
rect 209294 166294 209362 166350
rect 209418 166294 209488 166350
rect 209168 166226 209488 166294
rect 209168 166170 209238 166226
rect 209294 166170 209362 166226
rect 209418 166170 209488 166226
rect 209168 166102 209488 166170
rect 209168 166046 209238 166102
rect 209294 166046 209362 166102
rect 209418 166046 209488 166102
rect 209168 165978 209488 166046
rect 209168 165922 209238 165978
rect 209294 165922 209362 165978
rect 209418 165922 209488 165978
rect 209168 165888 209488 165922
rect 239888 166350 240208 166384
rect 239888 166294 239958 166350
rect 240014 166294 240082 166350
rect 240138 166294 240208 166350
rect 239888 166226 240208 166294
rect 239888 166170 239958 166226
rect 240014 166170 240082 166226
rect 240138 166170 240208 166226
rect 239888 166102 240208 166170
rect 239888 166046 239958 166102
rect 240014 166046 240082 166102
rect 240138 166046 240208 166102
rect 239888 165978 240208 166046
rect 239888 165922 239958 165978
rect 240014 165922 240082 165978
rect 240138 165922 240208 165978
rect 239888 165888 240208 165922
rect 270608 166350 270928 166384
rect 270608 166294 270678 166350
rect 270734 166294 270802 166350
rect 270858 166294 270928 166350
rect 270608 166226 270928 166294
rect 270608 166170 270678 166226
rect 270734 166170 270802 166226
rect 270858 166170 270928 166226
rect 270608 166102 270928 166170
rect 270608 166046 270678 166102
rect 270734 166046 270802 166102
rect 270858 166046 270928 166102
rect 270608 165978 270928 166046
rect 270608 165922 270678 165978
rect 270734 165922 270802 165978
rect 270858 165922 270928 165978
rect 270608 165888 270928 165922
rect 174076 157378 174132 157388
rect 193808 154350 194128 154384
rect 193808 154294 193878 154350
rect 193934 154294 194002 154350
rect 194058 154294 194128 154350
rect 193808 154226 194128 154294
rect 193808 154170 193878 154226
rect 193934 154170 194002 154226
rect 194058 154170 194128 154226
rect 193808 154102 194128 154170
rect 193808 154046 193878 154102
rect 193934 154046 194002 154102
rect 194058 154046 194128 154102
rect 193808 153978 194128 154046
rect 193808 153922 193878 153978
rect 193934 153922 194002 153978
rect 194058 153922 194128 153978
rect 193808 153888 194128 153922
rect 224528 154350 224848 154384
rect 224528 154294 224598 154350
rect 224654 154294 224722 154350
rect 224778 154294 224848 154350
rect 224528 154226 224848 154294
rect 224528 154170 224598 154226
rect 224654 154170 224722 154226
rect 224778 154170 224848 154226
rect 224528 154102 224848 154170
rect 224528 154046 224598 154102
rect 224654 154046 224722 154102
rect 224778 154046 224848 154102
rect 224528 153978 224848 154046
rect 224528 153922 224598 153978
rect 224654 153922 224722 153978
rect 224778 153922 224848 153978
rect 224528 153888 224848 153922
rect 255248 154350 255568 154384
rect 255248 154294 255318 154350
rect 255374 154294 255442 154350
rect 255498 154294 255568 154350
rect 255248 154226 255568 154294
rect 255248 154170 255318 154226
rect 255374 154170 255442 154226
rect 255498 154170 255568 154226
rect 255248 154102 255568 154170
rect 255248 154046 255318 154102
rect 255374 154046 255442 154102
rect 255498 154046 255568 154102
rect 255248 153978 255568 154046
rect 255248 153922 255318 153978
rect 255374 153922 255442 153978
rect 255498 153922 255568 153978
rect 255248 153888 255568 153922
rect 178448 148350 178768 148384
rect 178448 148294 178518 148350
rect 178574 148294 178642 148350
rect 178698 148294 178768 148350
rect 178448 148226 178768 148294
rect 178448 148170 178518 148226
rect 178574 148170 178642 148226
rect 178698 148170 178768 148226
rect 178448 148102 178768 148170
rect 178448 148046 178518 148102
rect 178574 148046 178642 148102
rect 178698 148046 178768 148102
rect 178448 147978 178768 148046
rect 178448 147922 178518 147978
rect 178574 147922 178642 147978
rect 178698 147922 178768 147978
rect 178448 147888 178768 147922
rect 209168 148350 209488 148384
rect 209168 148294 209238 148350
rect 209294 148294 209362 148350
rect 209418 148294 209488 148350
rect 209168 148226 209488 148294
rect 209168 148170 209238 148226
rect 209294 148170 209362 148226
rect 209418 148170 209488 148226
rect 209168 148102 209488 148170
rect 209168 148046 209238 148102
rect 209294 148046 209362 148102
rect 209418 148046 209488 148102
rect 209168 147978 209488 148046
rect 209168 147922 209238 147978
rect 209294 147922 209362 147978
rect 209418 147922 209488 147978
rect 209168 147888 209488 147922
rect 239888 148350 240208 148384
rect 239888 148294 239958 148350
rect 240014 148294 240082 148350
rect 240138 148294 240208 148350
rect 239888 148226 240208 148294
rect 239888 148170 239958 148226
rect 240014 148170 240082 148226
rect 240138 148170 240208 148226
rect 239888 148102 240208 148170
rect 239888 148046 239958 148102
rect 240014 148046 240082 148102
rect 240138 148046 240208 148102
rect 239888 147978 240208 148046
rect 239888 147922 239958 147978
rect 240014 147922 240082 147978
rect 240138 147922 240208 147978
rect 239888 147888 240208 147922
rect 270608 148350 270928 148384
rect 270608 148294 270678 148350
rect 270734 148294 270802 148350
rect 270858 148294 270928 148350
rect 270608 148226 270928 148294
rect 270608 148170 270678 148226
rect 270734 148170 270802 148226
rect 270858 148170 270928 148226
rect 270608 148102 270928 148170
rect 270608 148046 270678 148102
rect 270734 148046 270802 148102
rect 270858 148046 270928 148102
rect 270608 147978 270928 148046
rect 270608 147922 270678 147978
rect 270734 147922 270802 147978
rect 270858 147922 270928 147978
rect 270608 147888 270928 147922
rect 193808 136350 194128 136384
rect 193808 136294 193878 136350
rect 193934 136294 194002 136350
rect 194058 136294 194128 136350
rect 193808 136226 194128 136294
rect 193808 136170 193878 136226
rect 193934 136170 194002 136226
rect 194058 136170 194128 136226
rect 193808 136102 194128 136170
rect 193808 136046 193878 136102
rect 193934 136046 194002 136102
rect 194058 136046 194128 136102
rect 193808 135978 194128 136046
rect 193808 135922 193878 135978
rect 193934 135922 194002 135978
rect 194058 135922 194128 135978
rect 193808 135888 194128 135922
rect 224528 136350 224848 136384
rect 224528 136294 224598 136350
rect 224654 136294 224722 136350
rect 224778 136294 224848 136350
rect 224528 136226 224848 136294
rect 224528 136170 224598 136226
rect 224654 136170 224722 136226
rect 224778 136170 224848 136226
rect 224528 136102 224848 136170
rect 224528 136046 224598 136102
rect 224654 136046 224722 136102
rect 224778 136046 224848 136102
rect 224528 135978 224848 136046
rect 224528 135922 224598 135978
rect 224654 135922 224722 135978
rect 224778 135922 224848 135978
rect 224528 135888 224848 135922
rect 255248 136350 255568 136384
rect 255248 136294 255318 136350
rect 255374 136294 255442 136350
rect 255498 136294 255568 136350
rect 255248 136226 255568 136294
rect 255248 136170 255318 136226
rect 255374 136170 255442 136226
rect 255498 136170 255568 136226
rect 255248 136102 255568 136170
rect 255248 136046 255318 136102
rect 255374 136046 255442 136102
rect 255498 136046 255568 136102
rect 255248 135978 255568 136046
rect 255248 135922 255318 135978
rect 255374 135922 255442 135978
rect 255498 135922 255568 135978
rect 255248 135888 255568 135922
rect 178448 130350 178768 130384
rect 178448 130294 178518 130350
rect 178574 130294 178642 130350
rect 178698 130294 178768 130350
rect 178448 130226 178768 130294
rect 178448 130170 178518 130226
rect 178574 130170 178642 130226
rect 178698 130170 178768 130226
rect 178448 130102 178768 130170
rect 178448 130046 178518 130102
rect 178574 130046 178642 130102
rect 178698 130046 178768 130102
rect 178448 129978 178768 130046
rect 178448 129922 178518 129978
rect 178574 129922 178642 129978
rect 178698 129922 178768 129978
rect 178448 129888 178768 129922
rect 209168 130350 209488 130384
rect 209168 130294 209238 130350
rect 209294 130294 209362 130350
rect 209418 130294 209488 130350
rect 209168 130226 209488 130294
rect 209168 130170 209238 130226
rect 209294 130170 209362 130226
rect 209418 130170 209488 130226
rect 209168 130102 209488 130170
rect 209168 130046 209238 130102
rect 209294 130046 209362 130102
rect 209418 130046 209488 130102
rect 209168 129978 209488 130046
rect 209168 129922 209238 129978
rect 209294 129922 209362 129978
rect 209418 129922 209488 129978
rect 209168 129888 209488 129922
rect 239888 130350 240208 130384
rect 239888 130294 239958 130350
rect 240014 130294 240082 130350
rect 240138 130294 240208 130350
rect 239888 130226 240208 130294
rect 239888 130170 239958 130226
rect 240014 130170 240082 130226
rect 240138 130170 240208 130226
rect 239888 130102 240208 130170
rect 239888 130046 239958 130102
rect 240014 130046 240082 130102
rect 240138 130046 240208 130102
rect 239888 129978 240208 130046
rect 239888 129922 239958 129978
rect 240014 129922 240082 129978
rect 240138 129922 240208 129978
rect 239888 129888 240208 129922
rect 270608 130350 270928 130384
rect 270608 130294 270678 130350
rect 270734 130294 270802 130350
rect 270858 130294 270928 130350
rect 270608 130226 270928 130294
rect 270608 130170 270678 130226
rect 270734 130170 270802 130226
rect 270858 130170 270928 130226
rect 270608 130102 270928 130170
rect 270608 130046 270678 130102
rect 270734 130046 270802 130102
rect 270858 130046 270928 130102
rect 270608 129978 270928 130046
rect 270608 129922 270678 129978
rect 270734 129922 270802 129978
rect 270858 129922 270928 129978
rect 270608 129888 270928 129922
rect 193808 118350 194128 118384
rect 193808 118294 193878 118350
rect 193934 118294 194002 118350
rect 194058 118294 194128 118350
rect 193808 118226 194128 118294
rect 193808 118170 193878 118226
rect 193934 118170 194002 118226
rect 194058 118170 194128 118226
rect 193808 118102 194128 118170
rect 193808 118046 193878 118102
rect 193934 118046 194002 118102
rect 194058 118046 194128 118102
rect 193808 117978 194128 118046
rect 193808 117922 193878 117978
rect 193934 117922 194002 117978
rect 194058 117922 194128 117978
rect 193808 117888 194128 117922
rect 224528 118350 224848 118384
rect 224528 118294 224598 118350
rect 224654 118294 224722 118350
rect 224778 118294 224848 118350
rect 224528 118226 224848 118294
rect 224528 118170 224598 118226
rect 224654 118170 224722 118226
rect 224778 118170 224848 118226
rect 224528 118102 224848 118170
rect 224528 118046 224598 118102
rect 224654 118046 224722 118102
rect 224778 118046 224848 118102
rect 224528 117978 224848 118046
rect 224528 117922 224598 117978
rect 224654 117922 224722 117978
rect 224778 117922 224848 117978
rect 224528 117888 224848 117922
rect 255248 118350 255568 118384
rect 255248 118294 255318 118350
rect 255374 118294 255442 118350
rect 255498 118294 255568 118350
rect 255248 118226 255568 118294
rect 255248 118170 255318 118226
rect 255374 118170 255442 118226
rect 255498 118170 255568 118226
rect 255248 118102 255568 118170
rect 255248 118046 255318 118102
rect 255374 118046 255442 118102
rect 255498 118046 255568 118102
rect 255248 117978 255568 118046
rect 255248 117922 255318 117978
rect 255374 117922 255442 117978
rect 255498 117922 255568 117978
rect 255248 117888 255568 117922
rect 178448 112350 178768 112384
rect 178448 112294 178518 112350
rect 178574 112294 178642 112350
rect 178698 112294 178768 112350
rect 178448 112226 178768 112294
rect 178448 112170 178518 112226
rect 178574 112170 178642 112226
rect 178698 112170 178768 112226
rect 178448 112102 178768 112170
rect 178448 112046 178518 112102
rect 178574 112046 178642 112102
rect 178698 112046 178768 112102
rect 178448 111978 178768 112046
rect 178448 111922 178518 111978
rect 178574 111922 178642 111978
rect 178698 111922 178768 111978
rect 178448 111888 178768 111922
rect 209168 112350 209488 112384
rect 209168 112294 209238 112350
rect 209294 112294 209362 112350
rect 209418 112294 209488 112350
rect 209168 112226 209488 112294
rect 209168 112170 209238 112226
rect 209294 112170 209362 112226
rect 209418 112170 209488 112226
rect 209168 112102 209488 112170
rect 209168 112046 209238 112102
rect 209294 112046 209362 112102
rect 209418 112046 209488 112102
rect 209168 111978 209488 112046
rect 209168 111922 209238 111978
rect 209294 111922 209362 111978
rect 209418 111922 209488 111978
rect 209168 111888 209488 111922
rect 239888 112350 240208 112384
rect 239888 112294 239958 112350
rect 240014 112294 240082 112350
rect 240138 112294 240208 112350
rect 239888 112226 240208 112294
rect 239888 112170 239958 112226
rect 240014 112170 240082 112226
rect 240138 112170 240208 112226
rect 239888 112102 240208 112170
rect 239888 112046 239958 112102
rect 240014 112046 240082 112102
rect 240138 112046 240208 112102
rect 239888 111978 240208 112046
rect 239888 111922 239958 111978
rect 240014 111922 240082 111978
rect 240138 111922 240208 111978
rect 239888 111888 240208 111922
rect 270608 112350 270928 112384
rect 270608 112294 270678 112350
rect 270734 112294 270802 112350
rect 270858 112294 270928 112350
rect 270608 112226 270928 112294
rect 270608 112170 270678 112226
rect 270734 112170 270802 112226
rect 270858 112170 270928 112226
rect 270608 112102 270928 112170
rect 270608 112046 270678 112102
rect 270734 112046 270802 112102
rect 270858 112046 270928 112102
rect 270608 111978 270928 112046
rect 270608 111922 270678 111978
rect 270734 111922 270802 111978
rect 270858 111922 270928 111978
rect 270608 111888 270928 111922
rect 271516 108298 271572 108308
rect 174636 105252 174692 105262
rect 174692 105196 174804 105238
rect 174636 105182 174804 105196
rect 174748 99540 174804 105182
rect 174748 99474 174804 99484
rect 189738 94350 190358 104970
rect 189738 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 190358 94350
rect 189738 94226 190358 94294
rect 189738 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 190358 94226
rect 189738 94102 190358 94170
rect 189738 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 190358 94102
rect 189738 93978 190358 94046
rect 189738 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 190358 93978
rect 189532 86518 189588 86528
rect 181468 81478 181524 81488
rect 181468 80276 181524 81422
rect 189532 80612 189588 86462
rect 189532 80546 189588 80556
rect 181468 80210 181524 80220
rect 173852 78978 173908 78988
rect 189738 76350 190358 93922
rect 189738 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 190358 76350
rect 189738 76226 190358 76294
rect 189738 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 190358 76226
rect 189738 76102 190358 76170
rect 189738 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 190358 76102
rect 189738 75978 190358 76046
rect 189738 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 190358 75978
rect 189738 74766 190358 75922
rect 193458 99923 194078 99964
rect 193458 99867 193554 99923
rect 193610 99867 193678 99923
rect 193734 99867 193802 99923
rect 193858 99867 193926 99923
rect 193982 99867 194078 99923
rect 193458 82350 194078 99867
rect 220458 94350 221078 104970
rect 243516 101998 243572 102008
rect 226604 101818 226660 101828
rect 220458 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 221078 94350
rect 220458 94226 221078 94294
rect 220458 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 221078 94226
rect 220458 94102 221078 94170
rect 220458 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 221078 94102
rect 220458 93978 221078 94046
rect 220458 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 221078 93978
rect 206556 88498 206612 88508
rect 193458 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 194078 82350
rect 193458 82226 194078 82294
rect 193458 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 194078 82226
rect 193458 82102 194078 82170
rect 193458 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 194078 82102
rect 193458 81978 194078 82046
rect 193458 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 194078 81978
rect 193458 74766 194078 81922
rect 202524 88318 202580 88328
rect 202524 80612 202580 88262
rect 202524 80546 202580 80556
rect 204876 88138 204932 88148
rect 204876 80612 204932 88082
rect 204876 80546 204932 80556
rect 206556 80612 206612 88442
rect 206556 80546 206612 80556
rect 213948 85078 214004 85088
rect 213948 80612 214004 85022
rect 213948 80546 214004 80556
rect 214844 84898 214900 84908
rect 214844 80612 214900 84842
rect 214844 80546 214900 80556
rect 220458 76350 221078 93922
rect 220458 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 221078 76350
rect 220458 76226 221078 76294
rect 220458 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 221078 76226
rect 220458 76102 221078 76170
rect 220458 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 221078 76102
rect 220458 75978 221078 76046
rect 220458 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 221078 75978
rect 220458 74766 221078 75922
rect 224178 99923 224798 99964
rect 224178 99867 224274 99923
rect 224330 99867 224398 99923
rect 224454 99867 224522 99923
rect 224578 99867 224646 99923
rect 224702 99867 224798 99923
rect 224178 82350 224798 99867
rect 224178 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 224798 82350
rect 224178 82226 224798 82294
rect 224178 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 224798 82226
rect 224178 82102 224798 82170
rect 224178 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 224798 82102
rect 224178 81978 224798 82046
rect 224178 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 224798 81978
rect 224178 74766 224798 81922
rect 226604 80612 226660 101762
rect 226604 80546 226660 80556
rect 226716 101638 226772 101648
rect 226716 80500 226772 101582
rect 235116 98578 235172 98588
rect 233436 98398 233492 98408
rect 230076 98218 230132 98228
rect 228396 96598 228452 96608
rect 228396 80612 228452 96542
rect 228396 80546 228452 80556
rect 229964 92458 230020 92468
rect 229964 80612 230020 92402
rect 229964 80546 230020 80556
rect 226716 80434 226772 80444
rect 230076 80500 230132 98162
rect 232092 89938 232148 89948
rect 232092 80612 232148 89882
rect 232092 80546 232148 80556
rect 233436 80612 233492 98342
rect 235116 80612 235172 98522
rect 241836 96778 241892 96788
rect 233436 80546 233492 80556
rect 234780 80578 234836 80588
rect 230076 80434 230132 80444
rect 235116 80546 235172 80556
rect 236796 94978 236852 94988
rect 236796 80612 236852 94922
rect 236796 80546 236852 80556
rect 238476 93178 238532 93188
rect 238476 80612 238532 93122
rect 238476 80546 238532 80556
rect 241836 80612 241892 96722
rect 241836 80546 241892 80556
rect 243516 80612 243572 101942
rect 251178 94350 251798 104970
rect 267932 104158 267988 104168
rect 251178 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 251798 94350
rect 251178 94226 251798 94294
rect 251178 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 251798 94226
rect 251178 94102 251798 94170
rect 251178 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 251798 94102
rect 251178 93978 251798 94046
rect 251178 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 251798 93978
rect 243516 80546 243572 80556
rect 245196 91558 245252 91568
rect 245196 80612 245252 91502
rect 249564 89218 249620 89228
rect 245196 80546 245252 80556
rect 246876 87418 246932 87428
rect 246876 80612 246932 87362
rect 246876 80546 246932 80556
rect 249564 80612 249620 89162
rect 249564 80546 249620 80556
rect 229964 80398 230020 80408
rect 229964 79716 230020 80342
rect 231420 80218 231476 80228
rect 229964 79650 230020 79660
rect 230748 79858 230804 79868
rect 230748 79380 230804 79802
rect 231420 79604 231476 80162
rect 231420 79538 231476 79548
rect 232764 80038 232820 80048
rect 232764 79492 232820 79982
rect 234780 79828 234836 80522
rect 234780 79762 234836 79772
rect 232764 79426 232820 79436
rect 230748 79314 230804 79324
rect 227388 79044 227444 79054
rect 227276 78958 227444 78988
rect 227332 78932 227444 78958
rect 227276 78892 227332 78902
rect 250908 78058 250964 78068
rect 250908 77364 250964 78002
rect 250908 77298 250964 77308
rect 251178 76350 251798 93922
rect 254898 99923 255518 99964
rect 254898 99867 254994 99923
rect 255050 99867 255118 99923
rect 255174 99867 255242 99923
rect 255298 99867 255366 99923
rect 255422 99867 255518 99923
rect 254716 91198 254772 91208
rect 253484 91018 253540 91028
rect 251916 90838 251972 90848
rect 251916 80612 251972 90782
rect 251916 80546 251972 80556
rect 252924 80938 252980 80948
rect 252924 79716 252980 80882
rect 253484 80612 253540 90962
rect 253484 80546 253540 80556
rect 254492 82738 254548 82748
rect 254492 80500 254548 82682
rect 254716 80612 254772 91142
rect 254716 80546 254772 80556
rect 254898 82350 255518 99867
rect 266476 97748 266532 97758
rect 266252 97636 266308 97646
rect 254898 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 255518 82350
rect 254898 82226 255518 82294
rect 254898 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 255518 82226
rect 254898 82102 255518 82170
rect 254898 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 255518 82102
rect 254898 81978 255518 82046
rect 254898 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 255518 81978
rect 254492 80434 254548 80444
rect 252924 79650 252980 79660
rect 251178 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 251798 76350
rect 251178 76226 251798 76294
rect 251178 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 251798 76226
rect 251178 76102 251798 76170
rect 251178 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 251798 76102
rect 251178 75978 251798 76046
rect 251178 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 251798 75978
rect 251178 74766 251798 75922
rect 254898 74766 255518 81922
rect 259644 89398 259700 89408
rect 256956 80758 257012 80768
rect 256956 79716 257012 80702
rect 259644 80612 259700 89342
rect 259644 80546 259700 80556
rect 265244 87780 265300 87790
rect 256956 79650 257012 79660
rect 169708 73938 169764 73948
rect 185808 64350 186128 64384
rect 185808 64294 185878 64350
rect 185934 64294 186002 64350
rect 186058 64294 186128 64350
rect 185808 64226 186128 64294
rect 185808 64170 185878 64226
rect 185934 64170 186002 64226
rect 186058 64170 186128 64226
rect 185808 64102 186128 64170
rect 185808 64046 185878 64102
rect 185934 64046 186002 64102
rect 186058 64046 186128 64102
rect 185808 63978 186128 64046
rect 185808 63922 185878 63978
rect 185934 63922 186002 63978
rect 186058 63922 186128 63978
rect 185808 63888 186128 63922
rect 216528 64350 216848 64384
rect 216528 64294 216598 64350
rect 216654 64294 216722 64350
rect 216778 64294 216848 64350
rect 216528 64226 216848 64294
rect 216528 64170 216598 64226
rect 216654 64170 216722 64226
rect 216778 64170 216848 64226
rect 216528 64102 216848 64170
rect 216528 64046 216598 64102
rect 216654 64046 216722 64102
rect 216778 64046 216848 64102
rect 216528 63978 216848 64046
rect 216528 63922 216598 63978
rect 216654 63922 216722 63978
rect 216778 63922 216848 63978
rect 216528 63888 216848 63922
rect 247248 64350 247568 64384
rect 247248 64294 247318 64350
rect 247374 64294 247442 64350
rect 247498 64294 247568 64350
rect 247248 64226 247568 64294
rect 247248 64170 247318 64226
rect 247374 64170 247442 64226
rect 247498 64170 247568 64226
rect 247248 64102 247568 64170
rect 247248 64046 247318 64102
rect 247374 64046 247442 64102
rect 247498 64046 247568 64102
rect 247248 63978 247568 64046
rect 247248 63922 247318 63978
rect 247374 63922 247442 63978
rect 247498 63922 247568 63978
rect 247248 63888 247568 63922
rect 170448 58350 170768 58384
rect 170448 58294 170518 58350
rect 170574 58294 170642 58350
rect 170698 58294 170768 58350
rect 170448 58226 170768 58294
rect 170448 58170 170518 58226
rect 170574 58170 170642 58226
rect 170698 58170 170768 58226
rect 170448 58102 170768 58170
rect 170448 58046 170518 58102
rect 170574 58046 170642 58102
rect 170698 58046 170768 58102
rect 170448 57978 170768 58046
rect 170448 57922 170518 57978
rect 170574 57922 170642 57978
rect 170698 57922 170768 57978
rect 170448 57888 170768 57922
rect 201168 58350 201488 58384
rect 201168 58294 201238 58350
rect 201294 58294 201362 58350
rect 201418 58294 201488 58350
rect 201168 58226 201488 58294
rect 201168 58170 201238 58226
rect 201294 58170 201362 58226
rect 201418 58170 201488 58226
rect 201168 58102 201488 58170
rect 201168 58046 201238 58102
rect 201294 58046 201362 58102
rect 201418 58046 201488 58102
rect 201168 57978 201488 58046
rect 201168 57922 201238 57978
rect 201294 57922 201362 57978
rect 201418 57922 201488 57978
rect 201168 57888 201488 57922
rect 231888 58350 232208 58384
rect 231888 58294 231958 58350
rect 232014 58294 232082 58350
rect 232138 58294 232208 58350
rect 231888 58226 232208 58294
rect 231888 58170 231958 58226
rect 232014 58170 232082 58226
rect 232138 58170 232208 58226
rect 231888 58102 232208 58170
rect 231888 58046 231958 58102
rect 232014 58046 232082 58102
rect 232138 58046 232208 58102
rect 231888 57978 232208 58046
rect 231888 57922 231958 57978
rect 232014 57922 232082 57978
rect 232138 57922 232208 57978
rect 231888 57888 232208 57922
rect 262608 58350 262928 58384
rect 262608 58294 262678 58350
rect 262734 58294 262802 58350
rect 262858 58294 262928 58350
rect 262608 58226 262928 58294
rect 262608 58170 262678 58226
rect 262734 58170 262802 58226
rect 262858 58170 262928 58226
rect 262608 58102 262928 58170
rect 262608 58046 262678 58102
rect 262734 58046 262802 58102
rect 262858 58046 262928 58102
rect 262608 57978 262928 58046
rect 262608 57922 262678 57978
rect 262734 57922 262802 57978
rect 262858 57922 262928 57978
rect 262608 57888 262928 57922
rect 264572 54658 264628 54668
rect 185808 46350 186128 46384
rect 185808 46294 185878 46350
rect 185934 46294 186002 46350
rect 186058 46294 186128 46350
rect 185808 46226 186128 46294
rect 185808 46170 185878 46226
rect 185934 46170 186002 46226
rect 186058 46170 186128 46226
rect 185808 46102 186128 46170
rect 185808 46046 185878 46102
rect 185934 46046 186002 46102
rect 186058 46046 186128 46102
rect 185808 45978 186128 46046
rect 185808 45922 185878 45978
rect 185934 45922 186002 45978
rect 186058 45922 186128 45978
rect 185808 45888 186128 45922
rect 216528 46350 216848 46384
rect 216528 46294 216598 46350
rect 216654 46294 216722 46350
rect 216778 46294 216848 46350
rect 216528 46226 216848 46294
rect 216528 46170 216598 46226
rect 216654 46170 216722 46226
rect 216778 46170 216848 46226
rect 216528 46102 216848 46170
rect 216528 46046 216598 46102
rect 216654 46046 216722 46102
rect 216778 46046 216848 46102
rect 216528 45978 216848 46046
rect 216528 45922 216598 45978
rect 216654 45922 216722 45978
rect 216778 45922 216848 45978
rect 216528 45888 216848 45922
rect 247248 46350 247568 46384
rect 247248 46294 247318 46350
rect 247374 46294 247442 46350
rect 247498 46294 247568 46350
rect 247248 46226 247568 46294
rect 247248 46170 247318 46226
rect 247374 46170 247442 46226
rect 247498 46170 247568 46226
rect 247248 46102 247568 46170
rect 247248 46046 247318 46102
rect 247374 46046 247442 46102
rect 247498 46046 247568 46102
rect 247248 45978 247568 46046
rect 247248 45922 247318 45978
rect 247374 45922 247442 45978
rect 247498 45922 247568 45978
rect 247248 45888 247568 45922
rect 170448 40350 170768 40384
rect 170448 40294 170518 40350
rect 170574 40294 170642 40350
rect 170698 40294 170768 40350
rect 170448 40226 170768 40294
rect 170448 40170 170518 40226
rect 170574 40170 170642 40226
rect 170698 40170 170768 40226
rect 170448 40102 170768 40170
rect 170448 40046 170518 40102
rect 170574 40046 170642 40102
rect 170698 40046 170768 40102
rect 170448 39978 170768 40046
rect 170448 39922 170518 39978
rect 170574 39922 170642 39978
rect 170698 39922 170768 39978
rect 170448 39888 170768 39922
rect 201168 40350 201488 40384
rect 201168 40294 201238 40350
rect 201294 40294 201362 40350
rect 201418 40294 201488 40350
rect 201168 40226 201488 40294
rect 201168 40170 201238 40226
rect 201294 40170 201362 40226
rect 201418 40170 201488 40226
rect 201168 40102 201488 40170
rect 201168 40046 201238 40102
rect 201294 40046 201362 40102
rect 201418 40046 201488 40102
rect 201168 39978 201488 40046
rect 201168 39922 201238 39978
rect 201294 39922 201362 39978
rect 201418 39922 201488 39978
rect 201168 39888 201488 39922
rect 231888 40350 232208 40384
rect 231888 40294 231958 40350
rect 232014 40294 232082 40350
rect 232138 40294 232208 40350
rect 231888 40226 232208 40294
rect 231888 40170 231958 40226
rect 232014 40170 232082 40226
rect 232138 40170 232208 40226
rect 231888 40102 232208 40170
rect 231888 40046 231958 40102
rect 232014 40046 232082 40102
rect 232138 40046 232208 40102
rect 231888 39978 232208 40046
rect 231888 39922 231958 39978
rect 232014 39922 232082 39978
rect 232138 39922 232208 39978
rect 231888 39888 232208 39922
rect 262608 40350 262928 40384
rect 262608 40294 262678 40350
rect 262734 40294 262802 40350
rect 262858 40294 262928 40350
rect 262608 40226 262928 40294
rect 262608 40170 262678 40226
rect 262734 40170 262802 40226
rect 262858 40170 262928 40226
rect 262608 40102 262928 40170
rect 262608 40046 262678 40102
rect 262734 40046 262802 40102
rect 262858 40046 262928 40102
rect 262608 39978 262928 40046
rect 262608 39922 262678 39978
rect 262734 39922 262802 39978
rect 262858 39922 262928 39978
rect 262608 39888 262928 39922
rect 185808 28350 186128 28384
rect 185808 28294 185878 28350
rect 185934 28294 186002 28350
rect 186058 28294 186128 28350
rect 185808 28226 186128 28294
rect 185808 28170 185878 28226
rect 185934 28170 186002 28226
rect 186058 28170 186128 28226
rect 185808 28102 186128 28170
rect 185808 28046 185878 28102
rect 185934 28046 186002 28102
rect 186058 28046 186128 28102
rect 185808 27978 186128 28046
rect 185808 27922 185878 27978
rect 185934 27922 186002 27978
rect 186058 27922 186128 27978
rect 185808 27888 186128 27922
rect 216528 28350 216848 28384
rect 216528 28294 216598 28350
rect 216654 28294 216722 28350
rect 216778 28294 216848 28350
rect 216528 28226 216848 28294
rect 216528 28170 216598 28226
rect 216654 28170 216722 28226
rect 216778 28170 216848 28226
rect 216528 28102 216848 28170
rect 216528 28046 216598 28102
rect 216654 28046 216722 28102
rect 216778 28046 216848 28102
rect 216528 27978 216848 28046
rect 216528 27922 216598 27978
rect 216654 27922 216722 27978
rect 216778 27922 216848 27978
rect 216528 27888 216848 27922
rect 247248 28350 247568 28384
rect 247248 28294 247318 28350
rect 247374 28294 247442 28350
rect 247498 28294 247568 28350
rect 247248 28226 247568 28294
rect 247248 28170 247318 28226
rect 247374 28170 247442 28226
rect 247498 28170 247568 28226
rect 247248 28102 247568 28170
rect 247248 28046 247318 28102
rect 247374 28046 247442 28102
rect 247498 28046 247568 28102
rect 247248 27978 247568 28046
rect 247248 27922 247318 27978
rect 247374 27922 247442 27978
rect 247498 27922 247568 27978
rect 247248 27888 247568 27922
rect 170448 22350 170768 22384
rect 170448 22294 170518 22350
rect 170574 22294 170642 22350
rect 170698 22294 170768 22350
rect 170448 22226 170768 22294
rect 170448 22170 170518 22226
rect 170574 22170 170642 22226
rect 170698 22170 170768 22226
rect 170448 22102 170768 22170
rect 170448 22046 170518 22102
rect 170574 22046 170642 22102
rect 170698 22046 170768 22102
rect 170448 21978 170768 22046
rect 170448 21922 170518 21978
rect 170574 21922 170642 21978
rect 170698 21922 170768 21978
rect 170448 21888 170768 21922
rect 201168 22350 201488 22384
rect 201168 22294 201238 22350
rect 201294 22294 201362 22350
rect 201418 22294 201488 22350
rect 201168 22226 201488 22294
rect 201168 22170 201238 22226
rect 201294 22170 201362 22226
rect 201418 22170 201488 22226
rect 201168 22102 201488 22170
rect 201168 22046 201238 22102
rect 201294 22046 201362 22102
rect 201418 22046 201488 22102
rect 201168 21978 201488 22046
rect 201168 21922 201238 21978
rect 201294 21922 201362 21978
rect 201418 21922 201488 21978
rect 201168 21888 201488 21922
rect 231888 22350 232208 22384
rect 231888 22294 231958 22350
rect 232014 22294 232082 22350
rect 232138 22294 232208 22350
rect 231888 22226 232208 22294
rect 231888 22170 231958 22226
rect 232014 22170 232082 22226
rect 232138 22170 232208 22226
rect 231888 22102 232208 22170
rect 231888 22046 231958 22102
rect 232014 22046 232082 22102
rect 232138 22046 232208 22102
rect 231888 21978 232208 22046
rect 231888 21922 231958 21978
rect 232014 21922 232082 21978
rect 232138 21922 232208 21978
rect 231888 21888 232208 21922
rect 262608 22350 262928 22384
rect 262608 22294 262678 22350
rect 262734 22294 262802 22350
rect 262858 22294 262928 22350
rect 262608 22226 262928 22294
rect 262608 22170 262678 22226
rect 262734 22170 262802 22226
rect 262858 22170 262928 22226
rect 262608 22102 262928 22170
rect 262608 22046 262678 22102
rect 262734 22046 262802 22102
rect 262858 22046 262928 22102
rect 262608 21978 262928 22046
rect 262608 21922 262678 21978
rect 262734 21922 262802 21978
rect 262858 21922 262928 21978
rect 262608 21888 262928 21922
rect 241948 21358 242004 21368
rect 240604 21178 240660 21188
rect 240380 20998 240436 21008
rect 231196 19918 231252 19928
rect 187068 13618 187124 13628
rect 169596 13372 169652 13382
rect 186844 13412 186900 13422
rect 185724 13078 185780 13086
rect 185724 13076 186340 13078
rect 185780 13022 186340 13076
rect 185724 13010 185780 13020
rect 186284 12898 186340 13022
rect 186284 12852 186452 12898
rect 186284 12842 186396 12852
rect 186396 12786 186452 12796
rect 185052 12516 185108 12526
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 184940 12292 184996 12302
rect 184940 5878 184996 12236
rect 184940 5812 184996 5822
rect 185052 3358 185108 12460
rect 186172 12292 186228 12302
rect 186172 9298 186228 12236
rect 186172 9232 186228 9242
rect 186508 12292 186564 12302
rect 186508 6058 186564 12236
rect 186844 11818 186900 13356
rect 187068 13412 187124 13562
rect 187068 13346 187124 13356
rect 186844 11752 186900 11762
rect 188188 12292 188244 12302
rect 188188 7498 188244 12236
rect 188188 7432 188244 7442
rect 186508 5992 186564 6002
rect 185052 3292 185108 3302
rect 189738 4350 190358 19842
rect 190428 13188 190484 13198
rect 190428 12538 190484 13132
rect 190428 12482 190596 12538
rect 190428 12292 190484 12302
rect 190428 7678 190484 12236
rect 190540 11998 190596 12482
rect 190540 11932 190596 11942
rect 190428 7612 190484 7622
rect 193458 10350 194078 19842
rect 219548 17220 219604 17230
rect 219548 16884 219604 17164
rect 219548 16818 219604 16828
rect 217308 16138 217364 16148
rect 217308 16034 217364 16044
rect 218652 13618 218708 13628
rect 209692 13438 209748 13450
rect 209468 13412 209524 13422
rect 209468 13078 209524 13356
rect 210140 13438 210196 13450
rect 209692 13346 209748 13356
rect 209916 13412 209972 13422
rect 209916 13258 209972 13356
rect 210140 13346 210196 13356
rect 218652 13412 218708 13562
rect 218652 13346 218708 13356
rect 209916 13192 209972 13202
rect 209468 13012 209524 13022
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 185612 1204 185668 1214
rect 185612 644 185668 1148
rect 185612 578 185668 588
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 -1120 194078 9922
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 4350 221078 19842
rect 222460 17780 222516 17790
rect 222460 16884 222516 17724
rect 222460 16818 222516 16828
rect 222908 17668 222964 17678
rect 222908 16884 222964 17612
rect 222908 16818 222964 16828
rect 223132 17444 223188 17454
rect 223132 16660 223188 17388
rect 223356 17332 223412 17342
rect 223356 16884 223412 17276
rect 223356 16818 223412 16828
rect 223132 16594 223188 16604
rect 221340 14980 221396 14990
rect 221340 13978 221396 14924
rect 221340 13912 221396 13922
rect 222236 14980 222292 14990
rect 222236 13798 222292 14924
rect 222236 13732 222292 13742
rect 222012 12964 222068 12974
rect 222012 9658 222068 12908
rect 222012 9592 222068 9602
rect 223356 12292 223412 12302
rect 223356 6418 223412 12236
rect 223356 6352 223412 6362
rect 224178 10350 224798 19842
rect 228844 17556 228900 17566
rect 228844 16884 228900 17500
rect 226268 16858 226324 16868
rect 228844 16818 228900 16828
rect 230748 17218 230804 17228
rect 226268 16772 226324 16802
rect 226268 16706 226324 16716
rect 230748 16772 230804 17162
rect 230748 16706 230804 16716
rect 231196 16772 231252 19862
rect 239260 19558 239316 19568
rect 231196 16706 231252 16716
rect 236572 19378 236628 19388
rect 236572 16772 236628 19322
rect 236572 16706 236628 16716
rect 236796 17038 236852 17048
rect 226044 16100 226100 16110
rect 226044 15958 226100 16044
rect 226044 15892 226100 15902
rect 236124 13412 236180 13422
rect 231420 12740 231476 12750
rect 225036 12404 225092 12414
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 -1120 224798 9922
rect 224924 12292 224980 12302
rect 224924 6058 224980 12236
rect 225036 6238 225092 12348
rect 226604 12404 226660 12414
rect 226604 8398 226660 12348
rect 226604 8332 226660 8342
rect 226716 12292 226772 12302
rect 225036 6172 225092 6182
rect 224924 5992 224980 6002
rect 226716 5878 226772 12236
rect 228396 12292 228452 12302
rect 228396 7678 228452 12236
rect 228396 7612 228452 7622
rect 230076 12292 230132 12302
rect 230076 7498 230132 12236
rect 231420 9298 231476 12684
rect 231420 9232 231476 9242
rect 231644 12292 231700 12302
rect 231644 8428 231700 12236
rect 236124 11638 236180 13356
rect 236124 11572 236180 11582
rect 236796 10836 236852 16982
rect 239260 16772 239316 19502
rect 239260 16706 239316 16716
rect 240380 16772 240436 20942
rect 240380 16706 240436 16716
rect 240604 16772 240660 21122
rect 241948 19918 242004 21302
rect 241948 19852 242004 19862
rect 243740 19918 243796 19928
rect 241948 19738 242004 19748
rect 241724 17892 241780 17902
rect 241724 16884 241780 17836
rect 241724 16818 241780 16828
rect 240604 16706 240660 16716
rect 241948 16660 242004 19682
rect 243740 16772 243796 19862
rect 243740 16706 243796 16716
rect 245084 17578 245140 17588
rect 245084 16772 245140 17522
rect 245084 16706 245140 16716
rect 241948 16594 242004 16604
rect 245308 16324 245364 16334
rect 245308 16230 245364 16262
rect 238588 15238 238644 15248
rect 238476 12404 238532 12414
rect 238364 12292 238420 12302
rect 238364 12178 238420 12236
rect 236796 10770 236852 10780
rect 238252 12122 238420 12178
rect 231644 8372 231812 8428
rect 230076 7432 230132 7442
rect 231756 6598 231812 8372
rect 238252 8038 238308 12122
rect 238252 7972 238308 7982
rect 238364 11844 238420 11854
rect 231756 6532 231812 6542
rect 226716 5812 226772 5822
rect 238364 2818 238420 11788
rect 238364 2752 238420 2762
rect 238476 838 238532 12348
rect 238588 12180 238644 15182
rect 243068 14980 243124 14990
rect 243068 14338 243124 14924
rect 243068 14272 243124 14282
rect 241500 13412 241556 13422
rect 239148 13188 239204 13198
rect 239148 12404 239204 13132
rect 239148 12338 239204 12348
rect 241052 12852 241108 12862
rect 240156 12292 240212 12302
rect 240156 12178 240212 12236
rect 238588 12114 238644 12124
rect 240044 12122 240212 12178
rect 240044 2458 240100 12122
rect 240044 2392 240100 2402
rect 240156 11844 240212 11854
rect 238476 772 238532 782
rect 240156 658 240212 11788
rect 241052 7858 241108 12796
rect 241500 11458 241556 13356
rect 243516 13412 243572 13422
rect 242396 12852 242452 12862
rect 241500 11392 241556 11402
rect 241724 12292 241780 12302
rect 241052 7792 241108 7802
rect 241724 3178 241780 12236
rect 242396 9478 242452 12796
rect 242396 9412 242452 9422
rect 243292 12404 243348 12414
rect 241724 3112 241780 3122
rect 240156 592 240212 602
rect 243292 298 243348 12348
rect 243292 232 243348 242
rect 243404 11844 243460 11854
rect 243404 118 243460 11788
rect 243516 11818 243572 13356
rect 245980 13412 246036 13422
rect 245980 12898 246036 13356
rect 245980 12832 246036 12842
rect 249452 12740 249508 12750
rect 245196 12404 245252 12414
rect 243516 11752 243572 11762
rect 245084 12180 245140 12190
rect 245084 4798 245140 12124
rect 245084 4732 245140 4742
rect 245196 3358 245252 12348
rect 246876 12180 246932 12190
rect 246876 4978 246932 12124
rect 249452 12180 249508 12684
rect 249452 12114 249508 12124
rect 246876 4912 246932 4922
rect 245196 3292 245252 3302
rect 251178 4350 251798 19842
rect 252812 18004 252868 18014
rect 252028 17780 252084 17790
rect 252028 14644 252084 17724
rect 252028 14578 252084 14588
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 243404 52 243460 62
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 -160 251798 3922
rect 252812 1764 252868 17948
rect 252812 1698 252868 1708
rect 254898 10350 255518 19842
rect 256956 18452 257012 18462
rect 256844 17668 256900 17678
rect 256844 15092 256900 17612
rect 256956 17218 257012 18396
rect 256956 17152 257012 17162
rect 256844 15026 256900 15036
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 -1120 255518 9922
rect 264572 8260 264628 54602
rect 265244 31948 265300 87724
rect 265916 72660 265972 72670
rect 265916 69412 265972 72604
rect 265916 69346 265972 69356
rect 265916 66052 265972 66062
rect 265916 64036 265972 65996
rect 265916 63970 265972 63980
rect 265916 37156 265972 37166
rect 265916 35140 265972 37100
rect 265916 35074 265972 35084
rect 265020 31892 265300 31948
rect 266140 34468 266196 34478
rect 265020 26908 265076 31892
rect 265916 31780 265972 31790
rect 265916 28420 265972 31724
rect 266140 31556 266196 34412
rect 266140 31490 266196 31500
rect 265916 28354 265972 28364
rect 264796 26852 265076 26908
rect 264572 8194 264628 8204
rect 264684 20098 264740 20108
rect 264684 3332 264740 20042
rect 264796 11788 264852 26852
rect 265916 26404 265972 26414
rect 265468 23158 265524 23166
rect 265244 23156 265524 23158
rect 265244 23102 265468 23156
rect 265244 21898 265300 23102
rect 265468 23090 265524 23100
rect 265916 22148 265972 26348
rect 265916 22082 265972 22092
rect 265020 21842 265300 21898
rect 265020 18004 265076 21842
rect 265020 17938 265076 17948
rect 265916 19684 265972 19694
rect 265468 17444 265524 17454
rect 265468 12538 265524 17388
rect 265916 14308 265972 19628
rect 265916 14242 265972 14252
rect 265468 12472 265524 12482
rect 264796 11732 265300 11788
rect 265244 6356 265300 11732
rect 265244 6290 265300 6300
rect 265468 10164 265524 10174
rect 264684 3266 264740 3276
rect 265468 2818 265524 10108
rect 266252 6692 266308 97580
rect 266364 85798 266420 85808
rect 266364 17578 266420 85742
rect 266364 17512 266420 17522
rect 266476 8148 266532 97692
rect 267932 83748 267988 104102
rect 270620 92820 270676 92830
rect 270620 90748 270676 92764
rect 270620 90692 271012 90748
rect 269612 89124 269668 89134
rect 268156 87598 268212 87608
rect 267932 83682 267988 83692
rect 268044 85258 268100 85268
rect 266588 82740 266644 82750
rect 266588 21358 266644 82684
rect 266588 21292 266644 21302
rect 266700 78484 266756 78494
rect 266700 19918 266756 78428
rect 267932 77338 267988 77348
rect 267820 76804 267876 76814
rect 266924 73018 266980 73028
rect 266700 19852 266756 19862
rect 266812 69778 266868 69788
rect 266812 12964 266868 69722
rect 266924 17892 266980 72962
rect 267036 25060 267092 25070
rect 267036 20580 267092 25004
rect 267036 20514 267092 20524
rect 266924 17826 266980 17836
rect 267820 15958 267876 76748
rect 267820 15892 267876 15902
rect 267932 13438 267988 77282
rect 267932 13372 267988 13382
rect 266812 12898 266868 12908
rect 266476 8082 266532 8092
rect 267148 9716 267204 9726
rect 266252 6626 266308 6636
rect 265468 2752 265524 2762
rect 267148 2638 267204 9660
rect 268044 5124 268100 85202
rect 268156 16318 268212 87542
rect 268828 85978 268884 85988
rect 268380 85876 268436 85886
rect 268156 16252 268212 16262
rect 268268 84178 268324 84188
rect 268156 14196 268212 14206
rect 268156 10052 268212 14140
rect 268268 13258 268324 84122
rect 268380 14338 268436 85820
rect 268828 85764 268884 85922
rect 268828 85698 268884 85708
rect 268940 82918 268996 82928
rect 268940 82404 268996 82862
rect 268940 82338 268996 82348
rect 268716 77698 268772 77708
rect 268604 74098 268660 74108
rect 268380 14272 268436 14282
rect 268492 73198 268548 73208
rect 268268 13192 268324 13202
rect 268156 9986 268212 9996
rect 268044 5058 268100 5068
rect 268492 5012 268548 73142
rect 268604 14196 268660 74042
rect 268604 14130 268660 14140
rect 268604 13978 268660 13988
rect 268604 13188 268660 13922
rect 268604 13122 268660 13132
rect 268716 13076 268772 77642
rect 268828 75460 268884 75470
rect 268828 72100 268884 75404
rect 268828 72034 268884 72044
rect 268940 73892 268996 73902
rect 268940 70756 268996 73836
rect 268940 70690 268996 70700
rect 268828 69188 268884 69198
rect 268828 66724 268884 69132
rect 268828 66658 268884 66668
rect 268828 39844 268884 39854
rect 268828 37828 268884 39788
rect 268828 37762 268884 37772
rect 268828 33124 268884 33134
rect 268828 29988 268884 33068
rect 268828 29922 268884 29932
rect 268940 30436 268996 30446
rect 268828 29092 268884 29102
rect 268828 25284 268884 29036
rect 268940 26852 268996 30380
rect 268940 26786 268996 26796
rect 268828 25218 268884 25228
rect 268940 23716 268996 23726
rect 268828 22372 268884 22382
rect 268828 17444 268884 22316
rect 268940 19012 268996 23660
rect 268940 18946 268996 18956
rect 268828 17378 268884 17388
rect 268940 18340 268996 18350
rect 268716 13010 268772 13020
rect 268940 13078 268996 18284
rect 269052 17556 269108 17566
rect 269052 16318 269108 17500
rect 269052 16252 269108 16262
rect 269612 15148 269668 89068
rect 268940 13012 268996 13022
rect 269500 15092 269668 15148
rect 269724 88004 269780 88014
rect 269164 11060 269220 11070
rect 269164 8428 269220 11004
rect 269500 10164 269556 15092
rect 269724 14698 269780 87948
rect 270284 87668 270340 87678
rect 269948 86698 270004 86708
rect 269612 14642 269780 14698
rect 269836 77140 269892 77150
rect 269612 11458 269668 14642
rect 269612 11392 269668 11402
rect 269724 14420 269780 14430
rect 269500 10098 269556 10108
rect 269724 8596 269780 14364
rect 269724 8530 269780 8540
rect 269164 8372 269332 8428
rect 269276 8306 269332 8316
rect 268492 4946 268548 4956
rect 267148 2572 267204 2582
rect 269836 2100 269892 77084
rect 269948 12898 270004 86642
rect 270172 81844 270228 81854
rect 270060 70756 270116 70766
rect 270060 68516 270116 70700
rect 270060 68450 270116 68460
rect 270060 67620 270116 67630
rect 270060 65380 270116 67564
rect 270060 65314 270116 65324
rect 270060 38500 270116 38510
rect 270060 36260 270116 38444
rect 270060 36194 270116 36204
rect 270060 35588 270116 35598
rect 270060 33124 270116 35532
rect 270060 33058 270116 33068
rect 270060 27748 270116 27758
rect 270060 23716 270116 27692
rect 270060 23650 270116 23660
rect 270060 21028 270116 21038
rect 270060 15876 270116 20972
rect 270060 15810 270116 15820
rect 269948 12832 270004 12842
rect 270172 12292 270228 81788
rect 270284 21178 270340 87612
rect 270620 87556 270676 87566
rect 270508 79604 270564 79614
rect 270508 76804 270564 79548
rect 270620 77252 270676 87500
rect 270956 85708 271012 90692
rect 270956 85652 271236 85708
rect 270844 84084 270900 84094
rect 270620 77186 270676 77196
rect 270732 83098 270788 83108
rect 270732 76978 270788 83042
rect 270620 76922 270788 76978
rect 270620 76916 270676 76922
rect 270620 76850 270676 76860
rect 270508 76738 270564 76748
rect 270844 76618 270900 84028
rect 270284 21112 270340 21122
rect 270508 76562 270900 76618
rect 271068 83972 271124 83982
rect 270508 20998 270564 76562
rect 271068 76438 271124 83916
rect 270620 76382 271124 76438
rect 270620 76356 270676 76382
rect 270620 76290 270676 76300
rect 271180 73948 271236 85652
rect 270732 73892 271236 73948
rect 271292 80948 271348 80958
rect 270732 55468 270788 73892
rect 270508 20932 270564 20942
rect 270620 55412 270788 55468
rect 270508 15204 270564 15214
rect 270508 13978 270564 15148
rect 270284 13922 270564 13978
rect 270284 12898 270340 13922
rect 270620 13618 270676 55412
rect 271292 19558 271348 80892
rect 271516 78260 271572 108242
rect 272972 104158 273028 236796
rect 272972 104092 273028 104102
rect 273308 88564 273364 88574
rect 271516 78194 271572 78204
rect 272972 87892 273028 87902
rect 271632 76350 271952 76384
rect 271632 76294 271702 76350
rect 271758 76294 271826 76350
rect 271882 76294 271952 76350
rect 271632 76226 271952 76294
rect 271632 76170 271702 76226
rect 271758 76170 271826 76226
rect 271882 76170 271952 76226
rect 271632 76102 271952 76170
rect 271632 76046 271702 76102
rect 271758 76046 271826 76102
rect 271882 76046 271952 76102
rect 271632 75978 271952 76046
rect 271632 75922 271702 75978
rect 271758 75922 271826 75978
rect 271882 75922 271952 75978
rect 271632 75888 271952 75922
rect 271632 58350 271952 58384
rect 271632 58294 271702 58350
rect 271758 58294 271826 58350
rect 271882 58294 271952 58350
rect 271632 58226 271952 58294
rect 271632 58170 271702 58226
rect 271758 58170 271826 58226
rect 271882 58170 271952 58226
rect 271632 58102 271952 58170
rect 271632 58046 271702 58102
rect 271758 58046 271826 58102
rect 271882 58046 271952 58102
rect 271632 57978 271952 58046
rect 271632 57922 271702 57978
rect 271758 57922 271826 57978
rect 271882 57922 271952 57978
rect 271632 57888 271952 57922
rect 271632 40350 271952 40384
rect 271632 40294 271702 40350
rect 271758 40294 271826 40350
rect 271882 40294 271952 40350
rect 271632 40226 271952 40294
rect 271632 40170 271702 40226
rect 271758 40170 271826 40226
rect 271882 40170 271952 40226
rect 271632 40102 271952 40170
rect 271632 40046 271702 40102
rect 271758 40046 271826 40102
rect 271882 40046 271952 40102
rect 271632 39978 271952 40046
rect 271632 39922 271702 39978
rect 271758 39922 271826 39978
rect 271882 39922 271952 39978
rect 271632 39888 271952 39922
rect 271632 22350 271952 22384
rect 271632 22294 271702 22350
rect 271758 22294 271826 22350
rect 271882 22294 271952 22350
rect 271632 22226 271952 22294
rect 271632 22170 271702 22226
rect 271758 22170 271826 22226
rect 271882 22170 271952 22226
rect 271632 22102 271952 22170
rect 271632 22046 271702 22102
rect 271758 22046 271826 22102
rect 271882 22046 271952 22102
rect 271632 21978 271952 22046
rect 271632 21922 271702 21978
rect 271758 21922 271826 21978
rect 271882 21922 271952 21978
rect 271632 21888 271952 21922
rect 271292 19492 271348 19502
rect 272972 19378 273028 87836
rect 273084 85988 273140 85998
rect 273084 54658 273140 85932
rect 273084 54592 273140 54602
rect 273196 83748 273252 83758
rect 273196 19738 273252 83692
rect 273308 73198 273364 88508
rect 273532 86324 273588 86334
rect 273308 73132 273364 73142
rect 273420 78260 273476 78270
rect 273420 20098 273476 78204
rect 273532 73018 273588 86268
rect 273868 81478 273924 290612
rect 281898 274350 282518 291922
rect 281898 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 282518 274350
rect 281898 274226 282518 274294
rect 281898 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 282518 274226
rect 281898 274102 282518 274170
rect 281898 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 282518 274102
rect 281898 273978 282518 274046
rect 281898 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 282518 273978
rect 281898 256350 282518 273922
rect 281898 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 282518 256350
rect 281898 256226 282518 256294
rect 281898 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 282518 256226
rect 281898 256102 282518 256170
rect 281898 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 282518 256102
rect 281898 255978 282518 256046
rect 281898 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 282518 255978
rect 281898 238350 282518 255922
rect 281898 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 282518 238350
rect 281898 238226 282518 238294
rect 281898 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 282518 238226
rect 281898 238102 282518 238170
rect 281898 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 282518 238102
rect 281898 237978 282518 238046
rect 281898 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 282518 237978
rect 281898 220350 282518 237922
rect 281898 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 282518 220350
rect 281898 220226 282518 220294
rect 281898 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 282518 220226
rect 281898 220102 282518 220170
rect 281898 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 282518 220102
rect 281898 219978 282518 220046
rect 281898 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 282518 219978
rect 281898 202350 282518 219922
rect 281898 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 282518 202350
rect 281898 202226 282518 202294
rect 281898 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 282518 202226
rect 281898 202102 282518 202170
rect 281898 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 282518 202102
rect 281898 201978 282518 202046
rect 281898 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 282518 201978
rect 281898 184350 282518 201922
rect 281898 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 282518 184350
rect 281898 184226 282518 184294
rect 281898 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 282518 184226
rect 281898 184102 282518 184170
rect 281898 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 282518 184102
rect 281898 183978 282518 184046
rect 281898 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 282518 183978
rect 281898 166350 282518 183922
rect 281898 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 282518 166350
rect 281898 166226 282518 166294
rect 281898 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 282518 166226
rect 281898 166102 282518 166170
rect 281898 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 282518 166102
rect 281898 165978 282518 166046
rect 281898 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 282518 165978
rect 281898 148350 282518 165922
rect 281898 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 282518 148350
rect 281898 148226 282518 148294
rect 281898 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 282518 148226
rect 281898 148102 282518 148170
rect 281898 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 282518 148102
rect 281898 147978 282518 148046
rect 281898 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 282518 147978
rect 281898 130350 282518 147922
rect 281898 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 282518 130350
rect 281898 130226 282518 130294
rect 281898 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 282518 130226
rect 281898 130102 282518 130170
rect 281898 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 282518 130102
rect 281898 129978 282518 130046
rect 281898 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 282518 129978
rect 281898 112350 282518 129922
rect 281898 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 282518 112350
rect 281898 112226 282518 112294
rect 281898 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 282518 112226
rect 281898 112102 282518 112170
rect 281898 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 282518 112102
rect 281898 111978 282518 112046
rect 281898 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 282518 111978
rect 281898 94350 282518 111922
rect 281898 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 282518 94350
rect 281898 94226 282518 94294
rect 281898 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 282518 94226
rect 281898 94102 282518 94170
rect 273980 94052 274036 94062
rect 273980 92458 274036 93996
rect 273980 92392 274036 92402
rect 281898 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 282518 94102
rect 281898 93978 282518 94046
rect 281898 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 282518 93978
rect 273868 81412 273924 81422
rect 273532 72952 273588 72962
rect 273644 81172 273700 81182
rect 273644 69778 273700 81116
rect 274092 80500 274148 80510
rect 274092 74098 274148 80444
rect 281898 79630 282518 93922
rect 282604 305284 282660 305294
rect 282604 86518 282660 305228
rect 282604 86452 282660 86462
rect 285618 298350 286238 306466
rect 296492 305396 296548 305406
rect 285618 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 286238 298350
rect 285618 298226 286238 298294
rect 285618 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 286238 298226
rect 285618 298102 286238 298170
rect 285618 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 286238 298102
rect 285618 297978 286238 298046
rect 285618 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 286238 297978
rect 285618 280350 286238 297922
rect 285618 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 286238 280350
rect 285618 280226 286238 280294
rect 285618 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 286238 280226
rect 285618 280102 286238 280170
rect 285618 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 286238 280102
rect 285618 279978 286238 280046
rect 285618 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 286238 279978
rect 285618 262350 286238 279922
rect 285618 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 286238 262350
rect 285618 262226 286238 262294
rect 285618 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 286238 262226
rect 285618 262102 286238 262170
rect 285618 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 286238 262102
rect 285618 261978 286238 262046
rect 285618 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 286238 261978
rect 285618 244350 286238 261922
rect 285618 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 286238 244350
rect 285618 244226 286238 244294
rect 285618 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 286238 244226
rect 285618 244102 286238 244170
rect 285618 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 286238 244102
rect 285618 243978 286238 244046
rect 285618 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 286238 243978
rect 285618 226350 286238 243922
rect 285618 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 286238 226350
rect 285618 226226 286238 226294
rect 285618 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 286238 226226
rect 285618 226102 286238 226170
rect 285618 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 286238 226102
rect 285618 225978 286238 226046
rect 285618 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 286238 225978
rect 285618 208350 286238 225922
rect 285618 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 286238 208350
rect 285618 208226 286238 208294
rect 285618 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 286238 208226
rect 285618 208102 286238 208170
rect 285618 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 286238 208102
rect 285618 207978 286238 208046
rect 285618 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 286238 207978
rect 285618 190350 286238 207922
rect 285618 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 286238 190350
rect 285618 190226 286238 190294
rect 285618 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 286238 190226
rect 285618 190102 286238 190170
rect 285618 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 286238 190102
rect 285618 189978 286238 190046
rect 285618 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 286238 189978
rect 285618 172350 286238 189922
rect 285618 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 286238 172350
rect 285618 172226 286238 172294
rect 285618 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 286238 172226
rect 285618 172102 286238 172170
rect 285618 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 286238 172102
rect 285618 171978 286238 172046
rect 285618 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 286238 171978
rect 285618 154350 286238 171922
rect 285618 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 286238 154350
rect 285618 154226 286238 154294
rect 285618 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 286238 154226
rect 285618 154102 286238 154170
rect 285618 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 286238 154102
rect 285618 153978 286238 154046
rect 285618 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 286238 153978
rect 285618 136350 286238 153922
rect 285618 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 286238 136350
rect 285618 136226 286238 136294
rect 285618 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 286238 136226
rect 285618 136102 286238 136170
rect 285618 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 286238 136102
rect 285618 135978 286238 136046
rect 285618 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 286238 135978
rect 285618 118350 286238 135922
rect 285618 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 286238 118350
rect 285618 118226 286238 118294
rect 285618 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 286238 118226
rect 285618 118102 286238 118170
rect 285618 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 286238 118102
rect 285618 117978 286238 118046
rect 285618 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 286238 117978
rect 285618 100350 286238 117922
rect 286300 305284 286356 305294
rect 286300 108298 286356 305228
rect 286300 108232 286356 108242
rect 290668 305284 290724 305294
rect 285618 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 286238 100350
rect 285618 100226 286238 100294
rect 285618 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 286238 100226
rect 285618 100102 286238 100170
rect 285618 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 286238 100102
rect 285618 99978 286238 100046
rect 285618 99922 285714 99978
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 286238 99978
rect 283836 85764 283892 85774
rect 283836 85258 283892 85708
rect 283836 85192 283892 85202
rect 285618 82350 286238 99922
rect 290668 88318 290724 305228
rect 290668 88252 290724 88262
rect 292348 305284 292404 305294
rect 292348 88138 292404 305228
rect 294140 305284 294196 305294
rect 294140 290668 294196 305228
rect 294028 290612 294196 290668
rect 294028 88498 294084 290612
rect 294028 88432 294084 88442
rect 292348 88072 292404 88082
rect 296492 85078 296548 305340
rect 296492 85012 296548 85022
rect 299068 305284 299124 305294
rect 299068 84898 299124 305228
rect 310828 305284 310884 305294
rect 310828 305038 310884 305228
rect 310828 304972 310884 304982
rect 309148 304052 309204 304062
rect 309148 303238 309204 303996
rect 309148 303172 309204 303182
rect 310604 301258 310660 301268
rect 310828 301258 310884 301268
rect 310660 301202 310772 301258
rect 310604 301192 310660 301202
rect 310716 300898 310772 301202
rect 310828 301140 310884 301202
rect 310828 301074 310884 301084
rect 310716 300842 310884 300898
rect 310828 290668 310884 300842
rect 312618 292350 313238 306466
rect 315084 301618 315140 301628
rect 312618 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 313238 292350
rect 312618 292226 313238 292294
rect 312618 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 313238 292226
rect 312618 292102 313238 292170
rect 312618 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 313238 292102
rect 312618 291978 313238 292046
rect 312618 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 313238 291978
rect 310828 290612 311668 290668
rect 311612 93380 311668 290612
rect 311612 93314 311668 93324
rect 312618 274350 313238 291922
rect 312618 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 313238 274350
rect 312618 274226 313238 274294
rect 312618 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 313238 274226
rect 312618 274102 313238 274170
rect 312618 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 313238 274102
rect 312618 273978 313238 274046
rect 312618 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 313238 273978
rect 312618 256350 313238 273922
rect 312618 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 313238 256350
rect 312618 256226 313238 256294
rect 312618 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 313238 256226
rect 312618 256102 313238 256170
rect 312618 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 313238 256102
rect 312618 255978 313238 256046
rect 312618 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 313238 255978
rect 312618 238350 313238 255922
rect 312618 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 313238 238350
rect 312618 238226 313238 238294
rect 312618 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 313238 238226
rect 312618 238102 313238 238170
rect 312618 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 313238 238102
rect 312618 237978 313238 238046
rect 312618 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 313238 237978
rect 312618 220350 313238 237922
rect 312618 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 313238 220350
rect 312618 220226 313238 220294
rect 312618 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 313238 220226
rect 312618 220102 313238 220170
rect 312618 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 313238 220102
rect 312618 219978 313238 220046
rect 312618 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 313238 219978
rect 312618 202350 313238 219922
rect 312618 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 313238 202350
rect 312618 202226 313238 202294
rect 312618 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 313238 202226
rect 312618 202102 313238 202170
rect 312618 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 313238 202102
rect 312618 201978 313238 202046
rect 312618 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 313238 201978
rect 312618 184350 313238 201922
rect 312618 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 313238 184350
rect 312618 184226 313238 184294
rect 312618 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 313238 184226
rect 312618 184102 313238 184170
rect 312618 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 313238 184102
rect 312618 183978 313238 184046
rect 312618 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 313238 183978
rect 312618 166350 313238 183922
rect 312618 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 313238 166350
rect 312618 166226 313238 166294
rect 312618 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 313238 166226
rect 312618 166102 313238 166170
rect 312618 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 313238 166102
rect 312618 165978 313238 166046
rect 312618 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 313238 165978
rect 312618 148350 313238 165922
rect 312618 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 313238 148350
rect 312618 148226 313238 148294
rect 312618 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 313238 148226
rect 312618 148102 313238 148170
rect 312618 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 313238 148102
rect 312618 147978 313238 148046
rect 312618 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 313238 147978
rect 312618 130350 313238 147922
rect 312618 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 313238 130350
rect 312618 130226 313238 130294
rect 312618 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 313238 130226
rect 312618 130102 313238 130170
rect 312618 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 313238 130102
rect 312618 129978 313238 130046
rect 312618 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 313238 129978
rect 312618 112350 313238 129922
rect 312618 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 313238 112350
rect 312618 112226 313238 112294
rect 312618 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 313238 112226
rect 312618 112102 313238 112170
rect 312618 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 313238 112102
rect 312618 111978 313238 112046
rect 312618 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 313238 111978
rect 312618 94350 313238 111922
rect 312618 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 313238 94350
rect 312618 94226 313238 94294
rect 312618 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 313238 94226
rect 312618 94102 313238 94170
rect 312618 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 313238 94102
rect 312618 93978 313238 94046
rect 312618 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 313238 93978
rect 299068 84832 299124 84842
rect 285618 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 286238 82350
rect 285618 82226 286238 82294
rect 285618 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 286238 82226
rect 285618 82102 286238 82170
rect 285618 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 286238 82102
rect 285618 81978 286238 82046
rect 285618 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 286238 81978
rect 285618 79630 286238 81922
rect 312618 79630 313238 93922
rect 314972 296548 315028 296558
rect 314972 78958 315028 296492
rect 315084 90132 315140 301562
rect 315084 90066 315140 90076
rect 316338 298350 316958 306466
rect 320684 305732 320740 305742
rect 320012 305508 320068 305518
rect 320012 304500 320068 305452
rect 320012 304434 320068 304444
rect 319004 303380 319060 303390
rect 319004 302518 319060 303324
rect 319004 302452 319060 302462
rect 320684 302158 320740 305676
rect 324156 305732 324212 305742
rect 322588 305060 322644 305070
rect 320796 304724 320852 304734
rect 320796 302338 320852 304668
rect 322588 302596 322644 305004
rect 324156 304858 324212 305676
rect 324156 304792 324212 304802
rect 324604 305732 324660 305742
rect 324604 303418 324660 305676
rect 324604 303352 324660 303362
rect 327292 305732 327348 305742
rect 324492 303238 324548 303248
rect 324492 302820 324548 303182
rect 327292 303238 327348 305676
rect 330428 305732 330484 305742
rect 327740 305038 327796 305048
rect 327740 304164 327796 304982
rect 327740 304098 327796 304108
rect 329196 304388 329252 304398
rect 327292 303172 327348 303182
rect 329196 302932 329252 304332
rect 330428 304138 330484 305676
rect 336476 305732 336532 305742
rect 331548 305620 331604 305630
rect 330428 304072 330484 304082
rect 330876 305508 330932 305518
rect 330876 303778 330932 305452
rect 330876 303712 330932 303722
rect 330988 304836 331044 304846
rect 330988 303716 331044 304780
rect 330988 303650 331044 303660
rect 329196 302866 329252 302876
rect 324492 302754 324548 302764
rect 322588 302530 322644 302540
rect 320796 302272 320852 302282
rect 329868 302338 329924 302348
rect 320684 302092 320740 302102
rect 329420 302158 329476 302168
rect 321692 301476 321748 301486
rect 316338 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 316958 298350
rect 316338 298226 316958 298294
rect 316338 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 316958 298226
rect 316338 298102 316958 298170
rect 316338 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 316958 298102
rect 316338 297978 316958 298046
rect 316338 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 316958 297978
rect 316338 280350 316958 297922
rect 316338 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 316958 280350
rect 316338 280226 316958 280294
rect 316338 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 316958 280226
rect 316338 280102 316958 280170
rect 316338 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 316958 280102
rect 316338 279978 316958 280046
rect 316338 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 316958 279978
rect 316338 262350 316958 279922
rect 316338 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 316958 262350
rect 316338 262226 316958 262294
rect 316338 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 316958 262226
rect 316338 262102 316958 262170
rect 316338 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 316958 262102
rect 316338 261978 316958 262046
rect 316338 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 316958 261978
rect 316338 244350 316958 261922
rect 316338 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 316958 244350
rect 316338 244226 316958 244294
rect 316338 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 316958 244226
rect 316338 244102 316958 244170
rect 316338 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 316958 244102
rect 316338 243978 316958 244046
rect 316338 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 316958 243978
rect 316338 226350 316958 243922
rect 316338 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 316958 226350
rect 316338 226226 316958 226294
rect 316338 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 316958 226226
rect 316338 226102 316958 226170
rect 316338 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 316958 226102
rect 316338 225978 316958 226046
rect 316338 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 316958 225978
rect 316338 208350 316958 225922
rect 316338 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 316958 208350
rect 316338 208226 316958 208294
rect 316338 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 316958 208226
rect 316338 208102 316958 208170
rect 316338 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 316958 208102
rect 316338 207978 316958 208046
rect 316338 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 316958 207978
rect 316338 190350 316958 207922
rect 316338 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 316958 190350
rect 316338 190226 316958 190294
rect 316338 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 316958 190226
rect 316338 190102 316958 190170
rect 316338 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 316958 190102
rect 316338 189978 316958 190046
rect 316338 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 316958 189978
rect 316338 172350 316958 189922
rect 316338 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 316958 172350
rect 316338 172226 316958 172294
rect 316338 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 316958 172226
rect 316338 172102 316958 172170
rect 316338 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 316958 172102
rect 316338 171978 316958 172046
rect 316338 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 316958 171978
rect 316338 154350 316958 171922
rect 316338 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 316958 154350
rect 316338 154226 316958 154294
rect 316338 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 316958 154226
rect 316338 154102 316958 154170
rect 316338 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 316958 154102
rect 316338 153978 316958 154046
rect 316338 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 316958 153978
rect 316338 136350 316958 153922
rect 316338 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 316958 136350
rect 316338 136226 316958 136294
rect 316338 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 316958 136226
rect 316338 136102 316958 136170
rect 316338 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 316958 136102
rect 316338 135978 316958 136046
rect 316338 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 316958 135978
rect 316338 118350 316958 135922
rect 316338 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 316958 118350
rect 316338 118226 316958 118294
rect 316338 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 316958 118226
rect 316338 118102 316958 118170
rect 316338 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 316958 118102
rect 316338 117978 316958 118046
rect 316338 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 316958 117978
rect 316338 100350 316958 117922
rect 316338 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 316958 100350
rect 316338 100226 316958 100294
rect 316338 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 316958 100226
rect 316338 100102 316958 100170
rect 316338 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 316958 100102
rect 316338 99978 316958 100046
rect 316338 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 316958 99978
rect 316338 82350 316958 99922
rect 318332 301438 318388 301448
rect 318332 90244 318388 301382
rect 318332 90178 318388 90188
rect 317436 88004 317492 88014
rect 317436 86698 317492 87948
rect 317436 86632 317492 86642
rect 317436 84358 317492 84368
rect 317436 83098 317492 84302
rect 321692 83412 321748 301420
rect 329420 300804 329476 302102
rect 329420 300738 329476 300748
rect 329868 300804 329924 302282
rect 329868 300738 329924 300748
rect 331548 300804 331604 305564
rect 334236 305172 334292 305182
rect 332556 302518 332612 302528
rect 332556 300916 332612 302462
rect 334236 301364 334292 305116
rect 336476 305038 336532 305676
rect 336476 304972 336532 304982
rect 342524 305732 342580 305742
rect 341404 304612 341460 304622
rect 336028 303940 336084 303950
rect 336028 303598 336084 303884
rect 336028 303532 336084 303542
rect 334236 301298 334292 301308
rect 341404 301140 341460 304556
rect 342524 304318 342580 305676
rect 342524 304252 342580 304262
rect 342972 305732 343028 305742
rect 342972 303958 343028 305676
rect 344652 304858 344708 304868
rect 344652 304164 344708 304802
rect 344652 304098 344708 304108
rect 342972 303892 343028 303902
rect 341404 301074 341460 301084
rect 342636 303418 342692 303428
rect 332556 300850 332612 300860
rect 331548 300738 331604 300748
rect 342636 300804 342692 303362
rect 344428 303238 344484 303248
rect 344316 302036 344372 302046
rect 344316 301618 344372 301980
rect 344316 301552 344372 301562
rect 344428 301028 344484 303182
rect 344428 300962 344484 300972
rect 342636 300738 342692 300748
rect 347058 298350 347678 306466
rect 352380 305732 352436 305742
rect 349580 305508 349636 305518
rect 347788 303778 347844 303788
rect 347788 302596 347844 303722
rect 347788 302530 347844 302540
rect 349580 300916 349636 305452
rect 351372 304138 351428 304148
rect 351036 303598 351092 303608
rect 351036 302932 351092 303542
rect 351036 302866 351092 302876
rect 349580 300850 349636 300860
rect 351372 300804 351428 304082
rect 352380 304138 352436 305676
rect 357756 305732 357812 305742
rect 352828 305396 352884 305406
rect 352828 304836 352884 305340
rect 352828 304770 352884 304780
rect 355852 305038 355908 305048
rect 352380 304072 352436 304082
rect 354396 304500 354452 304510
rect 354396 302596 354452 304444
rect 355852 304164 355908 304982
rect 357756 304858 357812 305676
rect 357756 304792 357812 304802
rect 360892 305732 360948 305742
rect 355852 304098 355908 304108
rect 357756 304318 357812 304328
rect 354396 302530 354452 302540
rect 357756 301364 357812 304262
rect 360892 303598 360948 305676
rect 369404 305732 369460 305742
rect 362684 305620 362740 305630
rect 361900 305060 361956 305070
rect 361900 304388 361956 305004
rect 361900 304322 361956 304332
rect 360892 303532 360948 303542
rect 362684 303238 362740 305564
rect 364588 304948 364644 304958
rect 362684 303172 362740 303182
rect 363468 303958 363524 303968
rect 363468 302484 363524 303902
rect 363468 302418 363524 302428
rect 364588 302338 364644 304892
rect 366268 304612 366324 304622
rect 366268 304052 366324 304556
rect 366268 303986 366324 303996
rect 369404 303958 369460 305676
rect 369404 303892 369460 303902
rect 371084 305284 371140 305294
rect 369516 302932 369572 302942
rect 364588 302272 364644 302282
rect 367612 302372 367668 302382
rect 357756 301298 357812 301308
rect 364812 301618 364868 301628
rect 351372 300738 351428 300748
rect 364812 300804 364868 301562
rect 367612 301618 367668 302316
rect 367612 301552 367668 301562
rect 369516 301364 369572 302876
rect 371084 301476 371140 305228
rect 376460 304858 376516 304868
rect 372988 304612 373044 304622
rect 371084 301410 371140 301420
rect 372428 304138 372484 304148
rect 369516 301298 369572 301308
rect 364812 300738 364868 300748
rect 372428 300804 372484 304082
rect 372428 300738 372484 300748
rect 372988 300804 373044 304556
rect 376460 304164 376516 304802
rect 376460 304098 376516 304108
rect 377580 304052 377636 304062
rect 377580 302372 377636 303996
rect 374556 302338 374612 302348
rect 377580 302306 377636 302316
rect 374332 302148 374388 302158
rect 374332 301798 374388 302092
rect 374332 301732 374388 301742
rect 374556 300916 374612 302282
rect 374556 300850 374612 300860
rect 372988 300738 373044 300748
rect 377778 298350 378398 306466
rect 379596 305732 379652 305742
rect 378812 305508 378868 305518
rect 378812 305172 378868 305452
rect 378812 305106 378868 305116
rect 379596 303778 379652 305676
rect 381052 305732 381108 305742
rect 381052 304858 381108 305676
rect 381052 304792 381108 304802
rect 394492 305284 394548 305294
rect 379596 303712 379652 303722
rect 383068 304724 383124 304734
rect 381388 303598 381444 303608
rect 379708 303238 379764 303248
rect 379708 300804 379764 303182
rect 381388 303156 381444 303542
rect 381388 303090 381444 303100
rect 383068 302484 383124 304668
rect 388444 304724 388500 304734
rect 388444 304164 388500 304668
rect 388444 304098 388500 304108
rect 389900 303958 389956 303968
rect 389900 303156 389956 303902
rect 394492 303238 394548 305228
rect 401548 304858 401604 304868
rect 394492 303172 394548 303182
rect 398076 304276 398132 304286
rect 389900 303090 389956 303100
rect 398076 302932 398132 304220
rect 401548 304164 401604 304802
rect 401548 304098 401604 304108
rect 405244 304164 405300 304174
rect 398412 303778 398468 303788
rect 398412 303156 398468 303722
rect 398412 303090 398468 303100
rect 398076 302866 398132 302876
rect 383068 302418 383124 302428
rect 393148 302260 393204 302270
rect 393148 302158 393204 302204
rect 393148 302092 393204 302102
rect 399756 302158 399812 302168
rect 394828 301798 394884 301808
rect 379708 300738 379764 300748
rect 388108 301618 388164 301628
rect 388108 300804 388164 301562
rect 388108 300738 388164 300748
rect 394828 300804 394884 301742
rect 394828 300738 394884 300748
rect 399756 300804 399812 302102
rect 399756 300738 399812 300748
rect 332332 298340 332388 298350
rect 332332 298004 332388 298284
rect 347058 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 347678 298350
rect 332332 297938 332388 297948
rect 337708 298228 337764 298238
rect 337708 297892 337764 298172
rect 337708 297826 337764 297836
rect 343532 298228 343588 298238
rect 343532 297892 343588 298172
rect 343532 297826 343588 297836
rect 347058 298226 347678 298294
rect 347058 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 347678 298226
rect 347058 298102 347678 298170
rect 347058 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 347678 298102
rect 347058 297978 347678 298046
rect 347058 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 347678 297978
rect 352716 298340 352772 298350
rect 352716 298004 352772 298284
rect 377778 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 378398 298350
rect 352716 297938 352772 297948
rect 356188 298228 356244 298238
rect 347058 297430 347678 297922
rect 356188 297892 356244 298172
rect 356188 297826 356244 297836
rect 371084 298228 371140 298238
rect 371084 297892 371140 298172
rect 371084 297826 371140 297836
rect 377778 298226 378398 298294
rect 384972 298340 385028 298350
rect 377778 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 378398 298226
rect 377778 298102 378398 298170
rect 377778 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 378398 298102
rect 377778 297978 378398 298046
rect 377778 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 378398 297978
rect 377778 297430 378398 297922
rect 384860 298228 384916 298238
rect 384860 297892 384916 298172
rect 384972 298004 385028 298284
rect 384972 297938 385028 297948
rect 384860 297826 384916 297836
rect 405244 296772 405300 304108
rect 408498 298350 409118 306466
rect 414092 302428 414148 337708
rect 408498 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 409118 298350
rect 408498 298226 409118 298294
rect 408498 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 409118 298226
rect 408498 298102 409118 298170
rect 408498 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 409118 298102
rect 408498 297978 409118 298046
rect 408498 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 409118 297978
rect 408498 297430 409118 297922
rect 413980 302372 414148 302428
rect 414988 303238 415044 303248
rect 405244 296706 405300 296716
rect 413980 296660 414036 302372
rect 414988 300804 415044 303182
rect 415772 301588 415828 353948
rect 415996 339892 416052 339902
rect 415996 301700 416052 339836
rect 416108 304388 416164 364700
rect 417452 359380 417508 359390
rect 416668 347956 416724 347966
rect 416668 346948 416724 347900
rect 416668 346882 416724 346892
rect 416780 347284 416836 347294
rect 416780 343588 416836 347228
rect 416780 343522 416836 343532
rect 416668 341908 416724 341918
rect 416668 340228 416724 341852
rect 416668 340162 416724 340172
rect 416668 323764 416724 323774
rect 416668 320068 416724 323708
rect 416668 320002 416724 320012
rect 416108 304322 416164 304332
rect 417452 301924 417508 359324
rect 417564 350980 417620 373436
rect 417676 372148 417732 372158
rect 417676 353668 417732 372092
rect 417900 371476 417956 371486
rect 417676 353602 417732 353612
rect 417788 356692 417844 356702
rect 417564 350914 417620 350924
rect 417564 348628 417620 348638
rect 417564 313348 417620 348572
rect 417564 313282 417620 313292
rect 417676 345940 417732 345950
rect 417452 301858 417508 301868
rect 417676 301812 417732 345884
rect 417788 323428 417844 356636
rect 417900 348740 417956 371420
rect 418348 368788 418404 368798
rect 418348 365540 418404 368732
rect 418348 365474 418404 365484
rect 419020 366100 419076 366110
rect 417900 348674 417956 348684
rect 418012 353332 418068 353342
rect 418012 345380 418068 353276
rect 418236 350644 418292 350654
rect 418236 348628 418292 350588
rect 418236 348562 418292 348572
rect 418012 345314 418068 345324
rect 418236 345268 418292 345278
rect 418236 323540 418292 345212
rect 418236 323474 418292 323484
rect 417788 323362 417844 323372
rect 418012 323092 418068 323102
rect 417676 301746 417732 301756
rect 417788 321076 417844 321086
rect 415996 301634 416052 301644
rect 415772 301522 415828 301532
rect 414988 300738 415044 300748
rect 414092 298788 414148 298798
rect 414092 298116 414148 298732
rect 414092 298050 414148 298060
rect 413980 296594 414036 296604
rect 417788 296660 417844 321020
rect 418012 298788 418068 323036
rect 419020 311556 419076 366044
rect 419916 365428 419972 365438
rect 419804 360724 419860 360734
rect 419692 358036 419748 358046
rect 419468 333844 419524 333854
rect 419356 328468 419412 328478
rect 419244 325108 419300 325118
rect 419020 311490 419076 311500
rect 419132 321748 419188 321758
rect 418012 298722 418068 298732
rect 417788 296594 417844 296604
rect 324448 292350 324768 292384
rect 324448 292294 324518 292350
rect 324574 292294 324642 292350
rect 324698 292294 324768 292350
rect 324448 292226 324768 292294
rect 324448 292170 324518 292226
rect 324574 292170 324642 292226
rect 324698 292170 324768 292226
rect 324448 292102 324768 292170
rect 324448 292046 324518 292102
rect 324574 292046 324642 292102
rect 324698 292046 324768 292102
rect 324448 291978 324768 292046
rect 324448 291922 324518 291978
rect 324574 291922 324642 291978
rect 324698 291922 324768 291978
rect 324448 291888 324768 291922
rect 355168 292350 355488 292384
rect 355168 292294 355238 292350
rect 355294 292294 355362 292350
rect 355418 292294 355488 292350
rect 355168 292226 355488 292294
rect 355168 292170 355238 292226
rect 355294 292170 355362 292226
rect 355418 292170 355488 292226
rect 355168 292102 355488 292170
rect 355168 292046 355238 292102
rect 355294 292046 355362 292102
rect 355418 292046 355488 292102
rect 355168 291978 355488 292046
rect 355168 291922 355238 291978
rect 355294 291922 355362 291978
rect 355418 291922 355488 291978
rect 355168 291888 355488 291922
rect 385888 292350 386208 292384
rect 385888 292294 385958 292350
rect 386014 292294 386082 292350
rect 386138 292294 386208 292350
rect 385888 292226 386208 292294
rect 385888 292170 385958 292226
rect 386014 292170 386082 292226
rect 386138 292170 386208 292226
rect 385888 292102 386208 292170
rect 385888 292046 385958 292102
rect 386014 292046 386082 292102
rect 386138 292046 386208 292102
rect 385888 291978 386208 292046
rect 385888 291922 385958 291978
rect 386014 291922 386082 291978
rect 386138 291922 386208 291978
rect 385888 291888 386208 291922
rect 416608 292350 416928 292384
rect 416608 292294 416678 292350
rect 416734 292294 416802 292350
rect 416858 292294 416928 292350
rect 416608 292226 416928 292294
rect 416608 292170 416678 292226
rect 416734 292170 416802 292226
rect 416858 292170 416928 292226
rect 416608 292102 416928 292170
rect 416608 292046 416678 292102
rect 416734 292046 416802 292102
rect 416858 292046 416928 292102
rect 416608 291978 416928 292046
rect 416608 291922 416678 291978
rect 416734 291922 416802 291978
rect 416858 291922 416928 291978
rect 416608 291888 416928 291922
rect 339808 280350 340128 280384
rect 339808 280294 339878 280350
rect 339934 280294 340002 280350
rect 340058 280294 340128 280350
rect 339808 280226 340128 280294
rect 339808 280170 339878 280226
rect 339934 280170 340002 280226
rect 340058 280170 340128 280226
rect 339808 280102 340128 280170
rect 339808 280046 339878 280102
rect 339934 280046 340002 280102
rect 340058 280046 340128 280102
rect 339808 279978 340128 280046
rect 339808 279922 339878 279978
rect 339934 279922 340002 279978
rect 340058 279922 340128 279978
rect 339808 279888 340128 279922
rect 370528 280350 370848 280384
rect 370528 280294 370598 280350
rect 370654 280294 370722 280350
rect 370778 280294 370848 280350
rect 370528 280226 370848 280294
rect 370528 280170 370598 280226
rect 370654 280170 370722 280226
rect 370778 280170 370848 280226
rect 370528 280102 370848 280170
rect 370528 280046 370598 280102
rect 370654 280046 370722 280102
rect 370778 280046 370848 280102
rect 370528 279978 370848 280046
rect 370528 279922 370598 279978
rect 370654 279922 370722 279978
rect 370778 279922 370848 279978
rect 370528 279888 370848 279922
rect 401248 280350 401568 280384
rect 401248 280294 401318 280350
rect 401374 280294 401442 280350
rect 401498 280294 401568 280350
rect 401248 280226 401568 280294
rect 401248 280170 401318 280226
rect 401374 280170 401442 280226
rect 401498 280170 401568 280226
rect 401248 280102 401568 280170
rect 401248 280046 401318 280102
rect 401374 280046 401442 280102
rect 401498 280046 401568 280102
rect 401248 279978 401568 280046
rect 401248 279922 401318 279978
rect 401374 279922 401442 279978
rect 401498 279922 401568 279978
rect 401248 279888 401568 279922
rect 324448 274350 324768 274384
rect 324448 274294 324518 274350
rect 324574 274294 324642 274350
rect 324698 274294 324768 274350
rect 324448 274226 324768 274294
rect 324448 274170 324518 274226
rect 324574 274170 324642 274226
rect 324698 274170 324768 274226
rect 324448 274102 324768 274170
rect 324448 274046 324518 274102
rect 324574 274046 324642 274102
rect 324698 274046 324768 274102
rect 324448 273978 324768 274046
rect 324448 273922 324518 273978
rect 324574 273922 324642 273978
rect 324698 273922 324768 273978
rect 324448 273888 324768 273922
rect 355168 274350 355488 274384
rect 355168 274294 355238 274350
rect 355294 274294 355362 274350
rect 355418 274294 355488 274350
rect 355168 274226 355488 274294
rect 355168 274170 355238 274226
rect 355294 274170 355362 274226
rect 355418 274170 355488 274226
rect 355168 274102 355488 274170
rect 355168 274046 355238 274102
rect 355294 274046 355362 274102
rect 355418 274046 355488 274102
rect 355168 273978 355488 274046
rect 355168 273922 355238 273978
rect 355294 273922 355362 273978
rect 355418 273922 355488 273978
rect 355168 273888 355488 273922
rect 385888 274350 386208 274384
rect 385888 274294 385958 274350
rect 386014 274294 386082 274350
rect 386138 274294 386208 274350
rect 385888 274226 386208 274294
rect 385888 274170 385958 274226
rect 386014 274170 386082 274226
rect 386138 274170 386208 274226
rect 385888 274102 386208 274170
rect 385888 274046 385958 274102
rect 386014 274046 386082 274102
rect 386138 274046 386208 274102
rect 385888 273978 386208 274046
rect 385888 273922 385958 273978
rect 386014 273922 386082 273978
rect 386138 273922 386208 273978
rect 385888 273888 386208 273922
rect 416608 274350 416928 274384
rect 416608 274294 416678 274350
rect 416734 274294 416802 274350
rect 416858 274294 416928 274350
rect 416608 274226 416928 274294
rect 416608 274170 416678 274226
rect 416734 274170 416802 274226
rect 416858 274170 416928 274226
rect 416608 274102 416928 274170
rect 416608 274046 416678 274102
rect 416734 274046 416802 274102
rect 416858 274046 416928 274102
rect 416608 273978 416928 274046
rect 416608 273922 416678 273978
rect 416734 273922 416802 273978
rect 416858 273922 416928 273978
rect 416608 273888 416928 273922
rect 339808 262350 340128 262384
rect 339808 262294 339878 262350
rect 339934 262294 340002 262350
rect 340058 262294 340128 262350
rect 339808 262226 340128 262294
rect 339808 262170 339878 262226
rect 339934 262170 340002 262226
rect 340058 262170 340128 262226
rect 339808 262102 340128 262170
rect 339808 262046 339878 262102
rect 339934 262046 340002 262102
rect 340058 262046 340128 262102
rect 339808 261978 340128 262046
rect 339808 261922 339878 261978
rect 339934 261922 340002 261978
rect 340058 261922 340128 261978
rect 339808 261888 340128 261922
rect 370528 262350 370848 262384
rect 370528 262294 370598 262350
rect 370654 262294 370722 262350
rect 370778 262294 370848 262350
rect 370528 262226 370848 262294
rect 370528 262170 370598 262226
rect 370654 262170 370722 262226
rect 370778 262170 370848 262226
rect 370528 262102 370848 262170
rect 370528 262046 370598 262102
rect 370654 262046 370722 262102
rect 370778 262046 370848 262102
rect 370528 261978 370848 262046
rect 370528 261922 370598 261978
rect 370654 261922 370722 261978
rect 370778 261922 370848 261978
rect 370528 261888 370848 261922
rect 401248 262350 401568 262384
rect 401248 262294 401318 262350
rect 401374 262294 401442 262350
rect 401498 262294 401568 262350
rect 401248 262226 401568 262294
rect 401248 262170 401318 262226
rect 401374 262170 401442 262226
rect 401498 262170 401568 262226
rect 401248 262102 401568 262170
rect 401248 262046 401318 262102
rect 401374 262046 401442 262102
rect 401498 262046 401568 262102
rect 401248 261978 401568 262046
rect 401248 261922 401318 261978
rect 401374 261922 401442 261978
rect 401498 261922 401568 261978
rect 401248 261888 401568 261922
rect 324448 256350 324768 256384
rect 324448 256294 324518 256350
rect 324574 256294 324642 256350
rect 324698 256294 324768 256350
rect 324448 256226 324768 256294
rect 324448 256170 324518 256226
rect 324574 256170 324642 256226
rect 324698 256170 324768 256226
rect 324448 256102 324768 256170
rect 324448 256046 324518 256102
rect 324574 256046 324642 256102
rect 324698 256046 324768 256102
rect 324448 255978 324768 256046
rect 324448 255922 324518 255978
rect 324574 255922 324642 255978
rect 324698 255922 324768 255978
rect 324448 255888 324768 255922
rect 355168 256350 355488 256384
rect 355168 256294 355238 256350
rect 355294 256294 355362 256350
rect 355418 256294 355488 256350
rect 355168 256226 355488 256294
rect 355168 256170 355238 256226
rect 355294 256170 355362 256226
rect 355418 256170 355488 256226
rect 355168 256102 355488 256170
rect 355168 256046 355238 256102
rect 355294 256046 355362 256102
rect 355418 256046 355488 256102
rect 355168 255978 355488 256046
rect 355168 255922 355238 255978
rect 355294 255922 355362 255978
rect 355418 255922 355488 255978
rect 355168 255888 355488 255922
rect 385888 256350 386208 256384
rect 385888 256294 385958 256350
rect 386014 256294 386082 256350
rect 386138 256294 386208 256350
rect 385888 256226 386208 256294
rect 385888 256170 385958 256226
rect 386014 256170 386082 256226
rect 386138 256170 386208 256226
rect 385888 256102 386208 256170
rect 385888 256046 385958 256102
rect 386014 256046 386082 256102
rect 386138 256046 386208 256102
rect 385888 255978 386208 256046
rect 385888 255922 385958 255978
rect 386014 255922 386082 255978
rect 386138 255922 386208 255978
rect 385888 255888 386208 255922
rect 416608 256350 416928 256384
rect 416608 256294 416678 256350
rect 416734 256294 416802 256350
rect 416858 256294 416928 256350
rect 416608 256226 416928 256294
rect 416608 256170 416678 256226
rect 416734 256170 416802 256226
rect 416858 256170 416928 256226
rect 416608 256102 416928 256170
rect 416608 256046 416678 256102
rect 416734 256046 416802 256102
rect 416858 256046 416928 256102
rect 416608 255978 416928 256046
rect 416608 255922 416678 255978
rect 416734 255922 416802 255978
rect 416858 255922 416928 255978
rect 416608 255888 416928 255922
rect 339808 244350 340128 244384
rect 339808 244294 339878 244350
rect 339934 244294 340002 244350
rect 340058 244294 340128 244350
rect 339808 244226 340128 244294
rect 339808 244170 339878 244226
rect 339934 244170 340002 244226
rect 340058 244170 340128 244226
rect 339808 244102 340128 244170
rect 339808 244046 339878 244102
rect 339934 244046 340002 244102
rect 340058 244046 340128 244102
rect 339808 243978 340128 244046
rect 339808 243922 339878 243978
rect 339934 243922 340002 243978
rect 340058 243922 340128 243978
rect 339808 243888 340128 243922
rect 370528 244350 370848 244384
rect 370528 244294 370598 244350
rect 370654 244294 370722 244350
rect 370778 244294 370848 244350
rect 370528 244226 370848 244294
rect 370528 244170 370598 244226
rect 370654 244170 370722 244226
rect 370778 244170 370848 244226
rect 370528 244102 370848 244170
rect 370528 244046 370598 244102
rect 370654 244046 370722 244102
rect 370778 244046 370848 244102
rect 370528 243978 370848 244046
rect 370528 243922 370598 243978
rect 370654 243922 370722 243978
rect 370778 243922 370848 243978
rect 370528 243888 370848 243922
rect 401248 244350 401568 244384
rect 401248 244294 401318 244350
rect 401374 244294 401442 244350
rect 401498 244294 401568 244350
rect 401248 244226 401568 244294
rect 401248 244170 401318 244226
rect 401374 244170 401442 244226
rect 401498 244170 401568 244226
rect 401248 244102 401568 244170
rect 401248 244046 401318 244102
rect 401374 244046 401442 244102
rect 401498 244046 401568 244102
rect 401248 243978 401568 244046
rect 401248 243922 401318 243978
rect 401374 243922 401442 243978
rect 401498 243922 401568 243978
rect 401248 243888 401568 243922
rect 324448 238350 324768 238384
rect 324448 238294 324518 238350
rect 324574 238294 324642 238350
rect 324698 238294 324768 238350
rect 324448 238226 324768 238294
rect 324448 238170 324518 238226
rect 324574 238170 324642 238226
rect 324698 238170 324768 238226
rect 324448 238102 324768 238170
rect 324448 238046 324518 238102
rect 324574 238046 324642 238102
rect 324698 238046 324768 238102
rect 324448 237978 324768 238046
rect 324448 237922 324518 237978
rect 324574 237922 324642 237978
rect 324698 237922 324768 237978
rect 324448 237888 324768 237922
rect 355168 238350 355488 238384
rect 355168 238294 355238 238350
rect 355294 238294 355362 238350
rect 355418 238294 355488 238350
rect 355168 238226 355488 238294
rect 355168 238170 355238 238226
rect 355294 238170 355362 238226
rect 355418 238170 355488 238226
rect 355168 238102 355488 238170
rect 355168 238046 355238 238102
rect 355294 238046 355362 238102
rect 355418 238046 355488 238102
rect 355168 237978 355488 238046
rect 355168 237922 355238 237978
rect 355294 237922 355362 237978
rect 355418 237922 355488 237978
rect 355168 237888 355488 237922
rect 385888 238350 386208 238384
rect 385888 238294 385958 238350
rect 386014 238294 386082 238350
rect 386138 238294 386208 238350
rect 385888 238226 386208 238294
rect 385888 238170 385958 238226
rect 386014 238170 386082 238226
rect 386138 238170 386208 238226
rect 385888 238102 386208 238170
rect 385888 238046 385958 238102
rect 386014 238046 386082 238102
rect 386138 238046 386208 238102
rect 385888 237978 386208 238046
rect 385888 237922 385958 237978
rect 386014 237922 386082 237978
rect 386138 237922 386208 237978
rect 385888 237888 386208 237922
rect 416608 238350 416928 238384
rect 416608 238294 416678 238350
rect 416734 238294 416802 238350
rect 416858 238294 416928 238350
rect 416608 238226 416928 238294
rect 416608 238170 416678 238226
rect 416734 238170 416802 238226
rect 416858 238170 416928 238226
rect 416608 238102 416928 238170
rect 416608 238046 416678 238102
rect 416734 238046 416802 238102
rect 416858 238046 416928 238102
rect 416608 237978 416928 238046
rect 416608 237922 416678 237978
rect 416734 237922 416802 237978
rect 416858 237922 416928 237978
rect 416608 237888 416928 237922
rect 339808 226350 340128 226384
rect 339808 226294 339878 226350
rect 339934 226294 340002 226350
rect 340058 226294 340128 226350
rect 339808 226226 340128 226294
rect 339808 226170 339878 226226
rect 339934 226170 340002 226226
rect 340058 226170 340128 226226
rect 339808 226102 340128 226170
rect 339808 226046 339878 226102
rect 339934 226046 340002 226102
rect 340058 226046 340128 226102
rect 339808 225978 340128 226046
rect 339808 225922 339878 225978
rect 339934 225922 340002 225978
rect 340058 225922 340128 225978
rect 339808 225888 340128 225922
rect 370528 226350 370848 226384
rect 370528 226294 370598 226350
rect 370654 226294 370722 226350
rect 370778 226294 370848 226350
rect 370528 226226 370848 226294
rect 370528 226170 370598 226226
rect 370654 226170 370722 226226
rect 370778 226170 370848 226226
rect 370528 226102 370848 226170
rect 370528 226046 370598 226102
rect 370654 226046 370722 226102
rect 370778 226046 370848 226102
rect 370528 225978 370848 226046
rect 370528 225922 370598 225978
rect 370654 225922 370722 225978
rect 370778 225922 370848 225978
rect 370528 225888 370848 225922
rect 401248 226350 401568 226384
rect 401248 226294 401318 226350
rect 401374 226294 401442 226350
rect 401498 226294 401568 226350
rect 401248 226226 401568 226294
rect 401248 226170 401318 226226
rect 401374 226170 401442 226226
rect 401498 226170 401568 226226
rect 401248 226102 401568 226170
rect 401248 226046 401318 226102
rect 401374 226046 401442 226102
rect 401498 226046 401568 226102
rect 401248 225978 401568 226046
rect 401248 225922 401318 225978
rect 401374 225922 401442 225978
rect 401498 225922 401568 225978
rect 401248 225888 401568 225922
rect 324448 220350 324768 220384
rect 324448 220294 324518 220350
rect 324574 220294 324642 220350
rect 324698 220294 324768 220350
rect 324448 220226 324768 220294
rect 324448 220170 324518 220226
rect 324574 220170 324642 220226
rect 324698 220170 324768 220226
rect 324448 220102 324768 220170
rect 324448 220046 324518 220102
rect 324574 220046 324642 220102
rect 324698 220046 324768 220102
rect 324448 219978 324768 220046
rect 324448 219922 324518 219978
rect 324574 219922 324642 219978
rect 324698 219922 324768 219978
rect 324448 219888 324768 219922
rect 355168 220350 355488 220384
rect 355168 220294 355238 220350
rect 355294 220294 355362 220350
rect 355418 220294 355488 220350
rect 355168 220226 355488 220294
rect 355168 220170 355238 220226
rect 355294 220170 355362 220226
rect 355418 220170 355488 220226
rect 355168 220102 355488 220170
rect 355168 220046 355238 220102
rect 355294 220046 355362 220102
rect 355418 220046 355488 220102
rect 355168 219978 355488 220046
rect 355168 219922 355238 219978
rect 355294 219922 355362 219978
rect 355418 219922 355488 219978
rect 355168 219888 355488 219922
rect 385888 220350 386208 220384
rect 385888 220294 385958 220350
rect 386014 220294 386082 220350
rect 386138 220294 386208 220350
rect 385888 220226 386208 220294
rect 385888 220170 385958 220226
rect 386014 220170 386082 220226
rect 386138 220170 386208 220226
rect 385888 220102 386208 220170
rect 385888 220046 385958 220102
rect 386014 220046 386082 220102
rect 386138 220046 386208 220102
rect 385888 219978 386208 220046
rect 385888 219922 385958 219978
rect 386014 219922 386082 219978
rect 386138 219922 386208 219978
rect 385888 219888 386208 219922
rect 416608 220350 416928 220384
rect 416608 220294 416678 220350
rect 416734 220294 416802 220350
rect 416858 220294 416928 220350
rect 416608 220226 416928 220294
rect 416608 220170 416678 220226
rect 416734 220170 416802 220226
rect 416858 220170 416928 220226
rect 416608 220102 416928 220170
rect 416608 220046 416678 220102
rect 416734 220046 416802 220102
rect 416858 220046 416928 220102
rect 416608 219978 416928 220046
rect 416608 219922 416678 219978
rect 416734 219922 416802 219978
rect 416858 219922 416928 219978
rect 416608 219888 416928 219922
rect 339808 208350 340128 208384
rect 339808 208294 339878 208350
rect 339934 208294 340002 208350
rect 340058 208294 340128 208350
rect 339808 208226 340128 208294
rect 339808 208170 339878 208226
rect 339934 208170 340002 208226
rect 340058 208170 340128 208226
rect 339808 208102 340128 208170
rect 339808 208046 339878 208102
rect 339934 208046 340002 208102
rect 340058 208046 340128 208102
rect 339808 207978 340128 208046
rect 339808 207922 339878 207978
rect 339934 207922 340002 207978
rect 340058 207922 340128 207978
rect 339808 207888 340128 207922
rect 370528 208350 370848 208384
rect 370528 208294 370598 208350
rect 370654 208294 370722 208350
rect 370778 208294 370848 208350
rect 370528 208226 370848 208294
rect 370528 208170 370598 208226
rect 370654 208170 370722 208226
rect 370778 208170 370848 208226
rect 370528 208102 370848 208170
rect 370528 208046 370598 208102
rect 370654 208046 370722 208102
rect 370778 208046 370848 208102
rect 370528 207978 370848 208046
rect 370528 207922 370598 207978
rect 370654 207922 370722 207978
rect 370778 207922 370848 207978
rect 370528 207888 370848 207922
rect 401248 208350 401568 208384
rect 401248 208294 401318 208350
rect 401374 208294 401442 208350
rect 401498 208294 401568 208350
rect 401248 208226 401568 208294
rect 401248 208170 401318 208226
rect 401374 208170 401442 208226
rect 401498 208170 401568 208226
rect 401248 208102 401568 208170
rect 401248 208046 401318 208102
rect 401374 208046 401442 208102
rect 401498 208046 401568 208102
rect 401248 207978 401568 208046
rect 401248 207922 401318 207978
rect 401374 207922 401442 207978
rect 401498 207922 401568 207978
rect 401248 207888 401568 207922
rect 324448 202350 324768 202384
rect 324448 202294 324518 202350
rect 324574 202294 324642 202350
rect 324698 202294 324768 202350
rect 324448 202226 324768 202294
rect 324448 202170 324518 202226
rect 324574 202170 324642 202226
rect 324698 202170 324768 202226
rect 324448 202102 324768 202170
rect 324448 202046 324518 202102
rect 324574 202046 324642 202102
rect 324698 202046 324768 202102
rect 324448 201978 324768 202046
rect 324448 201922 324518 201978
rect 324574 201922 324642 201978
rect 324698 201922 324768 201978
rect 324448 201888 324768 201922
rect 355168 202350 355488 202384
rect 355168 202294 355238 202350
rect 355294 202294 355362 202350
rect 355418 202294 355488 202350
rect 355168 202226 355488 202294
rect 355168 202170 355238 202226
rect 355294 202170 355362 202226
rect 355418 202170 355488 202226
rect 355168 202102 355488 202170
rect 355168 202046 355238 202102
rect 355294 202046 355362 202102
rect 355418 202046 355488 202102
rect 355168 201978 355488 202046
rect 355168 201922 355238 201978
rect 355294 201922 355362 201978
rect 355418 201922 355488 201978
rect 355168 201888 355488 201922
rect 385888 202350 386208 202384
rect 385888 202294 385958 202350
rect 386014 202294 386082 202350
rect 386138 202294 386208 202350
rect 385888 202226 386208 202294
rect 385888 202170 385958 202226
rect 386014 202170 386082 202226
rect 386138 202170 386208 202226
rect 385888 202102 386208 202170
rect 385888 202046 385958 202102
rect 386014 202046 386082 202102
rect 386138 202046 386208 202102
rect 385888 201978 386208 202046
rect 385888 201922 385958 201978
rect 386014 201922 386082 201978
rect 386138 201922 386208 201978
rect 385888 201888 386208 201922
rect 416608 202350 416928 202384
rect 416608 202294 416678 202350
rect 416734 202294 416802 202350
rect 416858 202294 416928 202350
rect 416608 202226 416928 202294
rect 416608 202170 416678 202226
rect 416734 202170 416802 202226
rect 416858 202170 416928 202226
rect 416608 202102 416928 202170
rect 416608 202046 416678 202102
rect 416734 202046 416802 202102
rect 416858 202046 416928 202102
rect 416608 201978 416928 202046
rect 416608 201922 416678 201978
rect 416734 201922 416802 201978
rect 416858 201922 416928 201978
rect 416608 201888 416928 201922
rect 339808 190350 340128 190384
rect 339808 190294 339878 190350
rect 339934 190294 340002 190350
rect 340058 190294 340128 190350
rect 339808 190226 340128 190294
rect 339808 190170 339878 190226
rect 339934 190170 340002 190226
rect 340058 190170 340128 190226
rect 339808 190102 340128 190170
rect 339808 190046 339878 190102
rect 339934 190046 340002 190102
rect 340058 190046 340128 190102
rect 339808 189978 340128 190046
rect 339808 189922 339878 189978
rect 339934 189922 340002 189978
rect 340058 189922 340128 189978
rect 339808 189888 340128 189922
rect 370528 190350 370848 190384
rect 370528 190294 370598 190350
rect 370654 190294 370722 190350
rect 370778 190294 370848 190350
rect 370528 190226 370848 190294
rect 370528 190170 370598 190226
rect 370654 190170 370722 190226
rect 370778 190170 370848 190226
rect 370528 190102 370848 190170
rect 370528 190046 370598 190102
rect 370654 190046 370722 190102
rect 370778 190046 370848 190102
rect 370528 189978 370848 190046
rect 370528 189922 370598 189978
rect 370654 189922 370722 189978
rect 370778 189922 370848 189978
rect 370528 189888 370848 189922
rect 401248 190350 401568 190384
rect 401248 190294 401318 190350
rect 401374 190294 401442 190350
rect 401498 190294 401568 190350
rect 401248 190226 401568 190294
rect 401248 190170 401318 190226
rect 401374 190170 401442 190226
rect 401498 190170 401568 190226
rect 401248 190102 401568 190170
rect 401248 190046 401318 190102
rect 401374 190046 401442 190102
rect 401498 190046 401568 190102
rect 401248 189978 401568 190046
rect 401248 189922 401318 189978
rect 401374 189922 401442 189978
rect 401498 189922 401568 189978
rect 401248 189888 401568 189922
rect 324448 184350 324768 184384
rect 324448 184294 324518 184350
rect 324574 184294 324642 184350
rect 324698 184294 324768 184350
rect 324448 184226 324768 184294
rect 324448 184170 324518 184226
rect 324574 184170 324642 184226
rect 324698 184170 324768 184226
rect 324448 184102 324768 184170
rect 324448 184046 324518 184102
rect 324574 184046 324642 184102
rect 324698 184046 324768 184102
rect 324448 183978 324768 184046
rect 324448 183922 324518 183978
rect 324574 183922 324642 183978
rect 324698 183922 324768 183978
rect 324448 183888 324768 183922
rect 355168 184350 355488 184384
rect 355168 184294 355238 184350
rect 355294 184294 355362 184350
rect 355418 184294 355488 184350
rect 355168 184226 355488 184294
rect 355168 184170 355238 184226
rect 355294 184170 355362 184226
rect 355418 184170 355488 184226
rect 355168 184102 355488 184170
rect 355168 184046 355238 184102
rect 355294 184046 355362 184102
rect 355418 184046 355488 184102
rect 355168 183978 355488 184046
rect 355168 183922 355238 183978
rect 355294 183922 355362 183978
rect 355418 183922 355488 183978
rect 355168 183888 355488 183922
rect 385888 184350 386208 184384
rect 385888 184294 385958 184350
rect 386014 184294 386082 184350
rect 386138 184294 386208 184350
rect 385888 184226 386208 184294
rect 385888 184170 385958 184226
rect 386014 184170 386082 184226
rect 386138 184170 386208 184226
rect 385888 184102 386208 184170
rect 385888 184046 385958 184102
rect 386014 184046 386082 184102
rect 386138 184046 386208 184102
rect 385888 183978 386208 184046
rect 385888 183922 385958 183978
rect 386014 183922 386082 183978
rect 386138 183922 386208 183978
rect 385888 183888 386208 183922
rect 416608 184350 416928 184384
rect 416608 184294 416678 184350
rect 416734 184294 416802 184350
rect 416858 184294 416928 184350
rect 416608 184226 416928 184294
rect 416608 184170 416678 184226
rect 416734 184170 416802 184226
rect 416858 184170 416928 184226
rect 416608 184102 416928 184170
rect 416608 184046 416678 184102
rect 416734 184046 416802 184102
rect 416858 184046 416928 184102
rect 416608 183978 416928 184046
rect 416608 183922 416678 183978
rect 416734 183922 416802 183978
rect 416858 183922 416928 183978
rect 416608 183888 416928 183922
rect 339808 172350 340128 172384
rect 339808 172294 339878 172350
rect 339934 172294 340002 172350
rect 340058 172294 340128 172350
rect 339808 172226 340128 172294
rect 339808 172170 339878 172226
rect 339934 172170 340002 172226
rect 340058 172170 340128 172226
rect 339808 172102 340128 172170
rect 339808 172046 339878 172102
rect 339934 172046 340002 172102
rect 340058 172046 340128 172102
rect 339808 171978 340128 172046
rect 339808 171922 339878 171978
rect 339934 171922 340002 171978
rect 340058 171922 340128 171978
rect 339808 171888 340128 171922
rect 370528 172350 370848 172384
rect 370528 172294 370598 172350
rect 370654 172294 370722 172350
rect 370778 172294 370848 172350
rect 370528 172226 370848 172294
rect 370528 172170 370598 172226
rect 370654 172170 370722 172226
rect 370778 172170 370848 172226
rect 370528 172102 370848 172170
rect 370528 172046 370598 172102
rect 370654 172046 370722 172102
rect 370778 172046 370848 172102
rect 370528 171978 370848 172046
rect 370528 171922 370598 171978
rect 370654 171922 370722 171978
rect 370778 171922 370848 171978
rect 370528 171888 370848 171922
rect 401248 172350 401568 172384
rect 401248 172294 401318 172350
rect 401374 172294 401442 172350
rect 401498 172294 401568 172350
rect 401248 172226 401568 172294
rect 401248 172170 401318 172226
rect 401374 172170 401442 172226
rect 401498 172170 401568 172226
rect 401248 172102 401568 172170
rect 401248 172046 401318 172102
rect 401374 172046 401442 172102
rect 401498 172046 401568 172102
rect 401248 171978 401568 172046
rect 401248 171922 401318 171978
rect 401374 171922 401442 171978
rect 401498 171922 401568 171978
rect 401248 171888 401568 171922
rect 324448 166350 324768 166384
rect 324448 166294 324518 166350
rect 324574 166294 324642 166350
rect 324698 166294 324768 166350
rect 324448 166226 324768 166294
rect 324448 166170 324518 166226
rect 324574 166170 324642 166226
rect 324698 166170 324768 166226
rect 324448 166102 324768 166170
rect 324448 166046 324518 166102
rect 324574 166046 324642 166102
rect 324698 166046 324768 166102
rect 324448 165978 324768 166046
rect 324448 165922 324518 165978
rect 324574 165922 324642 165978
rect 324698 165922 324768 165978
rect 324448 165888 324768 165922
rect 355168 166350 355488 166384
rect 355168 166294 355238 166350
rect 355294 166294 355362 166350
rect 355418 166294 355488 166350
rect 355168 166226 355488 166294
rect 355168 166170 355238 166226
rect 355294 166170 355362 166226
rect 355418 166170 355488 166226
rect 355168 166102 355488 166170
rect 355168 166046 355238 166102
rect 355294 166046 355362 166102
rect 355418 166046 355488 166102
rect 355168 165978 355488 166046
rect 355168 165922 355238 165978
rect 355294 165922 355362 165978
rect 355418 165922 355488 165978
rect 355168 165888 355488 165922
rect 385888 166350 386208 166384
rect 385888 166294 385958 166350
rect 386014 166294 386082 166350
rect 386138 166294 386208 166350
rect 385888 166226 386208 166294
rect 385888 166170 385958 166226
rect 386014 166170 386082 166226
rect 386138 166170 386208 166226
rect 385888 166102 386208 166170
rect 385888 166046 385958 166102
rect 386014 166046 386082 166102
rect 386138 166046 386208 166102
rect 385888 165978 386208 166046
rect 385888 165922 385958 165978
rect 386014 165922 386082 165978
rect 386138 165922 386208 165978
rect 385888 165888 386208 165922
rect 416608 166350 416928 166384
rect 416608 166294 416678 166350
rect 416734 166294 416802 166350
rect 416858 166294 416928 166350
rect 416608 166226 416928 166294
rect 416608 166170 416678 166226
rect 416734 166170 416802 166226
rect 416858 166170 416928 166226
rect 416608 166102 416928 166170
rect 416608 166046 416678 166102
rect 416734 166046 416802 166102
rect 416858 166046 416928 166102
rect 416608 165978 416928 166046
rect 416608 165922 416678 165978
rect 416734 165922 416802 165978
rect 416858 165922 416928 165978
rect 416608 165888 416928 165922
rect 339808 154350 340128 154384
rect 339808 154294 339878 154350
rect 339934 154294 340002 154350
rect 340058 154294 340128 154350
rect 339808 154226 340128 154294
rect 339808 154170 339878 154226
rect 339934 154170 340002 154226
rect 340058 154170 340128 154226
rect 339808 154102 340128 154170
rect 339808 154046 339878 154102
rect 339934 154046 340002 154102
rect 340058 154046 340128 154102
rect 339808 153978 340128 154046
rect 339808 153922 339878 153978
rect 339934 153922 340002 153978
rect 340058 153922 340128 153978
rect 339808 153888 340128 153922
rect 370528 154350 370848 154384
rect 370528 154294 370598 154350
rect 370654 154294 370722 154350
rect 370778 154294 370848 154350
rect 370528 154226 370848 154294
rect 370528 154170 370598 154226
rect 370654 154170 370722 154226
rect 370778 154170 370848 154226
rect 370528 154102 370848 154170
rect 370528 154046 370598 154102
rect 370654 154046 370722 154102
rect 370778 154046 370848 154102
rect 370528 153978 370848 154046
rect 370528 153922 370598 153978
rect 370654 153922 370722 153978
rect 370778 153922 370848 153978
rect 370528 153888 370848 153922
rect 401248 154350 401568 154384
rect 401248 154294 401318 154350
rect 401374 154294 401442 154350
rect 401498 154294 401568 154350
rect 401248 154226 401568 154294
rect 401248 154170 401318 154226
rect 401374 154170 401442 154226
rect 401498 154170 401568 154226
rect 401248 154102 401568 154170
rect 401248 154046 401318 154102
rect 401374 154046 401442 154102
rect 401498 154046 401568 154102
rect 401248 153978 401568 154046
rect 401248 153922 401318 153978
rect 401374 153922 401442 153978
rect 401498 153922 401568 153978
rect 401248 153888 401568 153922
rect 324448 148350 324768 148384
rect 324448 148294 324518 148350
rect 324574 148294 324642 148350
rect 324698 148294 324768 148350
rect 324448 148226 324768 148294
rect 324448 148170 324518 148226
rect 324574 148170 324642 148226
rect 324698 148170 324768 148226
rect 324448 148102 324768 148170
rect 324448 148046 324518 148102
rect 324574 148046 324642 148102
rect 324698 148046 324768 148102
rect 324448 147978 324768 148046
rect 324448 147922 324518 147978
rect 324574 147922 324642 147978
rect 324698 147922 324768 147978
rect 324448 147888 324768 147922
rect 355168 148350 355488 148384
rect 355168 148294 355238 148350
rect 355294 148294 355362 148350
rect 355418 148294 355488 148350
rect 355168 148226 355488 148294
rect 355168 148170 355238 148226
rect 355294 148170 355362 148226
rect 355418 148170 355488 148226
rect 355168 148102 355488 148170
rect 355168 148046 355238 148102
rect 355294 148046 355362 148102
rect 355418 148046 355488 148102
rect 355168 147978 355488 148046
rect 355168 147922 355238 147978
rect 355294 147922 355362 147978
rect 355418 147922 355488 147978
rect 355168 147888 355488 147922
rect 385888 148350 386208 148384
rect 385888 148294 385958 148350
rect 386014 148294 386082 148350
rect 386138 148294 386208 148350
rect 385888 148226 386208 148294
rect 385888 148170 385958 148226
rect 386014 148170 386082 148226
rect 386138 148170 386208 148226
rect 385888 148102 386208 148170
rect 385888 148046 385958 148102
rect 386014 148046 386082 148102
rect 386138 148046 386208 148102
rect 385888 147978 386208 148046
rect 385888 147922 385958 147978
rect 386014 147922 386082 147978
rect 386138 147922 386208 147978
rect 385888 147888 386208 147922
rect 416608 148350 416928 148384
rect 416608 148294 416678 148350
rect 416734 148294 416802 148350
rect 416858 148294 416928 148350
rect 416608 148226 416928 148294
rect 416608 148170 416678 148226
rect 416734 148170 416802 148226
rect 416858 148170 416928 148226
rect 416608 148102 416928 148170
rect 416608 148046 416678 148102
rect 416734 148046 416802 148102
rect 416858 148046 416928 148102
rect 416608 147978 416928 148046
rect 416608 147922 416678 147978
rect 416734 147922 416802 147978
rect 416858 147922 416928 147978
rect 416608 147888 416928 147922
rect 339808 136350 340128 136384
rect 339808 136294 339878 136350
rect 339934 136294 340002 136350
rect 340058 136294 340128 136350
rect 339808 136226 340128 136294
rect 339808 136170 339878 136226
rect 339934 136170 340002 136226
rect 340058 136170 340128 136226
rect 339808 136102 340128 136170
rect 339808 136046 339878 136102
rect 339934 136046 340002 136102
rect 340058 136046 340128 136102
rect 339808 135978 340128 136046
rect 339808 135922 339878 135978
rect 339934 135922 340002 135978
rect 340058 135922 340128 135978
rect 339808 135888 340128 135922
rect 370528 136350 370848 136384
rect 370528 136294 370598 136350
rect 370654 136294 370722 136350
rect 370778 136294 370848 136350
rect 370528 136226 370848 136294
rect 370528 136170 370598 136226
rect 370654 136170 370722 136226
rect 370778 136170 370848 136226
rect 370528 136102 370848 136170
rect 370528 136046 370598 136102
rect 370654 136046 370722 136102
rect 370778 136046 370848 136102
rect 370528 135978 370848 136046
rect 370528 135922 370598 135978
rect 370654 135922 370722 135978
rect 370778 135922 370848 135978
rect 370528 135888 370848 135922
rect 401248 136350 401568 136384
rect 401248 136294 401318 136350
rect 401374 136294 401442 136350
rect 401498 136294 401568 136350
rect 401248 136226 401568 136294
rect 401248 136170 401318 136226
rect 401374 136170 401442 136226
rect 401498 136170 401568 136226
rect 401248 136102 401568 136170
rect 401248 136046 401318 136102
rect 401374 136046 401442 136102
rect 401498 136046 401568 136102
rect 401248 135978 401568 136046
rect 401248 135922 401318 135978
rect 401374 135922 401442 135978
rect 401498 135922 401568 135978
rect 401248 135888 401568 135922
rect 324448 130350 324768 130384
rect 324448 130294 324518 130350
rect 324574 130294 324642 130350
rect 324698 130294 324768 130350
rect 324448 130226 324768 130294
rect 324448 130170 324518 130226
rect 324574 130170 324642 130226
rect 324698 130170 324768 130226
rect 324448 130102 324768 130170
rect 324448 130046 324518 130102
rect 324574 130046 324642 130102
rect 324698 130046 324768 130102
rect 324448 129978 324768 130046
rect 324448 129922 324518 129978
rect 324574 129922 324642 129978
rect 324698 129922 324768 129978
rect 324448 129888 324768 129922
rect 355168 130350 355488 130384
rect 355168 130294 355238 130350
rect 355294 130294 355362 130350
rect 355418 130294 355488 130350
rect 355168 130226 355488 130294
rect 355168 130170 355238 130226
rect 355294 130170 355362 130226
rect 355418 130170 355488 130226
rect 355168 130102 355488 130170
rect 355168 130046 355238 130102
rect 355294 130046 355362 130102
rect 355418 130046 355488 130102
rect 355168 129978 355488 130046
rect 355168 129922 355238 129978
rect 355294 129922 355362 129978
rect 355418 129922 355488 129978
rect 355168 129888 355488 129922
rect 385888 130350 386208 130384
rect 385888 130294 385958 130350
rect 386014 130294 386082 130350
rect 386138 130294 386208 130350
rect 385888 130226 386208 130294
rect 385888 130170 385958 130226
rect 386014 130170 386082 130226
rect 386138 130170 386208 130226
rect 385888 130102 386208 130170
rect 385888 130046 385958 130102
rect 386014 130046 386082 130102
rect 386138 130046 386208 130102
rect 385888 129978 386208 130046
rect 385888 129922 385958 129978
rect 386014 129922 386082 129978
rect 386138 129922 386208 129978
rect 385888 129888 386208 129922
rect 416608 130350 416928 130384
rect 416608 130294 416678 130350
rect 416734 130294 416802 130350
rect 416858 130294 416928 130350
rect 416608 130226 416928 130294
rect 416608 130170 416678 130226
rect 416734 130170 416802 130226
rect 416858 130170 416928 130226
rect 416608 130102 416928 130170
rect 416608 130046 416678 130102
rect 416734 130046 416802 130102
rect 416858 130046 416928 130102
rect 416608 129978 416928 130046
rect 416608 129922 416678 129978
rect 416734 129922 416802 129978
rect 416858 129922 416928 129978
rect 416608 129888 416928 129922
rect 339808 118350 340128 118384
rect 339808 118294 339878 118350
rect 339934 118294 340002 118350
rect 340058 118294 340128 118350
rect 339808 118226 340128 118294
rect 339808 118170 339878 118226
rect 339934 118170 340002 118226
rect 340058 118170 340128 118226
rect 339808 118102 340128 118170
rect 339808 118046 339878 118102
rect 339934 118046 340002 118102
rect 340058 118046 340128 118102
rect 339808 117978 340128 118046
rect 339808 117922 339878 117978
rect 339934 117922 340002 117978
rect 340058 117922 340128 117978
rect 339808 117888 340128 117922
rect 370528 118350 370848 118384
rect 370528 118294 370598 118350
rect 370654 118294 370722 118350
rect 370778 118294 370848 118350
rect 370528 118226 370848 118294
rect 370528 118170 370598 118226
rect 370654 118170 370722 118226
rect 370778 118170 370848 118226
rect 370528 118102 370848 118170
rect 370528 118046 370598 118102
rect 370654 118046 370722 118102
rect 370778 118046 370848 118102
rect 370528 117978 370848 118046
rect 370528 117922 370598 117978
rect 370654 117922 370722 117978
rect 370778 117922 370848 117978
rect 370528 117888 370848 117922
rect 401248 118350 401568 118384
rect 401248 118294 401318 118350
rect 401374 118294 401442 118350
rect 401498 118294 401568 118350
rect 401248 118226 401568 118294
rect 401248 118170 401318 118226
rect 401374 118170 401442 118226
rect 401498 118170 401568 118226
rect 401248 118102 401568 118170
rect 401248 118046 401318 118102
rect 401374 118046 401442 118102
rect 401498 118046 401568 118102
rect 401248 117978 401568 118046
rect 401248 117922 401318 117978
rect 401374 117922 401442 117978
rect 401498 117922 401568 117978
rect 401248 117888 401568 117922
rect 324448 112350 324768 112384
rect 324448 112294 324518 112350
rect 324574 112294 324642 112350
rect 324698 112294 324768 112350
rect 324448 112226 324768 112294
rect 324448 112170 324518 112226
rect 324574 112170 324642 112226
rect 324698 112170 324768 112226
rect 324448 112102 324768 112170
rect 324448 112046 324518 112102
rect 324574 112046 324642 112102
rect 324698 112046 324768 112102
rect 324448 111978 324768 112046
rect 324448 111922 324518 111978
rect 324574 111922 324642 111978
rect 324698 111922 324768 111978
rect 324448 111888 324768 111922
rect 355168 112350 355488 112384
rect 355168 112294 355238 112350
rect 355294 112294 355362 112350
rect 355418 112294 355488 112350
rect 355168 112226 355488 112294
rect 355168 112170 355238 112226
rect 355294 112170 355362 112226
rect 355418 112170 355488 112226
rect 355168 112102 355488 112170
rect 355168 112046 355238 112102
rect 355294 112046 355362 112102
rect 355418 112046 355488 112102
rect 355168 111978 355488 112046
rect 355168 111922 355238 111978
rect 355294 111922 355362 111978
rect 355418 111922 355488 111978
rect 355168 111888 355488 111922
rect 385888 112350 386208 112384
rect 385888 112294 385958 112350
rect 386014 112294 386082 112350
rect 386138 112294 386208 112350
rect 385888 112226 386208 112294
rect 385888 112170 385958 112226
rect 386014 112170 386082 112226
rect 386138 112170 386208 112226
rect 385888 112102 386208 112170
rect 385888 112046 385958 112102
rect 386014 112046 386082 112102
rect 386138 112046 386208 112102
rect 385888 111978 386208 112046
rect 385888 111922 385958 111978
rect 386014 111922 386082 111978
rect 386138 111922 386208 111978
rect 385888 111888 386208 111922
rect 416608 112350 416928 112384
rect 416608 112294 416678 112350
rect 416734 112294 416802 112350
rect 416858 112294 416928 112350
rect 416608 112226 416928 112294
rect 416608 112170 416678 112226
rect 416734 112170 416802 112226
rect 416858 112170 416928 112226
rect 416608 112102 416928 112170
rect 416608 112046 416678 112102
rect 416734 112046 416802 112102
rect 416858 112046 416928 112102
rect 416608 111978 416928 112046
rect 416608 111922 416678 111978
rect 416734 111922 416802 111978
rect 416858 111922 416928 111978
rect 416608 111888 416928 111922
rect 321692 83346 321748 83356
rect 347058 100350 347678 102954
rect 347058 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 347678 100350
rect 347058 100226 347678 100294
rect 347058 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 347678 100226
rect 347058 100102 347678 100170
rect 347058 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 347678 100102
rect 347058 99978 347678 100046
rect 347058 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 347678 99978
rect 317436 83032 317492 83042
rect 316338 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 316958 82350
rect 316338 82226 316958 82294
rect 316338 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 316958 82226
rect 316338 82102 316958 82170
rect 316338 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 316958 82102
rect 316338 81978 316958 82046
rect 316338 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 316958 81978
rect 316338 79630 316958 81922
rect 347058 82350 347678 99922
rect 347058 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 347678 82350
rect 347058 82226 347678 82294
rect 347058 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 347678 82226
rect 347058 82102 347678 82170
rect 347058 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 347678 82102
rect 347058 81978 347678 82046
rect 347058 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 347678 81978
rect 347058 79630 347678 81922
rect 377778 100350 378398 102954
rect 377778 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 378398 100350
rect 377778 100226 378398 100294
rect 377778 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 378398 100226
rect 377778 100102 378398 100170
rect 377778 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 378398 100102
rect 377778 99978 378398 100046
rect 377778 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 378398 99978
rect 377778 82350 378398 99922
rect 377778 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 378398 82350
rect 377778 82226 378398 82294
rect 377778 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 378398 82226
rect 377778 82102 378398 82170
rect 377778 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 378398 82102
rect 377778 81978 378398 82046
rect 377778 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 378398 81978
rect 377778 79630 378398 81922
rect 408498 100350 409118 102954
rect 408498 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 409118 100350
rect 408498 100226 409118 100294
rect 408498 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 409118 100226
rect 408498 100102 409118 100170
rect 408498 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 409118 100102
rect 408498 99978 409118 100046
rect 408498 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 409118 99978
rect 408498 82350 409118 99922
rect 408498 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 409118 82350
rect 408498 82226 409118 82294
rect 408498 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 409118 82226
rect 408498 82102 409118 82170
rect 408498 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 409118 82102
rect 408498 81978 409118 82046
rect 408498 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 409118 81978
rect 408498 79630 409118 81922
rect 419132 81508 419188 321692
rect 419244 92932 419300 325052
rect 419356 110852 419412 328412
rect 419468 139524 419524 333788
rect 419580 322420 419636 322430
rect 419580 170548 419636 322364
rect 419692 268548 419748 357980
rect 419804 282884 419860 360668
rect 419916 307972 419972 365372
rect 420812 364084 420868 364094
rect 419916 307906 419972 307916
rect 420700 361396 420756 361406
rect 420700 286468 420756 361340
rect 420812 331940 420868 364028
rect 420924 358148 420980 374780
rect 422604 374164 422660 374174
rect 421036 370804 421092 370814
rect 421036 360388 421092 370748
rect 421036 360322 421092 360332
rect 422492 362068 422548 362078
rect 420924 358082 420980 358092
rect 421596 356020 421652 356030
rect 420924 351316 420980 351326
rect 420924 336868 420980 351260
rect 420924 336802 420980 336812
rect 421484 337204 421540 337214
rect 420812 331874 420868 331884
rect 421372 334516 421428 334526
rect 421260 331828 421316 331838
rect 421036 325780 421092 325790
rect 420700 286402 420756 286412
rect 420812 317716 420868 317726
rect 419804 282818 419860 282828
rect 420476 285684 420532 285694
rect 419692 268482 419748 268492
rect 419580 170482 419636 170492
rect 419468 139458 419524 139468
rect 419356 110786 419412 110796
rect 419244 92866 419300 92876
rect 419132 81442 419188 81452
rect 314972 78892 315028 78902
rect 302352 76350 302672 76384
rect 302352 76294 302422 76350
rect 302478 76294 302546 76350
rect 302602 76294 302672 76350
rect 302352 76226 302672 76294
rect 302352 76170 302422 76226
rect 302478 76170 302546 76226
rect 302602 76170 302672 76226
rect 302352 76102 302672 76170
rect 302352 76046 302422 76102
rect 302478 76046 302546 76102
rect 302602 76046 302672 76102
rect 302352 75978 302672 76046
rect 302352 75922 302422 75978
rect 302478 75922 302546 75978
rect 302602 75922 302672 75978
rect 302352 75888 302672 75922
rect 333072 76350 333392 76384
rect 333072 76294 333142 76350
rect 333198 76294 333266 76350
rect 333322 76294 333392 76350
rect 333072 76226 333392 76294
rect 333072 76170 333142 76226
rect 333198 76170 333266 76226
rect 333322 76170 333392 76226
rect 333072 76102 333392 76170
rect 333072 76046 333142 76102
rect 333198 76046 333266 76102
rect 333322 76046 333392 76102
rect 333072 75978 333392 76046
rect 333072 75922 333142 75978
rect 333198 75922 333266 75978
rect 333322 75922 333392 75978
rect 333072 75888 333392 75922
rect 363792 76350 364112 76384
rect 363792 76294 363862 76350
rect 363918 76294 363986 76350
rect 364042 76294 364112 76350
rect 363792 76226 364112 76294
rect 363792 76170 363862 76226
rect 363918 76170 363986 76226
rect 364042 76170 364112 76226
rect 363792 76102 364112 76170
rect 363792 76046 363862 76102
rect 363918 76046 363986 76102
rect 364042 76046 364112 76102
rect 363792 75978 364112 76046
rect 363792 75922 363862 75978
rect 363918 75922 363986 75978
rect 364042 75922 364112 75978
rect 363792 75888 364112 75922
rect 394512 76350 394832 76384
rect 394512 76294 394582 76350
rect 394638 76294 394706 76350
rect 394762 76294 394832 76350
rect 394512 76226 394832 76294
rect 394512 76170 394582 76226
rect 394638 76170 394706 76226
rect 394762 76170 394832 76226
rect 394512 76102 394832 76170
rect 394512 76046 394582 76102
rect 394638 76046 394706 76102
rect 394762 76046 394832 76102
rect 394512 75978 394832 76046
rect 394512 75922 394582 75978
rect 394638 75922 394706 75978
rect 394762 75922 394832 75978
rect 394512 75888 394832 75922
rect 274092 74032 274148 74042
rect 273644 69712 273700 69722
rect 286992 64350 287312 64384
rect 286992 64294 287062 64350
rect 287118 64294 287186 64350
rect 287242 64294 287312 64350
rect 286992 64226 287312 64294
rect 286992 64170 287062 64226
rect 287118 64170 287186 64226
rect 287242 64170 287312 64226
rect 286992 64102 287312 64170
rect 286992 64046 287062 64102
rect 287118 64046 287186 64102
rect 287242 64046 287312 64102
rect 286992 63978 287312 64046
rect 286992 63922 287062 63978
rect 287118 63922 287186 63978
rect 287242 63922 287312 63978
rect 286992 63888 287312 63922
rect 317712 64350 318032 64384
rect 317712 64294 317782 64350
rect 317838 64294 317906 64350
rect 317962 64294 318032 64350
rect 317712 64226 318032 64294
rect 317712 64170 317782 64226
rect 317838 64170 317906 64226
rect 317962 64170 318032 64226
rect 317712 64102 318032 64170
rect 317712 64046 317782 64102
rect 317838 64046 317906 64102
rect 317962 64046 318032 64102
rect 317712 63978 318032 64046
rect 317712 63922 317782 63978
rect 317838 63922 317906 63978
rect 317962 63922 318032 63978
rect 317712 63888 318032 63922
rect 348432 64350 348752 64384
rect 348432 64294 348502 64350
rect 348558 64294 348626 64350
rect 348682 64294 348752 64350
rect 348432 64226 348752 64294
rect 348432 64170 348502 64226
rect 348558 64170 348626 64226
rect 348682 64170 348752 64226
rect 348432 64102 348752 64170
rect 348432 64046 348502 64102
rect 348558 64046 348626 64102
rect 348682 64046 348752 64102
rect 348432 63978 348752 64046
rect 348432 63922 348502 63978
rect 348558 63922 348626 63978
rect 348682 63922 348752 63978
rect 348432 63888 348752 63922
rect 379152 64350 379472 64384
rect 379152 64294 379222 64350
rect 379278 64294 379346 64350
rect 379402 64294 379472 64350
rect 379152 64226 379472 64294
rect 379152 64170 379222 64226
rect 379278 64170 379346 64226
rect 379402 64170 379472 64226
rect 379152 64102 379472 64170
rect 379152 64046 379222 64102
rect 379278 64046 379346 64102
rect 379402 64046 379472 64102
rect 379152 63978 379472 64046
rect 379152 63922 379222 63978
rect 379278 63922 379346 63978
rect 379402 63922 379472 63978
rect 379152 63888 379472 63922
rect 409872 64350 410192 64384
rect 409872 64294 409942 64350
rect 409998 64294 410066 64350
rect 410122 64294 410192 64350
rect 409872 64226 410192 64294
rect 409872 64170 409942 64226
rect 409998 64170 410066 64226
rect 410122 64170 410192 64226
rect 409872 64102 410192 64170
rect 409872 64046 409942 64102
rect 409998 64046 410066 64102
rect 410122 64046 410192 64102
rect 409872 63978 410192 64046
rect 409872 63922 409942 63978
rect 409998 63922 410066 63978
rect 410122 63922 410192 63978
rect 409872 63888 410192 63922
rect 302352 58350 302672 58384
rect 302352 58294 302422 58350
rect 302478 58294 302546 58350
rect 302602 58294 302672 58350
rect 302352 58226 302672 58294
rect 302352 58170 302422 58226
rect 302478 58170 302546 58226
rect 302602 58170 302672 58226
rect 302352 58102 302672 58170
rect 302352 58046 302422 58102
rect 302478 58046 302546 58102
rect 302602 58046 302672 58102
rect 302352 57978 302672 58046
rect 302352 57922 302422 57978
rect 302478 57922 302546 57978
rect 302602 57922 302672 57978
rect 302352 57888 302672 57922
rect 333072 58350 333392 58384
rect 333072 58294 333142 58350
rect 333198 58294 333266 58350
rect 333322 58294 333392 58350
rect 333072 58226 333392 58294
rect 333072 58170 333142 58226
rect 333198 58170 333266 58226
rect 333322 58170 333392 58226
rect 333072 58102 333392 58170
rect 333072 58046 333142 58102
rect 333198 58046 333266 58102
rect 333322 58046 333392 58102
rect 333072 57978 333392 58046
rect 333072 57922 333142 57978
rect 333198 57922 333266 57978
rect 333322 57922 333392 57978
rect 333072 57888 333392 57922
rect 363792 58350 364112 58384
rect 363792 58294 363862 58350
rect 363918 58294 363986 58350
rect 364042 58294 364112 58350
rect 363792 58226 364112 58294
rect 363792 58170 363862 58226
rect 363918 58170 363986 58226
rect 364042 58170 364112 58226
rect 363792 58102 364112 58170
rect 363792 58046 363862 58102
rect 363918 58046 363986 58102
rect 364042 58046 364112 58102
rect 363792 57978 364112 58046
rect 363792 57922 363862 57978
rect 363918 57922 363986 57978
rect 364042 57922 364112 57978
rect 363792 57888 364112 57922
rect 394512 58350 394832 58384
rect 394512 58294 394582 58350
rect 394638 58294 394706 58350
rect 394762 58294 394832 58350
rect 394512 58226 394832 58294
rect 394512 58170 394582 58226
rect 394638 58170 394706 58226
rect 394762 58170 394832 58226
rect 394512 58102 394832 58170
rect 394512 58046 394582 58102
rect 394638 58046 394706 58102
rect 394762 58046 394832 58102
rect 394512 57978 394832 58046
rect 394512 57922 394582 57978
rect 394638 57922 394706 57978
rect 394762 57922 394832 57978
rect 394512 57888 394832 57922
rect 286992 46350 287312 46384
rect 286992 46294 287062 46350
rect 287118 46294 287186 46350
rect 287242 46294 287312 46350
rect 286992 46226 287312 46294
rect 286992 46170 287062 46226
rect 287118 46170 287186 46226
rect 287242 46170 287312 46226
rect 286992 46102 287312 46170
rect 286992 46046 287062 46102
rect 287118 46046 287186 46102
rect 287242 46046 287312 46102
rect 286992 45978 287312 46046
rect 286992 45922 287062 45978
rect 287118 45922 287186 45978
rect 287242 45922 287312 45978
rect 286992 45888 287312 45922
rect 317712 46350 318032 46384
rect 317712 46294 317782 46350
rect 317838 46294 317906 46350
rect 317962 46294 318032 46350
rect 317712 46226 318032 46294
rect 317712 46170 317782 46226
rect 317838 46170 317906 46226
rect 317962 46170 318032 46226
rect 317712 46102 318032 46170
rect 317712 46046 317782 46102
rect 317838 46046 317906 46102
rect 317962 46046 318032 46102
rect 317712 45978 318032 46046
rect 317712 45922 317782 45978
rect 317838 45922 317906 45978
rect 317962 45922 318032 45978
rect 317712 45888 318032 45922
rect 348432 46350 348752 46384
rect 348432 46294 348502 46350
rect 348558 46294 348626 46350
rect 348682 46294 348752 46350
rect 348432 46226 348752 46294
rect 348432 46170 348502 46226
rect 348558 46170 348626 46226
rect 348682 46170 348752 46226
rect 348432 46102 348752 46170
rect 348432 46046 348502 46102
rect 348558 46046 348626 46102
rect 348682 46046 348752 46102
rect 348432 45978 348752 46046
rect 348432 45922 348502 45978
rect 348558 45922 348626 45978
rect 348682 45922 348752 45978
rect 348432 45888 348752 45922
rect 379152 46350 379472 46384
rect 379152 46294 379222 46350
rect 379278 46294 379346 46350
rect 379402 46294 379472 46350
rect 379152 46226 379472 46294
rect 379152 46170 379222 46226
rect 379278 46170 379346 46226
rect 379402 46170 379472 46226
rect 379152 46102 379472 46170
rect 379152 46046 379222 46102
rect 379278 46046 379346 46102
rect 379402 46046 379472 46102
rect 379152 45978 379472 46046
rect 379152 45922 379222 45978
rect 379278 45922 379346 45978
rect 379402 45922 379472 45978
rect 379152 45888 379472 45922
rect 409872 46350 410192 46384
rect 409872 46294 409942 46350
rect 409998 46294 410066 46350
rect 410122 46294 410192 46350
rect 409872 46226 410192 46294
rect 409872 46170 409942 46226
rect 409998 46170 410066 46226
rect 410122 46170 410192 46226
rect 409872 46102 410192 46170
rect 409872 46046 409942 46102
rect 409998 46046 410066 46102
rect 410122 46046 410192 46102
rect 409872 45978 410192 46046
rect 409872 45922 409942 45978
rect 409998 45922 410066 45978
rect 410122 45922 410192 45978
rect 409872 45888 410192 45922
rect 302352 40350 302672 40384
rect 302352 40294 302422 40350
rect 302478 40294 302546 40350
rect 302602 40294 302672 40350
rect 302352 40226 302672 40294
rect 302352 40170 302422 40226
rect 302478 40170 302546 40226
rect 302602 40170 302672 40226
rect 302352 40102 302672 40170
rect 302352 40046 302422 40102
rect 302478 40046 302546 40102
rect 302602 40046 302672 40102
rect 302352 39978 302672 40046
rect 302352 39922 302422 39978
rect 302478 39922 302546 39978
rect 302602 39922 302672 39978
rect 302352 39888 302672 39922
rect 333072 40350 333392 40384
rect 333072 40294 333142 40350
rect 333198 40294 333266 40350
rect 333322 40294 333392 40350
rect 333072 40226 333392 40294
rect 333072 40170 333142 40226
rect 333198 40170 333266 40226
rect 333322 40170 333392 40226
rect 333072 40102 333392 40170
rect 333072 40046 333142 40102
rect 333198 40046 333266 40102
rect 333322 40046 333392 40102
rect 333072 39978 333392 40046
rect 333072 39922 333142 39978
rect 333198 39922 333266 39978
rect 333322 39922 333392 39978
rect 333072 39888 333392 39922
rect 363792 40350 364112 40384
rect 363792 40294 363862 40350
rect 363918 40294 363986 40350
rect 364042 40294 364112 40350
rect 363792 40226 364112 40294
rect 363792 40170 363862 40226
rect 363918 40170 363986 40226
rect 364042 40170 364112 40226
rect 363792 40102 364112 40170
rect 363792 40046 363862 40102
rect 363918 40046 363986 40102
rect 364042 40046 364112 40102
rect 363792 39978 364112 40046
rect 363792 39922 363862 39978
rect 363918 39922 363986 39978
rect 364042 39922 364112 39978
rect 363792 39888 364112 39922
rect 394512 40350 394832 40384
rect 394512 40294 394582 40350
rect 394638 40294 394706 40350
rect 394762 40294 394832 40350
rect 394512 40226 394832 40294
rect 394512 40170 394582 40226
rect 394638 40170 394706 40226
rect 394762 40170 394832 40226
rect 394512 40102 394832 40170
rect 394512 40046 394582 40102
rect 394638 40046 394706 40102
rect 394762 40046 394832 40102
rect 394512 39978 394832 40046
rect 394512 39922 394582 39978
rect 394638 39922 394706 39978
rect 394762 39922 394832 39978
rect 394512 39888 394832 39922
rect 286992 28350 287312 28384
rect 286992 28294 287062 28350
rect 287118 28294 287186 28350
rect 287242 28294 287312 28350
rect 286992 28226 287312 28294
rect 286992 28170 287062 28226
rect 287118 28170 287186 28226
rect 287242 28170 287312 28226
rect 286992 28102 287312 28170
rect 286992 28046 287062 28102
rect 287118 28046 287186 28102
rect 287242 28046 287312 28102
rect 286992 27978 287312 28046
rect 286992 27922 287062 27978
rect 287118 27922 287186 27978
rect 287242 27922 287312 27978
rect 286992 27888 287312 27922
rect 317712 28350 318032 28384
rect 317712 28294 317782 28350
rect 317838 28294 317906 28350
rect 317962 28294 318032 28350
rect 317712 28226 318032 28294
rect 317712 28170 317782 28226
rect 317838 28170 317906 28226
rect 317962 28170 318032 28226
rect 317712 28102 318032 28170
rect 317712 28046 317782 28102
rect 317838 28046 317906 28102
rect 317962 28046 318032 28102
rect 317712 27978 318032 28046
rect 317712 27922 317782 27978
rect 317838 27922 317906 27978
rect 317962 27922 318032 27978
rect 317712 27888 318032 27922
rect 348432 28350 348752 28384
rect 348432 28294 348502 28350
rect 348558 28294 348626 28350
rect 348682 28294 348752 28350
rect 348432 28226 348752 28294
rect 348432 28170 348502 28226
rect 348558 28170 348626 28226
rect 348682 28170 348752 28226
rect 348432 28102 348752 28170
rect 348432 28046 348502 28102
rect 348558 28046 348626 28102
rect 348682 28046 348752 28102
rect 348432 27978 348752 28046
rect 348432 27922 348502 27978
rect 348558 27922 348626 27978
rect 348682 27922 348752 27978
rect 348432 27888 348752 27922
rect 379152 28350 379472 28384
rect 379152 28294 379222 28350
rect 379278 28294 379346 28350
rect 379402 28294 379472 28350
rect 379152 28226 379472 28294
rect 379152 28170 379222 28226
rect 379278 28170 379346 28226
rect 379402 28170 379472 28226
rect 379152 28102 379472 28170
rect 379152 28046 379222 28102
rect 379278 28046 379346 28102
rect 379402 28046 379472 28102
rect 379152 27978 379472 28046
rect 379152 27922 379222 27978
rect 379278 27922 379346 27978
rect 379402 27922 379472 27978
rect 379152 27888 379472 27922
rect 409872 28350 410192 28384
rect 409872 28294 409942 28350
rect 409998 28294 410066 28350
rect 410122 28294 410192 28350
rect 409872 28226 410192 28294
rect 409872 28170 409942 28226
rect 409998 28170 410066 28226
rect 410122 28170 410192 28226
rect 409872 28102 410192 28170
rect 409872 28046 409942 28102
rect 409998 28046 410066 28102
rect 410122 28046 410192 28102
rect 409872 27978 410192 28046
rect 409872 27922 409942 27978
rect 409998 27922 410066 27978
rect 410122 27922 410192 27978
rect 409872 27888 410192 27922
rect 302352 22350 302672 22384
rect 302352 22294 302422 22350
rect 302478 22294 302546 22350
rect 302602 22294 302672 22350
rect 302352 22226 302672 22294
rect 302352 22170 302422 22226
rect 302478 22170 302546 22226
rect 302602 22170 302672 22226
rect 302352 22102 302672 22170
rect 302352 22046 302422 22102
rect 302478 22046 302546 22102
rect 302602 22046 302672 22102
rect 302352 21978 302672 22046
rect 302352 21922 302422 21978
rect 302478 21922 302546 21978
rect 302602 21922 302672 21978
rect 302352 21888 302672 21922
rect 333072 22350 333392 22384
rect 333072 22294 333142 22350
rect 333198 22294 333266 22350
rect 333322 22294 333392 22350
rect 333072 22226 333392 22294
rect 333072 22170 333142 22226
rect 333198 22170 333266 22226
rect 333322 22170 333392 22226
rect 333072 22102 333392 22170
rect 333072 22046 333142 22102
rect 333198 22046 333266 22102
rect 333322 22046 333392 22102
rect 333072 21978 333392 22046
rect 333072 21922 333142 21978
rect 333198 21922 333266 21978
rect 333322 21922 333392 21978
rect 333072 21888 333392 21922
rect 363792 22350 364112 22384
rect 363792 22294 363862 22350
rect 363918 22294 363986 22350
rect 364042 22294 364112 22350
rect 363792 22226 364112 22294
rect 363792 22170 363862 22226
rect 363918 22170 363986 22226
rect 364042 22170 364112 22226
rect 363792 22102 364112 22170
rect 363792 22046 363862 22102
rect 363918 22046 363986 22102
rect 364042 22046 364112 22102
rect 363792 21978 364112 22046
rect 363792 21922 363862 21978
rect 363918 21922 363986 21978
rect 364042 21922 364112 21978
rect 363792 21888 364112 21922
rect 394512 22350 394832 22384
rect 394512 22294 394582 22350
rect 394638 22294 394706 22350
rect 394762 22294 394832 22350
rect 394512 22226 394832 22294
rect 394512 22170 394582 22226
rect 394638 22170 394706 22226
rect 394762 22170 394832 22226
rect 394512 22102 394832 22170
rect 394512 22046 394582 22102
rect 394638 22046 394706 22102
rect 394762 22046 394832 22102
rect 394512 21978 394832 22046
rect 394512 21922 394582 21978
rect 394638 21922 394706 21978
rect 394762 21922 394832 21978
rect 394512 21888 394832 21922
rect 273420 20032 273476 20042
rect 273196 19672 273252 19682
rect 272972 19312 273028 19322
rect 273308 17038 273364 17048
rect 272860 16858 272916 16868
rect 272188 16138 272244 16148
rect 270508 13562 270676 13618
rect 272076 15238 272132 15248
rect 270508 13076 270564 13562
rect 270620 13412 270788 13438
rect 270676 13382 270788 13412
rect 270620 13346 270676 13356
rect 270732 13258 270788 13382
rect 270732 13202 271572 13258
rect 270620 13188 270676 13198
rect 270620 13078 270676 13132
rect 270620 13022 271460 13078
rect 270508 13010 270564 13020
rect 270284 12842 270564 12898
rect 270172 12226 270228 12236
rect 270396 12740 270452 12750
rect 270284 11284 270340 11294
rect 270284 10052 270340 11228
rect 270284 9986 270340 9996
rect 270396 2818 270452 12684
rect 270508 7028 270564 12842
rect 270620 12852 270676 12862
rect 270620 8428 270676 12796
rect 271404 8428 271460 13022
rect 271516 12898 271572 13202
rect 271516 12842 271684 12898
rect 270620 8372 271348 8428
rect 271404 8372 271572 8428
rect 270508 6962 270564 6972
rect 270396 2752 270452 2762
rect 269836 2034 269892 2044
rect 271292 478 271348 8372
rect 271516 4788 271572 8372
rect 271628 6356 271684 12842
rect 272076 9716 272132 15182
rect 272076 9650 272132 9660
rect 271628 6290 271684 6300
rect 271516 4722 271572 4732
rect 272188 4228 272244 16082
rect 272860 8428 272916 16802
rect 273196 16318 273252 16328
rect 272972 13798 273028 13808
rect 272972 9940 273028 13742
rect 272972 9874 273028 9884
rect 273084 12538 273140 12548
rect 272860 8372 273028 8428
rect 272972 6692 273028 8372
rect 272972 6626 273028 6636
rect 272188 4162 272244 4172
rect 273084 1540 273140 12482
rect 273196 4676 273252 16262
rect 273308 6916 273364 16982
rect 274092 13618 274148 13628
rect 273308 6850 273364 6860
rect 273420 11818 273476 11828
rect 273196 4610 273252 4620
rect 273420 2998 273476 11762
rect 273868 11638 273924 11648
rect 273868 10164 273924 11582
rect 273868 10098 273924 10108
rect 274092 8260 274148 13562
rect 420476 10500 420532 285628
rect 420476 10434 420532 10444
rect 420588 258692 420644 258702
rect 288988 9658 289044 9668
rect 274092 8194 274148 8204
rect 273420 2932 273476 2942
rect 281898 4350 282518 8578
rect 288988 6244 289044 9602
rect 288988 6178 289044 6188
rect 304108 8484 304164 8494
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 277228 2548 277284 2558
rect 277228 2458 277284 2492
rect 277228 2392 277284 2402
rect 273084 1474 273140 1484
rect 271292 412 271348 422
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 -160 282518 3922
rect 304108 2638 304164 8428
rect 304108 2572 304164 2582
rect 312618 4350 313238 8578
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 343338 4350 343958 8578
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 374058 4350 374678 8578
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 394044 6598 394100 6608
rect 394044 3444 394100 6542
rect 394044 3378 394100 3388
rect 404778 4350 405398 8578
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 420588 4340 420644 258636
rect 420700 91700 420756 91710
rect 420700 9380 420756 91644
rect 420812 85092 420868 317660
rect 420812 85026 420868 85036
rect 420924 315700 420980 315710
rect 420924 83300 420980 315644
rect 421036 96516 421092 325724
rect 421036 96450 421092 96460
rect 421148 298788 421204 298798
rect 420924 83234 420980 83244
rect 421036 86996 421092 87006
rect 420812 81172 420868 81182
rect 420812 67978 420868 81116
rect 420812 67912 420868 67922
rect 421036 9604 421092 86940
rect 421148 82180 421204 298732
rect 421260 128772 421316 331772
rect 421372 143108 421428 334460
rect 421484 173908 421540 337148
rect 421596 257796 421652 355964
rect 422492 330148 422548 362012
rect 422604 357028 422660 374108
rect 422604 356962 422660 356972
rect 423276 343252 423332 343262
rect 423164 340564 423220 340574
rect 423052 337876 423108 337886
rect 422492 330082 422548 330092
rect 422940 332500 422996 332510
rect 422716 329812 422772 329822
rect 422604 327124 422660 327134
rect 421596 257730 421652 257740
rect 422492 320404 422548 320414
rect 421484 173842 421540 173852
rect 421372 143042 421428 143052
rect 421260 128706 421316 128716
rect 422044 90356 422100 90366
rect 421932 87780 421988 87790
rect 421148 82114 421204 82124
rect 421484 87108 421540 87118
rect 421036 9538 421092 9548
rect 420700 9314 420756 9324
rect 421484 7924 421540 87052
rect 421484 7858 421540 7868
rect 421708 86884 421764 86894
rect 420588 4274 420644 4284
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 404778 -160 405398 3922
rect 421708 1652 421764 86828
rect 421820 86772 421876 86782
rect 421820 3332 421876 86716
rect 421932 4228 421988 87724
rect 422044 8036 422100 90300
rect 422268 86548 422324 86558
rect 422044 7970 422100 7980
rect 422156 83412 422212 83422
rect 421932 4162 421988 4172
rect 421820 3266 421876 3276
rect 422156 3108 422212 83356
rect 422268 7812 422324 86492
rect 422492 78372 422548 320348
rect 422604 103684 422660 327068
rect 422716 120148 422772 329756
rect 422716 120082 422772 120092
rect 422828 326452 422884 326462
rect 422828 105028 422884 326396
rect 422940 132356 422996 332444
rect 423052 161028 423108 337820
rect 423164 175364 423220 340508
rect 423276 189700 423332 343196
rect 423500 301078 423556 301088
rect 423276 189634 423332 189644
rect 423388 298340 423444 298350
rect 423164 175298 423220 175308
rect 423052 160962 423108 160972
rect 422940 132290 422996 132300
rect 422828 104962 422884 104972
rect 422604 103618 422660 103628
rect 422492 78306 422548 78316
rect 422268 7746 422324 7756
rect 422156 3042 422212 3052
rect 421708 1586 421764 1596
rect 423388 1540 423444 298284
rect 423500 5908 423556 301022
rect 423724 298900 423780 298910
rect 423612 298564 423668 298574
rect 423612 8148 423668 298508
rect 423724 8260 423780 298844
rect 424172 101998 424228 377132
rect 424396 344596 424452 344606
rect 424284 341236 424340 341246
rect 424284 178948 424340 341180
rect 424396 196868 424452 344540
rect 424508 329140 424564 329150
rect 424508 294868 424564 329084
rect 424508 294802 424564 294812
rect 424620 301924 424676 301934
rect 424620 275716 424676 301868
rect 424620 275650 424676 275660
rect 424396 196802 424452 196812
rect 424284 178882 424340 178892
rect 424172 101932 424228 101942
rect 425068 90244 425124 90254
rect 423724 8194 423780 8204
rect 423836 81060 423892 81070
rect 423612 8082 423668 8092
rect 423500 5842 423556 5852
rect 423836 4228 423892 81004
rect 423948 78260 424004 78270
rect 423948 10388 424004 78204
rect 423948 10322 424004 10332
rect 424172 13438 424228 13448
rect 424172 4900 424228 13382
rect 425068 6132 425124 90188
rect 425740 84196 425796 84206
rect 425628 82292 425684 82302
rect 425232 76350 425552 76384
rect 425232 76294 425302 76350
rect 425358 76294 425426 76350
rect 425482 76294 425552 76350
rect 425232 76226 425552 76294
rect 425232 76170 425302 76226
rect 425358 76170 425426 76226
rect 425482 76170 425552 76226
rect 425232 76102 425552 76170
rect 425232 76046 425302 76102
rect 425358 76046 425426 76102
rect 425482 76046 425552 76102
rect 425232 75978 425552 76046
rect 425232 75922 425302 75978
rect 425358 75922 425426 75978
rect 425482 75922 425552 75978
rect 425232 75888 425552 75922
rect 425232 58350 425552 58384
rect 425232 58294 425302 58350
rect 425358 58294 425426 58350
rect 425482 58294 425552 58350
rect 425232 58226 425552 58294
rect 425232 58170 425302 58226
rect 425358 58170 425426 58226
rect 425482 58170 425552 58226
rect 425232 58102 425552 58170
rect 425232 58046 425302 58102
rect 425358 58046 425426 58102
rect 425482 58046 425552 58102
rect 425232 57978 425552 58046
rect 425232 57922 425302 57978
rect 425358 57922 425426 57978
rect 425482 57922 425552 57978
rect 425232 57888 425552 57922
rect 425232 40350 425552 40384
rect 425232 40294 425302 40350
rect 425358 40294 425426 40350
rect 425482 40294 425552 40350
rect 425232 40226 425552 40294
rect 425232 40170 425302 40226
rect 425358 40170 425426 40226
rect 425482 40170 425552 40226
rect 425232 40102 425552 40170
rect 425232 40046 425302 40102
rect 425358 40046 425426 40102
rect 425482 40046 425552 40102
rect 425232 39978 425552 40046
rect 425232 39922 425302 39978
rect 425358 39922 425426 39978
rect 425482 39922 425552 39978
rect 425232 39888 425552 39922
rect 425232 22350 425552 22384
rect 425232 22294 425302 22350
rect 425358 22294 425426 22350
rect 425482 22294 425552 22350
rect 425232 22226 425552 22294
rect 425232 22170 425302 22226
rect 425358 22170 425426 22226
rect 425482 22170 425552 22226
rect 425232 22102 425552 22170
rect 425232 22046 425302 22102
rect 425358 22046 425426 22102
rect 425482 22046 425552 22102
rect 425232 21978 425552 22046
rect 425232 21922 425302 21978
rect 425358 21922 425426 21978
rect 425482 21922 425552 21978
rect 425232 21888 425552 21922
rect 425628 6356 425684 82236
rect 425740 10500 425796 84140
rect 425852 79858 425908 378812
rect 425964 370132 426020 370142
rect 425964 341908 426020 370076
rect 426412 349300 426468 349310
rect 425964 341842 426020 341852
rect 426300 346612 426356 346622
rect 426188 339220 426244 339230
rect 425964 324436 426020 324446
rect 425964 89348 426020 324380
rect 425964 89282 426020 89292
rect 426076 318388 426132 318398
rect 426076 86548 426132 318332
rect 426188 168196 426244 339164
rect 426300 207620 426356 346556
rect 426412 221956 426468 349244
rect 426412 221890 426468 221900
rect 426748 298676 426804 298686
rect 426300 207554 426356 207564
rect 426188 168130 426244 168140
rect 426076 86482 426132 86492
rect 425852 79792 425908 79802
rect 425740 10434 425796 10444
rect 426748 9268 426804 298620
rect 426748 9202 426804 9212
rect 426860 93380 426916 93390
rect 425628 6290 425684 6300
rect 426860 6244 426916 93324
rect 426972 91588 427028 91598
rect 426972 9492 427028 91532
rect 427532 80038 427588 394044
rect 434252 390628 434308 390638
rect 432684 388948 432740 388958
rect 432572 385588 432628 385598
rect 427980 369460 428036 369470
rect 427868 351988 427924 351998
rect 427756 343924 427812 343934
rect 427644 327796 427700 327806
rect 427644 107268 427700 327740
rect 427756 193284 427812 343868
rect 427868 236292 427924 351932
rect 427980 340340 428036 369404
rect 429436 367444 429492 367454
rect 427980 340274 428036 340284
rect 429212 352660 429268 352670
rect 427868 236226 427924 236236
rect 427980 317044 428036 317054
rect 427756 193218 427812 193228
rect 427644 107202 427700 107212
rect 427980 90748 428036 316988
rect 428540 299460 428596 299470
rect 428428 299236 428484 299246
rect 427980 90692 428148 90748
rect 427532 79972 427588 79982
rect 428092 75538 428148 90692
rect 428316 81284 428372 81294
rect 428092 75472 428148 75482
rect 428204 78148 428260 78158
rect 428204 13438 428260 78092
rect 428204 13372 428260 13382
rect 428316 12628 428372 81228
rect 428316 12562 428372 12572
rect 426972 9426 427028 9436
rect 426860 6178 426916 6188
rect 425068 6066 425124 6076
rect 424172 4834 424228 4844
rect 428428 4564 428484 299180
rect 428428 4498 428484 4508
rect 423836 4162 423892 4172
rect 428540 4228 428596 299404
rect 429212 239876 429268 352604
rect 429324 345380 429380 345390
rect 429324 243460 429380 345324
rect 429436 320180 429492 367388
rect 431228 357364 431284 357374
rect 429436 320114 429492 320124
rect 431004 335860 431060 335870
rect 429436 319060 429492 319070
rect 429436 303268 429492 319004
rect 429436 303202 429492 303212
rect 430892 315028 430948 315038
rect 429324 243394 429380 243404
rect 429212 239810 429268 239820
rect 429212 91028 429268 91038
rect 428652 75538 428708 75548
rect 428652 75460 428708 75482
rect 428652 75394 428708 75404
rect 429212 17668 429268 90972
rect 429660 88004 429716 88014
rect 429436 80612 429492 80622
rect 429436 29428 429492 80556
rect 429436 29362 429492 29372
rect 429212 17602 429268 17612
rect 429660 14308 429716 87948
rect 430892 49588 430948 314972
rect 431004 150276 431060 335804
rect 431116 323540 431172 323550
rect 431116 200452 431172 323484
rect 431228 264964 431284 357308
rect 431228 264898 431284 264908
rect 431788 299998 431844 300008
rect 431116 200386 431172 200396
rect 431004 150210 431060 150220
rect 430892 49522 430948 49532
rect 431228 89398 431284 89408
rect 431228 20020 431284 89342
rect 431228 19954 431284 19964
rect 429660 14242 429716 14252
rect 428540 4162 428596 4172
rect 431788 4228 431844 299942
rect 432460 91018 432516 91028
rect 432460 19908 432516 90962
rect 432572 89938 432628 385532
rect 432684 98578 432740 388892
rect 432908 372820 432964 372830
rect 432796 366772 432852 366782
rect 432796 334404 432852 366716
rect 432908 347396 432964 372764
rect 432908 347330 432964 347340
rect 433244 354676 433300 354686
rect 433132 346948 433188 346958
rect 433020 338548 433076 338558
rect 432796 334338 432852 334348
rect 432908 336532 432964 336542
rect 432684 98512 432740 98522
rect 432796 314356 432852 314366
rect 432572 89872 432628 89882
rect 432684 95844 432740 95854
rect 432684 20098 432740 95788
rect 432796 45332 432852 314300
rect 432908 153860 432964 336476
rect 433020 164612 433076 338492
rect 433132 214788 433188 346892
rect 433244 250628 433300 354620
rect 433244 250562 433300 250572
rect 433132 214722 433188 214732
rect 433020 164546 433076 164556
rect 432908 153794 432964 153804
rect 433132 91198 433188 91208
rect 433020 89218 433076 89228
rect 432796 45266 432852 45276
rect 432908 85978 432964 85988
rect 432684 20032 432740 20042
rect 432460 19842 432516 19852
rect 432908 14420 432964 85922
rect 433020 19796 433076 89162
rect 433020 19730 433076 19740
rect 433132 18116 433188 91142
rect 433356 90838 433412 90848
rect 433356 18340 433412 90782
rect 434252 80218 434308 390572
rect 435498 382350 436118 393242
rect 435498 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 436118 382350
rect 435498 382226 436118 382294
rect 435498 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 436118 382226
rect 435498 382102 436118 382170
rect 435498 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 436118 382102
rect 435498 381978 436118 382046
rect 435498 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 436118 381978
rect 434476 380660 434532 380670
rect 434252 80152 434308 80162
rect 434364 301258 434420 301268
rect 433356 18274 433412 18284
rect 433132 18050 433188 18060
rect 432908 14354 432964 14364
rect 434364 13300 434420 301202
rect 434476 80398 434532 380604
rect 435498 364350 436118 381922
rect 435498 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 436118 364350
rect 435498 364226 436118 364294
rect 435498 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 436118 364226
rect 435498 364102 436118 364170
rect 435498 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 436118 364102
rect 435498 363978 436118 364046
rect 435498 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 436118 363978
rect 434924 360052 434980 360062
rect 434812 342580 434868 342590
rect 434700 333172 434756 333182
rect 434588 331156 434644 331166
rect 434588 125188 434644 331100
rect 434700 135940 434756 333116
rect 434812 205044 434868 342524
rect 434924 279300 434980 359996
rect 434924 279234 434980 279244
rect 435498 346350 436118 363922
rect 435498 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 436118 346350
rect 435498 346226 436118 346294
rect 435498 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 436118 346226
rect 435498 346102 436118 346170
rect 435498 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 436118 346102
rect 435498 345978 436118 346046
rect 435498 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 436118 345978
rect 435498 328350 436118 345922
rect 435498 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 436118 328350
rect 435498 328226 436118 328294
rect 435498 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 436118 328226
rect 435498 328102 436118 328170
rect 435498 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 436118 328102
rect 435498 327978 436118 328046
rect 435498 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 436118 327978
rect 435498 310350 436118 327922
rect 435498 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 436118 310350
rect 435498 310226 436118 310294
rect 435498 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 436118 310226
rect 435498 310102 436118 310170
rect 435498 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 436118 310102
rect 435498 309978 436118 310046
rect 435498 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 436118 309978
rect 435498 292350 436118 309922
rect 435498 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 436118 292350
rect 435498 292226 436118 292294
rect 435498 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 436118 292226
rect 435498 292102 436118 292170
rect 435498 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 436118 292102
rect 435498 291978 436118 292046
rect 435498 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 436118 291978
rect 434812 204978 434868 204988
rect 435498 274350 436118 291922
rect 435498 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 436118 274350
rect 435498 274226 436118 274294
rect 435498 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 436118 274226
rect 435498 274102 436118 274170
rect 435498 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 436118 274102
rect 435498 273978 436118 274046
rect 435498 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 436118 273978
rect 435498 256350 436118 273922
rect 435498 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 436118 256350
rect 435498 256226 436118 256294
rect 435498 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 436118 256226
rect 435498 256102 436118 256170
rect 435498 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 436118 256102
rect 435498 255978 436118 256046
rect 435498 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 436118 255978
rect 435498 238350 436118 255922
rect 435498 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 436118 238350
rect 435498 238226 436118 238294
rect 435498 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 436118 238226
rect 435498 238102 436118 238170
rect 435498 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 436118 238102
rect 435498 237978 436118 238046
rect 435498 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 436118 237978
rect 435498 220350 436118 237922
rect 435498 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 436118 220350
rect 435498 220226 436118 220294
rect 435498 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 436118 220226
rect 435498 220102 436118 220170
rect 435498 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 436118 220102
rect 435498 219978 436118 220046
rect 435498 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 436118 219978
rect 434700 135874 434756 135884
rect 435498 202350 436118 219922
rect 435498 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 436118 202350
rect 435498 202226 436118 202294
rect 435498 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 436118 202226
rect 435498 202102 436118 202170
rect 435498 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 436118 202102
rect 435498 201978 436118 202046
rect 435498 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 436118 201978
rect 435498 184350 436118 201922
rect 435498 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 436118 184350
rect 435498 184226 436118 184294
rect 435498 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 436118 184226
rect 435498 184102 436118 184170
rect 435498 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 436118 184102
rect 435498 183978 436118 184046
rect 435498 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 436118 183978
rect 435498 166350 436118 183922
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 434588 125122 434644 125132
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 434476 80332 434532 80342
rect 435498 112350 436118 129922
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 435498 94350 436118 111922
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 434364 13234 434420 13244
rect 435498 76350 436118 93922
rect 436268 390740 436324 390750
rect 436268 93178 436324 390684
rect 437388 363412 437444 363422
rect 436604 355348 436660 355358
rect 436492 330484 436548 330494
rect 436268 93112 436324 93122
rect 436380 316372 436436 316382
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 435498 40350 436118 57922
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 431788 4162 431844 4172
rect 435498 4350 436118 21922
rect 436268 82918 436324 82928
rect 436268 7700 436324 82862
rect 436380 61348 436436 316316
rect 436492 121604 436548 330428
rect 436604 254212 436660 355292
rect 436604 254146 436660 254156
rect 436716 301812 436772 301822
rect 436716 204036 436772 301756
rect 436716 203970 436772 203980
rect 436828 299818 436884 299828
rect 436492 121538 436548 121548
rect 436380 61282 436436 61292
rect 436492 87598 436548 87608
rect 436492 16100 436548 87542
rect 436492 16034 436548 16044
rect 436604 84358 436660 84368
rect 436604 15958 436660 84302
rect 436604 15892 436660 15902
rect 436716 77698 436772 77708
rect 436716 12740 436772 77642
rect 436716 12674 436772 12684
rect 436268 7634 436324 7644
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 423388 1474 423444 1484
rect 435498 4102 436118 4170
rect 436828 4228 436884 299762
rect 437388 297220 437444 363356
rect 437388 297154 437444 297164
rect 437612 94978 437668 394156
rect 437724 390404 437780 390414
rect 437724 96778 437780 390348
rect 439218 388350 439838 393242
rect 439218 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 439838 388350
rect 439218 388226 439838 388294
rect 439218 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 439838 388226
rect 439218 388102 439838 388170
rect 439218 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 439838 388102
rect 439218 387978 439838 388046
rect 439218 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 439838 387978
rect 437948 373156 438004 373166
rect 437724 96712 437780 96722
rect 437836 300898 437892 300908
rect 437612 94912 437668 94922
rect 437836 17556 437892 300842
rect 437948 91558 438004 373100
rect 439218 370350 439838 387922
rect 439218 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 439838 370350
rect 439218 370226 439838 370294
rect 439218 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 439838 370226
rect 439218 370102 439838 370170
rect 439218 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 439838 370102
rect 439218 369978 439838 370046
rect 439218 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 439838 369978
rect 438396 362740 438452 362750
rect 438172 343588 438228 343598
rect 437948 91492 438004 91502
rect 438060 296660 438116 296670
rect 438060 71428 438116 296604
rect 438172 211204 438228 343532
rect 438284 335188 438340 335198
rect 438284 233492 438340 335132
rect 438396 293636 438452 362684
rect 439218 352350 439838 369922
rect 439218 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 439838 352350
rect 439218 352226 439838 352294
rect 439218 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 439838 352226
rect 439218 352102 439838 352170
rect 439218 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 439838 352102
rect 439218 351978 439838 352046
rect 439218 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 439838 351978
rect 438956 349972 439012 349982
rect 438396 293570 438452 293580
rect 438844 319732 438900 319742
rect 438844 248612 438900 319676
rect 438844 248546 438900 248556
rect 438284 233426 438340 233436
rect 438956 225540 439012 349916
rect 438956 225474 439012 225484
rect 439068 340228 439124 340238
rect 438172 211138 438228 211148
rect 439068 182532 439124 340172
rect 439068 182466 439124 182476
rect 439218 334350 439838 351922
rect 439218 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 439838 334350
rect 439218 334226 439838 334294
rect 439218 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 439838 334226
rect 439218 334102 439838 334170
rect 439218 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 439838 334102
rect 439218 333978 439838 334046
rect 439218 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 439838 333978
rect 439218 316350 439838 333922
rect 439218 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 439838 316350
rect 439218 316226 439838 316294
rect 439218 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 439838 316226
rect 439218 316102 439838 316170
rect 439218 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 439838 316102
rect 439218 315978 439838 316046
rect 439218 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 439838 315978
rect 439218 298350 439838 315922
rect 439218 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 439838 298350
rect 439218 298226 439838 298294
rect 439218 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 439838 298226
rect 439218 298102 439838 298170
rect 439218 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 439838 298102
rect 439218 297978 439838 298046
rect 439218 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 439838 297978
rect 439218 280350 439838 297922
rect 439218 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 439838 280350
rect 439218 280226 439838 280294
rect 439218 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 439838 280226
rect 439218 280102 439838 280170
rect 439218 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 439838 280102
rect 439218 279978 439838 280046
rect 439218 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 439838 279978
rect 439218 262350 439838 279922
rect 439218 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 439838 262350
rect 439218 262226 439838 262294
rect 439218 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 439838 262226
rect 439218 262102 439838 262170
rect 439218 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 439838 262102
rect 439218 261978 439838 262046
rect 439218 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 439838 261978
rect 439218 244350 439838 261922
rect 439218 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 439838 244350
rect 439218 244226 439838 244294
rect 439218 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 439838 244226
rect 439218 244102 439838 244170
rect 439218 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 439838 244102
rect 439218 243978 439838 244046
rect 439218 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 439838 243978
rect 439218 226350 439838 243922
rect 439218 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 439838 226350
rect 439218 226226 439838 226294
rect 439218 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 439838 226226
rect 439218 226102 439838 226170
rect 439218 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 439838 226102
rect 439218 225978 439838 226046
rect 439218 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 439838 225978
rect 439218 208350 439838 225922
rect 439218 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 439838 208350
rect 439218 208226 439838 208294
rect 439218 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 439838 208226
rect 439218 208102 439838 208170
rect 439218 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 439838 208102
rect 439218 207978 439838 208046
rect 439218 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 439838 207978
rect 439218 190350 439838 207922
rect 439218 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 439838 190350
rect 439218 190226 439838 190294
rect 439218 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 439838 190226
rect 439218 190102 439838 190170
rect 439218 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 439838 190102
rect 439218 189978 439838 190046
rect 439218 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 439838 189978
rect 439218 172350 439838 189922
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 439218 154350 439838 171922
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 439218 118350 439838 135922
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 439218 100350 439838 117922
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439068 82738 439124 82748
rect 438844 80938 438900 80948
rect 438060 71362 438116 71372
rect 438620 78058 438676 78068
rect 438620 20804 438676 78002
rect 438844 20916 438900 80882
rect 439068 21028 439124 82682
rect 439068 20962 439124 20972
rect 439218 82350 439838 99922
rect 439964 392338 440020 392348
rect 439964 98308 440020 392282
rect 440076 389060 440132 389070
rect 440076 98398 440132 389004
rect 441196 375396 441252 375406
rect 440972 368116 441028 368126
rect 440188 357028 440244 357038
rect 440188 354564 440244 356972
rect 440188 354498 440244 354508
rect 440188 348740 440244 348750
rect 440188 340228 440244 348684
rect 440188 340162 440244 340172
rect 440300 340340 440356 340350
rect 440300 337708 440356 340284
rect 440188 337652 440356 337708
rect 440188 329476 440244 337652
rect 440188 329410 440244 329420
rect 440748 331940 440804 331950
rect 440188 320180 440244 320190
rect 440188 318724 440244 320124
rect 440188 318658 440244 318668
rect 440748 300804 440804 331884
rect 440748 300738 440804 300748
rect 440860 330148 440916 330158
rect 440860 290052 440916 330092
rect 440972 322308 441028 368060
rect 441084 365540 441140 365550
rect 441084 325892 441140 365484
rect 441196 361732 441252 375340
rect 441196 361666 441252 361676
rect 441196 360388 441252 360398
rect 441196 336644 441252 360332
rect 442540 358708 442596 358718
rect 441308 353668 441364 353678
rect 441308 343812 441364 353612
rect 441308 343746 441364 343756
rect 441644 341908 441700 341918
rect 441196 336578 441252 336588
rect 441532 336868 441588 336878
rect 441084 325826 441140 325836
rect 441308 334404 441364 334414
rect 440972 322242 441028 322252
rect 441196 323428 441252 323438
rect 441084 320068 441140 320078
rect 440860 289986 440916 289996
rect 440972 303268 441028 303278
rect 440188 120148 440244 120158
rect 440188 118020 440244 120092
rect 440188 117954 440244 117964
rect 440188 105028 440244 105038
rect 440188 100100 440244 104972
rect 440188 100034 440244 100044
rect 440076 98332 440132 98342
rect 439964 98242 440020 98252
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 440076 87418 440132 87428
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 439218 46350 439838 63922
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 439218 28350 439838 45922
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 438844 20850 438900 20860
rect 438620 20738 438676 20748
rect 437836 17490 437892 17500
rect 436828 4162 436884 4172
rect 439218 10350 439838 27922
rect 439964 77338 440020 77348
rect 439964 15988 440020 77282
rect 440076 17668 440132 87362
rect 440412 81508 440468 81518
rect 440188 78372 440244 78382
rect 440188 67844 440244 78316
rect 440412 75012 440468 81452
rect 440412 74946 440468 74956
rect 440188 67778 440244 67788
rect 440972 60676 441028 303212
rect 441084 85764 441140 320012
rect 441196 261380 441252 323372
rect 441308 315140 441364 334348
rect 441308 315074 441364 315084
rect 441420 301700 441476 301710
rect 441196 261314 441252 261324
rect 441308 294868 441364 294878
rect 441084 85698 441140 85708
rect 441196 248612 441252 248622
rect 440972 60610 441028 60620
rect 441084 75460 441140 75470
rect 440972 49588 441028 49598
rect 440188 45332 440244 45342
rect 440188 39172 440244 45276
rect 440972 42756 441028 49532
rect 440972 42690 441028 42700
rect 440188 39106 440244 39116
rect 441084 35588 441140 75404
rect 441196 64260 441252 248556
rect 441308 114436 441364 294812
rect 441420 171780 441476 301644
rect 441532 232708 441588 336812
rect 441644 333060 441700 341852
rect 441644 332994 441700 333004
rect 441532 232642 441588 232652
rect 441644 313348 441700 313358
rect 441644 218372 441700 313292
rect 441756 301588 441812 301598
rect 441756 247044 441812 301532
rect 442540 272132 442596 358652
rect 442540 272066 442596 272076
rect 441756 246978 441812 246988
rect 441644 218306 441700 218316
rect 441756 233492 441812 233502
rect 441532 205044 441588 205054
rect 441532 186116 441588 204988
rect 441532 186050 441588 186060
rect 441420 171714 441476 171724
rect 441532 173908 441588 173918
rect 441308 114370 441364 114380
rect 441420 170548 441476 170558
rect 441196 64194 441252 64204
rect 441308 83300 441364 83310
rect 441196 61348 441252 61358
rect 441196 49924 441252 61292
rect 441196 49858 441252 49868
rect 441308 46340 441364 83244
rect 441420 78596 441476 170492
rect 441532 157444 441588 173852
rect 441532 157378 441588 157388
rect 441756 146692 441812 233436
rect 441756 146626 441812 146636
rect 441644 86548 441700 86558
rect 441420 78530 441476 78540
rect 441532 85092 441588 85102
rect 441532 53508 441588 85036
rect 441644 57092 441700 86492
rect 442652 80578 442708 394268
rect 443436 392980 443492 392990
rect 442876 392868 442932 392878
rect 442652 80512 442708 80522
rect 442764 300178 442820 300188
rect 441644 57026 441700 57036
rect 442652 67978 442708 67988
rect 441532 53442 441588 53452
rect 441308 46274 441364 46284
rect 441084 35522 441140 35532
rect 440076 17602 440132 17612
rect 442652 16772 442708 67922
rect 442652 16706 442708 16716
rect 439964 15922 440020 15932
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 -1120 439838 9922
rect 442764 4900 442820 300122
rect 442876 96598 442932 392812
rect 443212 392756 443268 392766
rect 443100 392518 443156 392528
rect 442876 96532 442932 96542
rect 442988 299012 443044 299022
rect 442876 84178 442932 84188
rect 442876 12628 442932 84122
rect 442876 12562 442932 12572
rect 442764 4834 442820 4844
rect 442988 4788 443044 298956
rect 443100 98218 443156 392462
rect 443212 101818 443268 392700
rect 443324 348628 443380 348638
rect 443324 229124 443380 348572
rect 443324 229058 443380 229068
rect 443212 101752 443268 101762
rect 443436 101638 443492 392924
rect 547708 386148 547764 590716
rect 547708 386082 547764 386092
rect 547820 575652 547876 575662
rect 547820 372260 547876 575596
rect 547932 575428 547988 575438
rect 547932 374612 547988 575372
rect 548044 392518 548100 590940
rect 548156 590884 548212 590894
rect 548156 392868 548212 590828
rect 548268 590548 548324 590558
rect 548268 392980 548324 590492
rect 548268 392914 548324 392924
rect 548156 392802 548212 392812
rect 548044 392452 548100 392462
rect 549388 389396 549444 591052
rect 549612 590660 549668 590670
rect 549388 389330 549444 389340
rect 549500 575540 549556 575550
rect 547932 374546 547988 374556
rect 549500 373940 549556 575484
rect 549612 392756 549668 590604
rect 549612 392690 549668 392700
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 558378 544350 558998 561922
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 558378 472350 558998 489922
rect 558378 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 558998 472350
rect 558378 472226 558998 472294
rect 558378 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 558998 472226
rect 558378 472102 558998 472170
rect 558378 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 558998 472102
rect 558378 471978 558998 472046
rect 558378 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 558998 471978
rect 558378 454350 558998 471922
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 549500 373874 549556 373884
rect 558378 382350 558998 399922
rect 558378 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 558998 382350
rect 558378 382226 558998 382294
rect 558378 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 558998 382226
rect 558378 382102 558998 382170
rect 558378 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 558998 382102
rect 558378 381978 558998 382046
rect 558378 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 558998 381978
rect 547820 372194 547876 372204
rect 558378 372094 558998 381922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 562098 550350 562718 567922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 562098 532350 562718 549922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 562098 478350 562718 495922
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 562098 460350 562718 477922
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 388350 562718 405922
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 562098 372094 562718 387922
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 589098 580350 589718 596784
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 589098 562350 589718 579922
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 589098 382350 589718 399922
rect 590492 588644 590548 588654
rect 590492 390628 590548 588588
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 590604 562212 590660 562222
rect 590604 394100 590660 562156
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 590604 394034 590660 394044
rect 590716 548996 590772 549006
rect 590492 390562 590548 390572
rect 590716 389060 590772 548940
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 590828 509348 590884 509358
rect 590828 392338 590884 509292
rect 590828 392272 590884 392282
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 590716 388994 590772 389004
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 463808 370350 464128 370384
rect 463808 370294 463878 370350
rect 463934 370294 464002 370350
rect 464058 370294 464128 370350
rect 463808 370226 464128 370294
rect 463808 370170 463878 370226
rect 463934 370170 464002 370226
rect 464058 370170 464128 370226
rect 463808 370102 464128 370170
rect 463808 370046 463878 370102
rect 463934 370046 464002 370102
rect 464058 370046 464128 370102
rect 463808 369978 464128 370046
rect 463808 369922 463878 369978
rect 463934 369922 464002 369978
rect 464058 369922 464128 369978
rect 463808 369888 464128 369922
rect 494528 370350 494848 370384
rect 494528 370294 494598 370350
rect 494654 370294 494722 370350
rect 494778 370294 494848 370350
rect 494528 370226 494848 370294
rect 494528 370170 494598 370226
rect 494654 370170 494722 370226
rect 494778 370170 494848 370226
rect 494528 370102 494848 370170
rect 494528 370046 494598 370102
rect 494654 370046 494722 370102
rect 494778 370046 494848 370102
rect 494528 369978 494848 370046
rect 494528 369922 494598 369978
rect 494654 369922 494722 369978
rect 494778 369922 494848 369978
rect 494528 369888 494848 369922
rect 525248 370350 525568 370384
rect 525248 370294 525318 370350
rect 525374 370294 525442 370350
rect 525498 370294 525568 370350
rect 525248 370226 525568 370294
rect 525248 370170 525318 370226
rect 525374 370170 525442 370226
rect 525498 370170 525568 370226
rect 525248 370102 525568 370170
rect 525248 370046 525318 370102
rect 525374 370046 525442 370102
rect 525498 370046 525568 370102
rect 525248 369978 525568 370046
rect 525248 369922 525318 369978
rect 525374 369922 525442 369978
rect 525498 369922 525568 369978
rect 525248 369888 525568 369922
rect 555968 370350 556288 370384
rect 555968 370294 556038 370350
rect 556094 370294 556162 370350
rect 556218 370294 556288 370350
rect 555968 370226 556288 370294
rect 555968 370170 556038 370226
rect 556094 370170 556162 370226
rect 556218 370170 556288 370226
rect 555968 370102 556288 370170
rect 555968 370046 556038 370102
rect 556094 370046 556162 370102
rect 556218 370046 556288 370102
rect 555968 369978 556288 370046
rect 555968 369922 556038 369978
rect 556094 369922 556162 369978
rect 556218 369922 556288 369978
rect 555968 369888 556288 369922
rect 448448 364350 448768 364384
rect 448448 364294 448518 364350
rect 448574 364294 448642 364350
rect 448698 364294 448768 364350
rect 448448 364226 448768 364294
rect 448448 364170 448518 364226
rect 448574 364170 448642 364226
rect 448698 364170 448768 364226
rect 448448 364102 448768 364170
rect 448448 364046 448518 364102
rect 448574 364046 448642 364102
rect 448698 364046 448768 364102
rect 448448 363978 448768 364046
rect 448448 363922 448518 363978
rect 448574 363922 448642 363978
rect 448698 363922 448768 363978
rect 448448 363888 448768 363922
rect 479168 364350 479488 364384
rect 479168 364294 479238 364350
rect 479294 364294 479362 364350
rect 479418 364294 479488 364350
rect 479168 364226 479488 364294
rect 479168 364170 479238 364226
rect 479294 364170 479362 364226
rect 479418 364170 479488 364226
rect 479168 364102 479488 364170
rect 479168 364046 479238 364102
rect 479294 364046 479362 364102
rect 479418 364046 479488 364102
rect 479168 363978 479488 364046
rect 479168 363922 479238 363978
rect 479294 363922 479362 363978
rect 479418 363922 479488 363978
rect 479168 363888 479488 363922
rect 509888 364350 510208 364384
rect 509888 364294 509958 364350
rect 510014 364294 510082 364350
rect 510138 364294 510208 364350
rect 509888 364226 510208 364294
rect 509888 364170 509958 364226
rect 510014 364170 510082 364226
rect 510138 364170 510208 364226
rect 509888 364102 510208 364170
rect 509888 364046 509958 364102
rect 510014 364046 510082 364102
rect 510138 364046 510208 364102
rect 509888 363978 510208 364046
rect 509888 363922 509958 363978
rect 510014 363922 510082 363978
rect 510138 363922 510208 363978
rect 509888 363888 510208 363922
rect 540608 364350 540928 364384
rect 540608 364294 540678 364350
rect 540734 364294 540802 364350
rect 540858 364294 540928 364350
rect 540608 364226 540928 364294
rect 540608 364170 540678 364226
rect 540734 364170 540802 364226
rect 540858 364170 540928 364226
rect 540608 364102 540928 364170
rect 540608 364046 540678 364102
rect 540734 364046 540802 364102
rect 540858 364046 540928 364102
rect 540608 363978 540928 364046
rect 540608 363922 540678 363978
rect 540734 363922 540802 363978
rect 540858 363922 540928 363978
rect 540608 363888 540928 363922
rect 571328 364350 571648 364384
rect 571328 364294 571398 364350
rect 571454 364294 571522 364350
rect 571578 364294 571648 364350
rect 571328 364226 571648 364294
rect 571328 364170 571398 364226
rect 571454 364170 571522 364226
rect 571578 364170 571648 364226
rect 571328 364102 571648 364170
rect 571328 364046 571398 364102
rect 571454 364046 571522 364102
rect 571578 364046 571648 364102
rect 571328 363978 571648 364046
rect 571328 363922 571398 363978
rect 571454 363922 571522 363978
rect 571578 363922 571648 363978
rect 571328 363888 571648 363922
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 463808 352350 464128 352384
rect 463808 352294 463878 352350
rect 463934 352294 464002 352350
rect 464058 352294 464128 352350
rect 463808 352226 464128 352294
rect 463808 352170 463878 352226
rect 463934 352170 464002 352226
rect 464058 352170 464128 352226
rect 463808 352102 464128 352170
rect 463808 352046 463878 352102
rect 463934 352046 464002 352102
rect 464058 352046 464128 352102
rect 463808 351978 464128 352046
rect 463808 351922 463878 351978
rect 463934 351922 464002 351978
rect 464058 351922 464128 351978
rect 463808 351888 464128 351922
rect 494528 352350 494848 352384
rect 494528 352294 494598 352350
rect 494654 352294 494722 352350
rect 494778 352294 494848 352350
rect 494528 352226 494848 352294
rect 494528 352170 494598 352226
rect 494654 352170 494722 352226
rect 494778 352170 494848 352226
rect 494528 352102 494848 352170
rect 494528 352046 494598 352102
rect 494654 352046 494722 352102
rect 494778 352046 494848 352102
rect 494528 351978 494848 352046
rect 494528 351922 494598 351978
rect 494654 351922 494722 351978
rect 494778 351922 494848 351978
rect 494528 351888 494848 351922
rect 525248 352350 525568 352384
rect 525248 352294 525318 352350
rect 525374 352294 525442 352350
rect 525498 352294 525568 352350
rect 525248 352226 525568 352294
rect 525248 352170 525318 352226
rect 525374 352170 525442 352226
rect 525498 352170 525568 352226
rect 525248 352102 525568 352170
rect 525248 352046 525318 352102
rect 525374 352046 525442 352102
rect 525498 352046 525568 352102
rect 525248 351978 525568 352046
rect 525248 351922 525318 351978
rect 525374 351922 525442 351978
rect 525498 351922 525568 351978
rect 525248 351888 525568 351922
rect 555968 352350 556288 352384
rect 555968 352294 556038 352350
rect 556094 352294 556162 352350
rect 556218 352294 556288 352350
rect 555968 352226 556288 352294
rect 555968 352170 556038 352226
rect 556094 352170 556162 352226
rect 556218 352170 556288 352226
rect 555968 352102 556288 352170
rect 555968 352046 556038 352102
rect 556094 352046 556162 352102
rect 556218 352046 556288 352102
rect 555968 351978 556288 352046
rect 555968 351922 556038 351978
rect 556094 351922 556162 351978
rect 556218 351922 556288 351978
rect 555968 351888 556288 351922
rect 448448 346350 448768 346384
rect 448448 346294 448518 346350
rect 448574 346294 448642 346350
rect 448698 346294 448768 346350
rect 448448 346226 448768 346294
rect 448448 346170 448518 346226
rect 448574 346170 448642 346226
rect 448698 346170 448768 346226
rect 448448 346102 448768 346170
rect 448448 346046 448518 346102
rect 448574 346046 448642 346102
rect 448698 346046 448768 346102
rect 448448 345978 448768 346046
rect 448448 345922 448518 345978
rect 448574 345922 448642 345978
rect 448698 345922 448768 345978
rect 448448 345888 448768 345922
rect 479168 346350 479488 346384
rect 479168 346294 479238 346350
rect 479294 346294 479362 346350
rect 479418 346294 479488 346350
rect 479168 346226 479488 346294
rect 479168 346170 479238 346226
rect 479294 346170 479362 346226
rect 479418 346170 479488 346226
rect 479168 346102 479488 346170
rect 479168 346046 479238 346102
rect 479294 346046 479362 346102
rect 479418 346046 479488 346102
rect 479168 345978 479488 346046
rect 479168 345922 479238 345978
rect 479294 345922 479362 345978
rect 479418 345922 479488 345978
rect 479168 345888 479488 345922
rect 509888 346350 510208 346384
rect 509888 346294 509958 346350
rect 510014 346294 510082 346350
rect 510138 346294 510208 346350
rect 509888 346226 510208 346294
rect 509888 346170 509958 346226
rect 510014 346170 510082 346226
rect 510138 346170 510208 346226
rect 509888 346102 510208 346170
rect 509888 346046 509958 346102
rect 510014 346046 510082 346102
rect 510138 346046 510208 346102
rect 509888 345978 510208 346046
rect 509888 345922 509958 345978
rect 510014 345922 510082 345978
rect 510138 345922 510208 345978
rect 509888 345888 510208 345922
rect 540608 346350 540928 346384
rect 540608 346294 540678 346350
rect 540734 346294 540802 346350
rect 540858 346294 540928 346350
rect 540608 346226 540928 346294
rect 540608 346170 540678 346226
rect 540734 346170 540802 346226
rect 540858 346170 540928 346226
rect 540608 346102 540928 346170
rect 540608 346046 540678 346102
rect 540734 346046 540802 346102
rect 540858 346046 540928 346102
rect 540608 345978 540928 346046
rect 540608 345922 540678 345978
rect 540734 345922 540802 345978
rect 540858 345922 540928 345978
rect 540608 345888 540928 345922
rect 571328 346350 571648 346384
rect 571328 346294 571398 346350
rect 571454 346294 571522 346350
rect 571578 346294 571648 346350
rect 571328 346226 571648 346294
rect 571328 346170 571398 346226
rect 571454 346170 571522 346226
rect 571578 346170 571648 346226
rect 571328 346102 571648 346170
rect 571328 346046 571398 346102
rect 571454 346046 571522 346102
rect 571578 346046 571648 346102
rect 571328 345978 571648 346046
rect 571328 345922 571398 345978
rect 571454 345922 571522 345978
rect 571578 345922 571648 345978
rect 571328 345888 571648 345922
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 463808 334350 464128 334384
rect 463808 334294 463878 334350
rect 463934 334294 464002 334350
rect 464058 334294 464128 334350
rect 463808 334226 464128 334294
rect 463808 334170 463878 334226
rect 463934 334170 464002 334226
rect 464058 334170 464128 334226
rect 463808 334102 464128 334170
rect 463808 334046 463878 334102
rect 463934 334046 464002 334102
rect 464058 334046 464128 334102
rect 463808 333978 464128 334046
rect 463808 333922 463878 333978
rect 463934 333922 464002 333978
rect 464058 333922 464128 333978
rect 463808 333888 464128 333922
rect 494528 334350 494848 334384
rect 494528 334294 494598 334350
rect 494654 334294 494722 334350
rect 494778 334294 494848 334350
rect 494528 334226 494848 334294
rect 494528 334170 494598 334226
rect 494654 334170 494722 334226
rect 494778 334170 494848 334226
rect 494528 334102 494848 334170
rect 494528 334046 494598 334102
rect 494654 334046 494722 334102
rect 494778 334046 494848 334102
rect 494528 333978 494848 334046
rect 494528 333922 494598 333978
rect 494654 333922 494722 333978
rect 494778 333922 494848 333978
rect 494528 333888 494848 333922
rect 525248 334350 525568 334384
rect 525248 334294 525318 334350
rect 525374 334294 525442 334350
rect 525498 334294 525568 334350
rect 525248 334226 525568 334294
rect 525248 334170 525318 334226
rect 525374 334170 525442 334226
rect 525498 334170 525568 334226
rect 525248 334102 525568 334170
rect 525248 334046 525318 334102
rect 525374 334046 525442 334102
rect 525498 334046 525568 334102
rect 525248 333978 525568 334046
rect 525248 333922 525318 333978
rect 525374 333922 525442 333978
rect 525498 333922 525568 333978
rect 525248 333888 525568 333922
rect 555968 334350 556288 334384
rect 555968 334294 556038 334350
rect 556094 334294 556162 334350
rect 556218 334294 556288 334350
rect 555968 334226 556288 334294
rect 555968 334170 556038 334226
rect 556094 334170 556162 334226
rect 556218 334170 556288 334226
rect 555968 334102 556288 334170
rect 555968 334046 556038 334102
rect 556094 334046 556162 334102
rect 556218 334046 556288 334102
rect 555968 333978 556288 334046
rect 555968 333922 556038 333978
rect 556094 333922 556162 333978
rect 556218 333922 556288 333978
rect 555968 333888 556288 333922
rect 448448 328350 448768 328384
rect 448448 328294 448518 328350
rect 448574 328294 448642 328350
rect 448698 328294 448768 328350
rect 448448 328226 448768 328294
rect 448448 328170 448518 328226
rect 448574 328170 448642 328226
rect 448698 328170 448768 328226
rect 448448 328102 448768 328170
rect 448448 328046 448518 328102
rect 448574 328046 448642 328102
rect 448698 328046 448768 328102
rect 448448 327978 448768 328046
rect 448448 327922 448518 327978
rect 448574 327922 448642 327978
rect 448698 327922 448768 327978
rect 448448 327888 448768 327922
rect 479168 328350 479488 328384
rect 479168 328294 479238 328350
rect 479294 328294 479362 328350
rect 479418 328294 479488 328350
rect 479168 328226 479488 328294
rect 479168 328170 479238 328226
rect 479294 328170 479362 328226
rect 479418 328170 479488 328226
rect 479168 328102 479488 328170
rect 479168 328046 479238 328102
rect 479294 328046 479362 328102
rect 479418 328046 479488 328102
rect 479168 327978 479488 328046
rect 479168 327922 479238 327978
rect 479294 327922 479362 327978
rect 479418 327922 479488 327978
rect 479168 327888 479488 327922
rect 509888 328350 510208 328384
rect 509888 328294 509958 328350
rect 510014 328294 510082 328350
rect 510138 328294 510208 328350
rect 509888 328226 510208 328294
rect 509888 328170 509958 328226
rect 510014 328170 510082 328226
rect 510138 328170 510208 328226
rect 509888 328102 510208 328170
rect 509888 328046 509958 328102
rect 510014 328046 510082 328102
rect 510138 328046 510208 328102
rect 509888 327978 510208 328046
rect 509888 327922 509958 327978
rect 510014 327922 510082 327978
rect 510138 327922 510208 327978
rect 509888 327888 510208 327922
rect 540608 328350 540928 328384
rect 540608 328294 540678 328350
rect 540734 328294 540802 328350
rect 540858 328294 540928 328350
rect 540608 328226 540928 328294
rect 540608 328170 540678 328226
rect 540734 328170 540802 328226
rect 540858 328170 540928 328226
rect 540608 328102 540928 328170
rect 540608 328046 540678 328102
rect 540734 328046 540802 328102
rect 540858 328046 540928 328102
rect 540608 327978 540928 328046
rect 540608 327922 540678 327978
rect 540734 327922 540802 327978
rect 540858 327922 540928 327978
rect 540608 327888 540928 327922
rect 571328 328350 571648 328384
rect 571328 328294 571398 328350
rect 571454 328294 571522 328350
rect 571578 328294 571648 328350
rect 571328 328226 571648 328294
rect 571328 328170 571398 328226
rect 571454 328170 571522 328226
rect 571578 328170 571648 328226
rect 571328 328102 571648 328170
rect 571328 328046 571398 328102
rect 571454 328046 571522 328102
rect 571578 328046 571648 328102
rect 571328 327978 571648 328046
rect 571328 327922 571398 327978
rect 571454 327922 571522 327978
rect 571578 327922 571648 327978
rect 571328 327888 571648 327922
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 463808 316350 464128 316384
rect 463808 316294 463878 316350
rect 463934 316294 464002 316350
rect 464058 316294 464128 316350
rect 463808 316226 464128 316294
rect 463808 316170 463878 316226
rect 463934 316170 464002 316226
rect 464058 316170 464128 316226
rect 463808 316102 464128 316170
rect 463808 316046 463878 316102
rect 463934 316046 464002 316102
rect 464058 316046 464128 316102
rect 463808 315978 464128 316046
rect 463808 315922 463878 315978
rect 463934 315922 464002 315978
rect 464058 315922 464128 315978
rect 463808 315888 464128 315922
rect 494528 316350 494848 316384
rect 494528 316294 494598 316350
rect 494654 316294 494722 316350
rect 494778 316294 494848 316350
rect 494528 316226 494848 316294
rect 494528 316170 494598 316226
rect 494654 316170 494722 316226
rect 494778 316170 494848 316226
rect 494528 316102 494848 316170
rect 494528 316046 494598 316102
rect 494654 316046 494722 316102
rect 494778 316046 494848 316102
rect 494528 315978 494848 316046
rect 494528 315922 494598 315978
rect 494654 315922 494722 315978
rect 494778 315922 494848 315978
rect 494528 315888 494848 315922
rect 525248 316350 525568 316384
rect 525248 316294 525318 316350
rect 525374 316294 525442 316350
rect 525498 316294 525568 316350
rect 525248 316226 525568 316294
rect 525248 316170 525318 316226
rect 525374 316170 525442 316226
rect 525498 316170 525568 316226
rect 525248 316102 525568 316170
rect 525248 316046 525318 316102
rect 525374 316046 525442 316102
rect 525498 316046 525568 316102
rect 525248 315978 525568 316046
rect 525248 315922 525318 315978
rect 525374 315922 525442 315978
rect 525498 315922 525568 315978
rect 525248 315888 525568 315922
rect 555968 316350 556288 316384
rect 555968 316294 556038 316350
rect 556094 316294 556162 316350
rect 556218 316294 556288 316350
rect 555968 316226 556288 316294
rect 555968 316170 556038 316226
rect 556094 316170 556162 316226
rect 556218 316170 556288 316226
rect 555968 316102 556288 316170
rect 555968 316046 556038 316102
rect 556094 316046 556162 316102
rect 556218 316046 556288 316102
rect 555968 315978 556288 316046
rect 555968 315922 556038 315978
rect 556094 315922 556162 315978
rect 556218 315922 556288 315978
rect 555968 315888 556288 315922
rect 448448 310350 448768 310384
rect 448448 310294 448518 310350
rect 448574 310294 448642 310350
rect 448698 310294 448768 310350
rect 448448 310226 448768 310294
rect 448448 310170 448518 310226
rect 448574 310170 448642 310226
rect 448698 310170 448768 310226
rect 448448 310102 448768 310170
rect 448448 310046 448518 310102
rect 448574 310046 448642 310102
rect 448698 310046 448768 310102
rect 448448 309978 448768 310046
rect 448448 309922 448518 309978
rect 448574 309922 448642 309978
rect 448698 309922 448768 309978
rect 448448 309888 448768 309922
rect 479168 310350 479488 310384
rect 479168 310294 479238 310350
rect 479294 310294 479362 310350
rect 479418 310294 479488 310350
rect 479168 310226 479488 310294
rect 479168 310170 479238 310226
rect 479294 310170 479362 310226
rect 479418 310170 479488 310226
rect 479168 310102 479488 310170
rect 479168 310046 479238 310102
rect 479294 310046 479362 310102
rect 479418 310046 479488 310102
rect 479168 309978 479488 310046
rect 479168 309922 479238 309978
rect 479294 309922 479362 309978
rect 479418 309922 479488 309978
rect 479168 309888 479488 309922
rect 509888 310350 510208 310384
rect 509888 310294 509958 310350
rect 510014 310294 510082 310350
rect 510138 310294 510208 310350
rect 509888 310226 510208 310294
rect 509888 310170 509958 310226
rect 510014 310170 510082 310226
rect 510138 310170 510208 310226
rect 509888 310102 510208 310170
rect 509888 310046 509958 310102
rect 510014 310046 510082 310102
rect 510138 310046 510208 310102
rect 509888 309978 510208 310046
rect 509888 309922 509958 309978
rect 510014 309922 510082 309978
rect 510138 309922 510208 309978
rect 509888 309888 510208 309922
rect 540608 310350 540928 310384
rect 540608 310294 540678 310350
rect 540734 310294 540802 310350
rect 540858 310294 540928 310350
rect 540608 310226 540928 310294
rect 540608 310170 540678 310226
rect 540734 310170 540802 310226
rect 540858 310170 540928 310226
rect 540608 310102 540928 310170
rect 540608 310046 540678 310102
rect 540734 310046 540802 310102
rect 540858 310046 540928 310102
rect 540608 309978 540928 310046
rect 540608 309922 540678 309978
rect 540734 309922 540802 309978
rect 540858 309922 540928 309978
rect 540608 309888 540928 309922
rect 571328 310350 571648 310384
rect 571328 310294 571398 310350
rect 571454 310294 571522 310350
rect 571578 310294 571648 310350
rect 571328 310226 571648 310294
rect 571328 310170 571398 310226
rect 571454 310170 571522 310226
rect 571578 310170 571648 310226
rect 571328 310102 571648 310170
rect 571328 310046 571398 310102
rect 571454 310046 571522 310102
rect 571578 310046 571648 310102
rect 571328 309978 571648 310046
rect 571328 309922 571398 309978
rect 571454 309922 571522 309978
rect 571578 309922 571648 309978
rect 571328 309888 571648 309922
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 463808 298350 464128 298384
rect 463808 298294 463878 298350
rect 463934 298294 464002 298350
rect 464058 298294 464128 298350
rect 463808 298226 464128 298294
rect 463808 298170 463878 298226
rect 463934 298170 464002 298226
rect 464058 298170 464128 298226
rect 463808 298102 464128 298170
rect 463808 298046 463878 298102
rect 463934 298046 464002 298102
rect 464058 298046 464128 298102
rect 463808 297978 464128 298046
rect 463808 297922 463878 297978
rect 463934 297922 464002 297978
rect 464058 297922 464128 297978
rect 463808 297888 464128 297922
rect 494528 298350 494848 298384
rect 494528 298294 494598 298350
rect 494654 298294 494722 298350
rect 494778 298294 494848 298350
rect 494528 298226 494848 298294
rect 494528 298170 494598 298226
rect 494654 298170 494722 298226
rect 494778 298170 494848 298226
rect 494528 298102 494848 298170
rect 494528 298046 494598 298102
rect 494654 298046 494722 298102
rect 494778 298046 494848 298102
rect 494528 297978 494848 298046
rect 494528 297922 494598 297978
rect 494654 297922 494722 297978
rect 494778 297922 494848 297978
rect 494528 297888 494848 297922
rect 525248 298350 525568 298384
rect 525248 298294 525318 298350
rect 525374 298294 525442 298350
rect 525498 298294 525568 298350
rect 525248 298226 525568 298294
rect 525248 298170 525318 298226
rect 525374 298170 525442 298226
rect 525498 298170 525568 298226
rect 525248 298102 525568 298170
rect 525248 298046 525318 298102
rect 525374 298046 525442 298102
rect 525498 298046 525568 298102
rect 525248 297978 525568 298046
rect 525248 297922 525318 297978
rect 525374 297922 525442 297978
rect 525498 297922 525568 297978
rect 525248 297888 525568 297922
rect 555968 298350 556288 298384
rect 555968 298294 556038 298350
rect 556094 298294 556162 298350
rect 556218 298294 556288 298350
rect 555968 298226 556288 298294
rect 555968 298170 556038 298226
rect 556094 298170 556162 298226
rect 556218 298170 556288 298226
rect 555968 298102 556288 298170
rect 555968 298046 556038 298102
rect 556094 298046 556162 298102
rect 556218 298046 556288 298102
rect 555968 297978 556288 298046
rect 555968 297922 556038 297978
rect 556094 297922 556162 297978
rect 556218 297922 556288 297978
rect 555968 297888 556288 297922
rect 448448 292350 448768 292384
rect 448448 292294 448518 292350
rect 448574 292294 448642 292350
rect 448698 292294 448768 292350
rect 448448 292226 448768 292294
rect 448448 292170 448518 292226
rect 448574 292170 448642 292226
rect 448698 292170 448768 292226
rect 448448 292102 448768 292170
rect 448448 292046 448518 292102
rect 448574 292046 448642 292102
rect 448698 292046 448768 292102
rect 448448 291978 448768 292046
rect 448448 291922 448518 291978
rect 448574 291922 448642 291978
rect 448698 291922 448768 291978
rect 448448 291888 448768 291922
rect 479168 292350 479488 292384
rect 479168 292294 479238 292350
rect 479294 292294 479362 292350
rect 479418 292294 479488 292350
rect 479168 292226 479488 292294
rect 479168 292170 479238 292226
rect 479294 292170 479362 292226
rect 479418 292170 479488 292226
rect 479168 292102 479488 292170
rect 479168 292046 479238 292102
rect 479294 292046 479362 292102
rect 479418 292046 479488 292102
rect 479168 291978 479488 292046
rect 479168 291922 479238 291978
rect 479294 291922 479362 291978
rect 479418 291922 479488 291978
rect 479168 291888 479488 291922
rect 509888 292350 510208 292384
rect 509888 292294 509958 292350
rect 510014 292294 510082 292350
rect 510138 292294 510208 292350
rect 509888 292226 510208 292294
rect 509888 292170 509958 292226
rect 510014 292170 510082 292226
rect 510138 292170 510208 292226
rect 509888 292102 510208 292170
rect 509888 292046 509958 292102
rect 510014 292046 510082 292102
rect 510138 292046 510208 292102
rect 509888 291978 510208 292046
rect 509888 291922 509958 291978
rect 510014 291922 510082 291978
rect 510138 291922 510208 291978
rect 509888 291888 510208 291922
rect 540608 292350 540928 292384
rect 540608 292294 540678 292350
rect 540734 292294 540802 292350
rect 540858 292294 540928 292350
rect 540608 292226 540928 292294
rect 540608 292170 540678 292226
rect 540734 292170 540802 292226
rect 540858 292170 540928 292226
rect 540608 292102 540928 292170
rect 540608 292046 540678 292102
rect 540734 292046 540802 292102
rect 540858 292046 540928 292102
rect 540608 291978 540928 292046
rect 540608 291922 540678 291978
rect 540734 291922 540802 291978
rect 540858 291922 540928 291978
rect 540608 291888 540928 291922
rect 571328 292350 571648 292384
rect 571328 292294 571398 292350
rect 571454 292294 571522 292350
rect 571578 292294 571648 292350
rect 571328 292226 571648 292294
rect 571328 292170 571398 292226
rect 571454 292170 571522 292226
rect 571578 292170 571648 292226
rect 571328 292102 571648 292170
rect 571328 292046 571398 292102
rect 571454 292046 571522 292102
rect 571578 292046 571648 292102
rect 571328 291978 571648 292046
rect 571328 291922 571398 291978
rect 571454 291922 571522 291978
rect 571578 291922 571648 291978
rect 571328 291888 571648 291922
rect 589098 292350 589718 309922
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 463808 280350 464128 280384
rect 463808 280294 463878 280350
rect 463934 280294 464002 280350
rect 464058 280294 464128 280350
rect 463808 280226 464128 280294
rect 463808 280170 463878 280226
rect 463934 280170 464002 280226
rect 464058 280170 464128 280226
rect 463808 280102 464128 280170
rect 463808 280046 463878 280102
rect 463934 280046 464002 280102
rect 464058 280046 464128 280102
rect 463808 279978 464128 280046
rect 463808 279922 463878 279978
rect 463934 279922 464002 279978
rect 464058 279922 464128 279978
rect 463808 279888 464128 279922
rect 494528 280350 494848 280384
rect 494528 280294 494598 280350
rect 494654 280294 494722 280350
rect 494778 280294 494848 280350
rect 494528 280226 494848 280294
rect 494528 280170 494598 280226
rect 494654 280170 494722 280226
rect 494778 280170 494848 280226
rect 494528 280102 494848 280170
rect 494528 280046 494598 280102
rect 494654 280046 494722 280102
rect 494778 280046 494848 280102
rect 494528 279978 494848 280046
rect 494528 279922 494598 279978
rect 494654 279922 494722 279978
rect 494778 279922 494848 279978
rect 494528 279888 494848 279922
rect 525248 280350 525568 280384
rect 525248 280294 525318 280350
rect 525374 280294 525442 280350
rect 525498 280294 525568 280350
rect 525248 280226 525568 280294
rect 525248 280170 525318 280226
rect 525374 280170 525442 280226
rect 525498 280170 525568 280226
rect 525248 280102 525568 280170
rect 525248 280046 525318 280102
rect 525374 280046 525442 280102
rect 525498 280046 525568 280102
rect 525248 279978 525568 280046
rect 525248 279922 525318 279978
rect 525374 279922 525442 279978
rect 525498 279922 525568 279978
rect 525248 279888 525568 279922
rect 555968 280350 556288 280384
rect 555968 280294 556038 280350
rect 556094 280294 556162 280350
rect 556218 280294 556288 280350
rect 555968 280226 556288 280294
rect 555968 280170 556038 280226
rect 556094 280170 556162 280226
rect 556218 280170 556288 280226
rect 555968 280102 556288 280170
rect 555968 280046 556038 280102
rect 556094 280046 556162 280102
rect 556218 280046 556288 280102
rect 555968 279978 556288 280046
rect 555968 279922 556038 279978
rect 556094 279922 556162 279978
rect 556218 279922 556288 279978
rect 555968 279888 556288 279922
rect 448448 274350 448768 274384
rect 448448 274294 448518 274350
rect 448574 274294 448642 274350
rect 448698 274294 448768 274350
rect 448448 274226 448768 274294
rect 448448 274170 448518 274226
rect 448574 274170 448642 274226
rect 448698 274170 448768 274226
rect 448448 274102 448768 274170
rect 448448 274046 448518 274102
rect 448574 274046 448642 274102
rect 448698 274046 448768 274102
rect 448448 273978 448768 274046
rect 448448 273922 448518 273978
rect 448574 273922 448642 273978
rect 448698 273922 448768 273978
rect 448448 273888 448768 273922
rect 479168 274350 479488 274384
rect 479168 274294 479238 274350
rect 479294 274294 479362 274350
rect 479418 274294 479488 274350
rect 479168 274226 479488 274294
rect 479168 274170 479238 274226
rect 479294 274170 479362 274226
rect 479418 274170 479488 274226
rect 479168 274102 479488 274170
rect 479168 274046 479238 274102
rect 479294 274046 479362 274102
rect 479418 274046 479488 274102
rect 479168 273978 479488 274046
rect 479168 273922 479238 273978
rect 479294 273922 479362 273978
rect 479418 273922 479488 273978
rect 479168 273888 479488 273922
rect 509888 274350 510208 274384
rect 509888 274294 509958 274350
rect 510014 274294 510082 274350
rect 510138 274294 510208 274350
rect 509888 274226 510208 274294
rect 509888 274170 509958 274226
rect 510014 274170 510082 274226
rect 510138 274170 510208 274226
rect 509888 274102 510208 274170
rect 509888 274046 509958 274102
rect 510014 274046 510082 274102
rect 510138 274046 510208 274102
rect 509888 273978 510208 274046
rect 509888 273922 509958 273978
rect 510014 273922 510082 273978
rect 510138 273922 510208 273978
rect 509888 273888 510208 273922
rect 540608 274350 540928 274384
rect 540608 274294 540678 274350
rect 540734 274294 540802 274350
rect 540858 274294 540928 274350
rect 540608 274226 540928 274294
rect 540608 274170 540678 274226
rect 540734 274170 540802 274226
rect 540858 274170 540928 274226
rect 540608 274102 540928 274170
rect 540608 274046 540678 274102
rect 540734 274046 540802 274102
rect 540858 274046 540928 274102
rect 540608 273978 540928 274046
rect 540608 273922 540678 273978
rect 540734 273922 540802 273978
rect 540858 273922 540928 273978
rect 540608 273888 540928 273922
rect 571328 274350 571648 274384
rect 571328 274294 571398 274350
rect 571454 274294 571522 274350
rect 571578 274294 571648 274350
rect 571328 274226 571648 274294
rect 571328 274170 571398 274226
rect 571454 274170 571522 274226
rect 571578 274170 571648 274226
rect 571328 274102 571648 274170
rect 571328 274046 571398 274102
rect 571454 274046 571522 274102
rect 571578 274046 571648 274102
rect 571328 273978 571648 274046
rect 571328 273922 571398 273978
rect 571454 273922 571522 273978
rect 571578 273922 571648 273978
rect 571328 273888 571648 273922
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 463808 262350 464128 262384
rect 463808 262294 463878 262350
rect 463934 262294 464002 262350
rect 464058 262294 464128 262350
rect 463808 262226 464128 262294
rect 463808 262170 463878 262226
rect 463934 262170 464002 262226
rect 464058 262170 464128 262226
rect 463808 262102 464128 262170
rect 463808 262046 463878 262102
rect 463934 262046 464002 262102
rect 464058 262046 464128 262102
rect 463808 261978 464128 262046
rect 463808 261922 463878 261978
rect 463934 261922 464002 261978
rect 464058 261922 464128 261978
rect 463808 261888 464128 261922
rect 494528 262350 494848 262384
rect 494528 262294 494598 262350
rect 494654 262294 494722 262350
rect 494778 262294 494848 262350
rect 494528 262226 494848 262294
rect 494528 262170 494598 262226
rect 494654 262170 494722 262226
rect 494778 262170 494848 262226
rect 494528 262102 494848 262170
rect 494528 262046 494598 262102
rect 494654 262046 494722 262102
rect 494778 262046 494848 262102
rect 494528 261978 494848 262046
rect 494528 261922 494598 261978
rect 494654 261922 494722 261978
rect 494778 261922 494848 261978
rect 494528 261888 494848 261922
rect 525248 262350 525568 262384
rect 525248 262294 525318 262350
rect 525374 262294 525442 262350
rect 525498 262294 525568 262350
rect 525248 262226 525568 262294
rect 525248 262170 525318 262226
rect 525374 262170 525442 262226
rect 525498 262170 525568 262226
rect 525248 262102 525568 262170
rect 525248 262046 525318 262102
rect 525374 262046 525442 262102
rect 525498 262046 525568 262102
rect 525248 261978 525568 262046
rect 525248 261922 525318 261978
rect 525374 261922 525442 261978
rect 525498 261922 525568 261978
rect 525248 261888 525568 261922
rect 555968 262350 556288 262384
rect 555968 262294 556038 262350
rect 556094 262294 556162 262350
rect 556218 262294 556288 262350
rect 555968 262226 556288 262294
rect 555968 262170 556038 262226
rect 556094 262170 556162 262226
rect 556218 262170 556288 262226
rect 555968 262102 556288 262170
rect 555968 262046 556038 262102
rect 556094 262046 556162 262102
rect 556218 262046 556288 262102
rect 555968 261978 556288 262046
rect 555968 261922 556038 261978
rect 556094 261922 556162 261978
rect 556218 261922 556288 261978
rect 555968 261888 556288 261922
rect 587132 258244 587188 258254
rect 448448 256350 448768 256384
rect 448448 256294 448518 256350
rect 448574 256294 448642 256350
rect 448698 256294 448768 256350
rect 448448 256226 448768 256294
rect 448448 256170 448518 256226
rect 448574 256170 448642 256226
rect 448698 256170 448768 256226
rect 448448 256102 448768 256170
rect 448448 256046 448518 256102
rect 448574 256046 448642 256102
rect 448698 256046 448768 256102
rect 448448 255978 448768 256046
rect 448448 255922 448518 255978
rect 448574 255922 448642 255978
rect 448698 255922 448768 255978
rect 448448 255888 448768 255922
rect 479168 256350 479488 256384
rect 479168 256294 479238 256350
rect 479294 256294 479362 256350
rect 479418 256294 479488 256350
rect 479168 256226 479488 256294
rect 479168 256170 479238 256226
rect 479294 256170 479362 256226
rect 479418 256170 479488 256226
rect 479168 256102 479488 256170
rect 479168 256046 479238 256102
rect 479294 256046 479362 256102
rect 479418 256046 479488 256102
rect 479168 255978 479488 256046
rect 479168 255922 479238 255978
rect 479294 255922 479362 255978
rect 479418 255922 479488 255978
rect 479168 255888 479488 255922
rect 509888 256350 510208 256384
rect 509888 256294 509958 256350
rect 510014 256294 510082 256350
rect 510138 256294 510208 256350
rect 509888 256226 510208 256294
rect 509888 256170 509958 256226
rect 510014 256170 510082 256226
rect 510138 256170 510208 256226
rect 509888 256102 510208 256170
rect 509888 256046 509958 256102
rect 510014 256046 510082 256102
rect 510138 256046 510208 256102
rect 509888 255978 510208 256046
rect 509888 255922 509958 255978
rect 510014 255922 510082 255978
rect 510138 255922 510208 255978
rect 509888 255888 510208 255922
rect 540608 256350 540928 256384
rect 540608 256294 540678 256350
rect 540734 256294 540802 256350
rect 540858 256294 540928 256350
rect 540608 256226 540928 256294
rect 540608 256170 540678 256226
rect 540734 256170 540802 256226
rect 540858 256170 540928 256226
rect 540608 256102 540928 256170
rect 540608 256046 540678 256102
rect 540734 256046 540802 256102
rect 540858 256046 540928 256102
rect 540608 255978 540928 256046
rect 540608 255922 540678 255978
rect 540734 255922 540802 255978
rect 540858 255922 540928 255978
rect 540608 255888 540928 255922
rect 571328 256350 571648 256384
rect 571328 256294 571398 256350
rect 571454 256294 571522 256350
rect 571578 256294 571648 256350
rect 571328 256226 571648 256294
rect 571328 256170 571398 256226
rect 571454 256170 571522 256226
rect 571578 256170 571648 256226
rect 571328 256102 571648 256170
rect 571328 256046 571398 256102
rect 571454 256046 571522 256102
rect 571578 256046 571648 256102
rect 571328 255978 571648 256046
rect 571328 255922 571398 255978
rect 571454 255922 571522 255978
rect 571578 255922 571648 255978
rect 571328 255888 571648 255922
rect 463808 244350 464128 244384
rect 463808 244294 463878 244350
rect 463934 244294 464002 244350
rect 464058 244294 464128 244350
rect 463808 244226 464128 244294
rect 463808 244170 463878 244226
rect 463934 244170 464002 244226
rect 464058 244170 464128 244226
rect 463808 244102 464128 244170
rect 463808 244046 463878 244102
rect 463934 244046 464002 244102
rect 464058 244046 464128 244102
rect 463808 243978 464128 244046
rect 463808 243922 463878 243978
rect 463934 243922 464002 243978
rect 464058 243922 464128 243978
rect 463808 243888 464128 243922
rect 494528 244350 494848 244384
rect 494528 244294 494598 244350
rect 494654 244294 494722 244350
rect 494778 244294 494848 244350
rect 494528 244226 494848 244294
rect 494528 244170 494598 244226
rect 494654 244170 494722 244226
rect 494778 244170 494848 244226
rect 494528 244102 494848 244170
rect 494528 244046 494598 244102
rect 494654 244046 494722 244102
rect 494778 244046 494848 244102
rect 494528 243978 494848 244046
rect 494528 243922 494598 243978
rect 494654 243922 494722 243978
rect 494778 243922 494848 243978
rect 494528 243888 494848 243922
rect 525248 244350 525568 244384
rect 525248 244294 525318 244350
rect 525374 244294 525442 244350
rect 525498 244294 525568 244350
rect 525248 244226 525568 244294
rect 525248 244170 525318 244226
rect 525374 244170 525442 244226
rect 525498 244170 525568 244226
rect 525248 244102 525568 244170
rect 525248 244046 525318 244102
rect 525374 244046 525442 244102
rect 525498 244046 525568 244102
rect 525248 243978 525568 244046
rect 525248 243922 525318 243978
rect 525374 243922 525442 243978
rect 525498 243922 525568 243978
rect 525248 243888 525568 243922
rect 555968 244350 556288 244384
rect 555968 244294 556038 244350
rect 556094 244294 556162 244350
rect 556218 244294 556288 244350
rect 555968 244226 556288 244294
rect 555968 244170 556038 244226
rect 556094 244170 556162 244226
rect 556218 244170 556288 244226
rect 555968 244102 556288 244170
rect 555968 244046 556038 244102
rect 556094 244046 556162 244102
rect 556218 244046 556288 244102
rect 555968 243978 556288 244046
rect 555968 243922 556038 243978
rect 556094 243922 556162 243978
rect 556218 243922 556288 243978
rect 555968 243888 556288 243922
rect 448448 238350 448768 238384
rect 448448 238294 448518 238350
rect 448574 238294 448642 238350
rect 448698 238294 448768 238350
rect 448448 238226 448768 238294
rect 448448 238170 448518 238226
rect 448574 238170 448642 238226
rect 448698 238170 448768 238226
rect 448448 238102 448768 238170
rect 448448 238046 448518 238102
rect 448574 238046 448642 238102
rect 448698 238046 448768 238102
rect 448448 237978 448768 238046
rect 448448 237922 448518 237978
rect 448574 237922 448642 237978
rect 448698 237922 448768 237978
rect 448448 237888 448768 237922
rect 479168 238350 479488 238384
rect 479168 238294 479238 238350
rect 479294 238294 479362 238350
rect 479418 238294 479488 238350
rect 479168 238226 479488 238294
rect 479168 238170 479238 238226
rect 479294 238170 479362 238226
rect 479418 238170 479488 238226
rect 479168 238102 479488 238170
rect 479168 238046 479238 238102
rect 479294 238046 479362 238102
rect 479418 238046 479488 238102
rect 479168 237978 479488 238046
rect 479168 237922 479238 237978
rect 479294 237922 479362 237978
rect 479418 237922 479488 237978
rect 479168 237888 479488 237922
rect 509888 238350 510208 238384
rect 509888 238294 509958 238350
rect 510014 238294 510082 238350
rect 510138 238294 510208 238350
rect 509888 238226 510208 238294
rect 509888 238170 509958 238226
rect 510014 238170 510082 238226
rect 510138 238170 510208 238226
rect 509888 238102 510208 238170
rect 509888 238046 509958 238102
rect 510014 238046 510082 238102
rect 510138 238046 510208 238102
rect 509888 237978 510208 238046
rect 509888 237922 509958 237978
rect 510014 237922 510082 237978
rect 510138 237922 510208 237978
rect 509888 237888 510208 237922
rect 540608 238350 540928 238384
rect 540608 238294 540678 238350
rect 540734 238294 540802 238350
rect 540858 238294 540928 238350
rect 540608 238226 540928 238294
rect 540608 238170 540678 238226
rect 540734 238170 540802 238226
rect 540858 238170 540928 238226
rect 540608 238102 540928 238170
rect 540608 238046 540678 238102
rect 540734 238046 540802 238102
rect 540858 238046 540928 238102
rect 540608 237978 540928 238046
rect 540608 237922 540678 237978
rect 540734 237922 540802 237978
rect 540858 237922 540928 237978
rect 540608 237888 540928 237922
rect 571328 238350 571648 238384
rect 571328 238294 571398 238350
rect 571454 238294 571522 238350
rect 571578 238294 571648 238350
rect 571328 238226 571648 238294
rect 571328 238170 571398 238226
rect 571454 238170 571522 238226
rect 571578 238170 571648 238226
rect 571328 238102 571648 238170
rect 571328 238046 571398 238102
rect 571454 238046 571522 238102
rect 571578 238046 571648 238102
rect 571328 237978 571648 238046
rect 571328 237922 571398 237978
rect 571454 237922 571522 237978
rect 571578 237922 571648 237978
rect 571328 237888 571648 237922
rect 463808 226350 464128 226384
rect 463808 226294 463878 226350
rect 463934 226294 464002 226350
rect 464058 226294 464128 226350
rect 463808 226226 464128 226294
rect 463808 226170 463878 226226
rect 463934 226170 464002 226226
rect 464058 226170 464128 226226
rect 463808 226102 464128 226170
rect 463808 226046 463878 226102
rect 463934 226046 464002 226102
rect 464058 226046 464128 226102
rect 463808 225978 464128 226046
rect 463808 225922 463878 225978
rect 463934 225922 464002 225978
rect 464058 225922 464128 225978
rect 463808 225888 464128 225922
rect 494528 226350 494848 226384
rect 494528 226294 494598 226350
rect 494654 226294 494722 226350
rect 494778 226294 494848 226350
rect 494528 226226 494848 226294
rect 494528 226170 494598 226226
rect 494654 226170 494722 226226
rect 494778 226170 494848 226226
rect 494528 226102 494848 226170
rect 494528 226046 494598 226102
rect 494654 226046 494722 226102
rect 494778 226046 494848 226102
rect 494528 225978 494848 226046
rect 494528 225922 494598 225978
rect 494654 225922 494722 225978
rect 494778 225922 494848 225978
rect 494528 225888 494848 225922
rect 525248 226350 525568 226384
rect 525248 226294 525318 226350
rect 525374 226294 525442 226350
rect 525498 226294 525568 226350
rect 525248 226226 525568 226294
rect 525248 226170 525318 226226
rect 525374 226170 525442 226226
rect 525498 226170 525568 226226
rect 525248 226102 525568 226170
rect 525248 226046 525318 226102
rect 525374 226046 525442 226102
rect 525498 226046 525568 226102
rect 525248 225978 525568 226046
rect 525248 225922 525318 225978
rect 525374 225922 525442 225978
rect 525498 225922 525568 225978
rect 525248 225888 525568 225922
rect 555968 226350 556288 226384
rect 555968 226294 556038 226350
rect 556094 226294 556162 226350
rect 556218 226294 556288 226350
rect 555968 226226 556288 226294
rect 555968 226170 556038 226226
rect 556094 226170 556162 226226
rect 556218 226170 556288 226226
rect 555968 226102 556288 226170
rect 555968 226046 556038 226102
rect 556094 226046 556162 226102
rect 556218 226046 556288 226102
rect 555968 225978 556288 226046
rect 555968 225922 556038 225978
rect 556094 225922 556162 225978
rect 556218 225922 556288 225978
rect 555968 225888 556288 225922
rect 448448 220350 448768 220384
rect 448448 220294 448518 220350
rect 448574 220294 448642 220350
rect 448698 220294 448768 220350
rect 448448 220226 448768 220294
rect 448448 220170 448518 220226
rect 448574 220170 448642 220226
rect 448698 220170 448768 220226
rect 448448 220102 448768 220170
rect 448448 220046 448518 220102
rect 448574 220046 448642 220102
rect 448698 220046 448768 220102
rect 448448 219978 448768 220046
rect 448448 219922 448518 219978
rect 448574 219922 448642 219978
rect 448698 219922 448768 219978
rect 448448 219888 448768 219922
rect 479168 220350 479488 220384
rect 479168 220294 479238 220350
rect 479294 220294 479362 220350
rect 479418 220294 479488 220350
rect 479168 220226 479488 220294
rect 479168 220170 479238 220226
rect 479294 220170 479362 220226
rect 479418 220170 479488 220226
rect 479168 220102 479488 220170
rect 479168 220046 479238 220102
rect 479294 220046 479362 220102
rect 479418 220046 479488 220102
rect 479168 219978 479488 220046
rect 479168 219922 479238 219978
rect 479294 219922 479362 219978
rect 479418 219922 479488 219978
rect 479168 219888 479488 219922
rect 509888 220350 510208 220384
rect 509888 220294 509958 220350
rect 510014 220294 510082 220350
rect 510138 220294 510208 220350
rect 509888 220226 510208 220294
rect 509888 220170 509958 220226
rect 510014 220170 510082 220226
rect 510138 220170 510208 220226
rect 509888 220102 510208 220170
rect 509888 220046 509958 220102
rect 510014 220046 510082 220102
rect 510138 220046 510208 220102
rect 509888 219978 510208 220046
rect 509888 219922 509958 219978
rect 510014 219922 510082 219978
rect 510138 219922 510208 219978
rect 509888 219888 510208 219922
rect 540608 220350 540928 220384
rect 540608 220294 540678 220350
rect 540734 220294 540802 220350
rect 540858 220294 540928 220350
rect 540608 220226 540928 220294
rect 540608 220170 540678 220226
rect 540734 220170 540802 220226
rect 540858 220170 540928 220226
rect 540608 220102 540928 220170
rect 540608 220046 540678 220102
rect 540734 220046 540802 220102
rect 540858 220046 540928 220102
rect 540608 219978 540928 220046
rect 540608 219922 540678 219978
rect 540734 219922 540802 219978
rect 540858 219922 540928 219978
rect 540608 219888 540928 219922
rect 571328 220350 571648 220384
rect 571328 220294 571398 220350
rect 571454 220294 571522 220350
rect 571578 220294 571648 220350
rect 571328 220226 571648 220294
rect 571328 220170 571398 220226
rect 571454 220170 571522 220226
rect 571578 220170 571648 220226
rect 571328 220102 571648 220170
rect 571328 220046 571398 220102
rect 571454 220046 571522 220102
rect 571578 220046 571648 220102
rect 571328 219978 571648 220046
rect 571328 219922 571398 219978
rect 571454 219922 571522 219978
rect 571578 219922 571648 219978
rect 571328 219888 571648 219922
rect 463808 208350 464128 208384
rect 463808 208294 463878 208350
rect 463934 208294 464002 208350
rect 464058 208294 464128 208350
rect 463808 208226 464128 208294
rect 463808 208170 463878 208226
rect 463934 208170 464002 208226
rect 464058 208170 464128 208226
rect 463808 208102 464128 208170
rect 463808 208046 463878 208102
rect 463934 208046 464002 208102
rect 464058 208046 464128 208102
rect 463808 207978 464128 208046
rect 463808 207922 463878 207978
rect 463934 207922 464002 207978
rect 464058 207922 464128 207978
rect 463808 207888 464128 207922
rect 494528 208350 494848 208384
rect 494528 208294 494598 208350
rect 494654 208294 494722 208350
rect 494778 208294 494848 208350
rect 494528 208226 494848 208294
rect 494528 208170 494598 208226
rect 494654 208170 494722 208226
rect 494778 208170 494848 208226
rect 494528 208102 494848 208170
rect 494528 208046 494598 208102
rect 494654 208046 494722 208102
rect 494778 208046 494848 208102
rect 494528 207978 494848 208046
rect 494528 207922 494598 207978
rect 494654 207922 494722 207978
rect 494778 207922 494848 207978
rect 494528 207888 494848 207922
rect 525248 208350 525568 208384
rect 525248 208294 525318 208350
rect 525374 208294 525442 208350
rect 525498 208294 525568 208350
rect 525248 208226 525568 208294
rect 525248 208170 525318 208226
rect 525374 208170 525442 208226
rect 525498 208170 525568 208226
rect 525248 208102 525568 208170
rect 525248 208046 525318 208102
rect 525374 208046 525442 208102
rect 525498 208046 525568 208102
rect 525248 207978 525568 208046
rect 525248 207922 525318 207978
rect 525374 207922 525442 207978
rect 525498 207922 525568 207978
rect 525248 207888 525568 207922
rect 555968 208350 556288 208384
rect 555968 208294 556038 208350
rect 556094 208294 556162 208350
rect 556218 208294 556288 208350
rect 555968 208226 556288 208294
rect 555968 208170 556038 208226
rect 556094 208170 556162 208226
rect 556218 208170 556288 208226
rect 555968 208102 556288 208170
rect 555968 208046 556038 208102
rect 556094 208046 556162 208102
rect 556218 208046 556288 208102
rect 555968 207978 556288 208046
rect 555968 207922 556038 207978
rect 556094 207922 556162 207978
rect 556218 207922 556288 207978
rect 555968 207888 556288 207922
rect 448448 202350 448768 202384
rect 448448 202294 448518 202350
rect 448574 202294 448642 202350
rect 448698 202294 448768 202350
rect 448448 202226 448768 202294
rect 448448 202170 448518 202226
rect 448574 202170 448642 202226
rect 448698 202170 448768 202226
rect 448448 202102 448768 202170
rect 448448 202046 448518 202102
rect 448574 202046 448642 202102
rect 448698 202046 448768 202102
rect 448448 201978 448768 202046
rect 448448 201922 448518 201978
rect 448574 201922 448642 201978
rect 448698 201922 448768 201978
rect 448448 201888 448768 201922
rect 479168 202350 479488 202384
rect 479168 202294 479238 202350
rect 479294 202294 479362 202350
rect 479418 202294 479488 202350
rect 479168 202226 479488 202294
rect 479168 202170 479238 202226
rect 479294 202170 479362 202226
rect 479418 202170 479488 202226
rect 479168 202102 479488 202170
rect 479168 202046 479238 202102
rect 479294 202046 479362 202102
rect 479418 202046 479488 202102
rect 479168 201978 479488 202046
rect 479168 201922 479238 201978
rect 479294 201922 479362 201978
rect 479418 201922 479488 201978
rect 479168 201888 479488 201922
rect 509888 202350 510208 202384
rect 509888 202294 509958 202350
rect 510014 202294 510082 202350
rect 510138 202294 510208 202350
rect 509888 202226 510208 202294
rect 509888 202170 509958 202226
rect 510014 202170 510082 202226
rect 510138 202170 510208 202226
rect 509888 202102 510208 202170
rect 509888 202046 509958 202102
rect 510014 202046 510082 202102
rect 510138 202046 510208 202102
rect 509888 201978 510208 202046
rect 509888 201922 509958 201978
rect 510014 201922 510082 201978
rect 510138 201922 510208 201978
rect 509888 201888 510208 201922
rect 540608 202350 540928 202384
rect 540608 202294 540678 202350
rect 540734 202294 540802 202350
rect 540858 202294 540928 202350
rect 540608 202226 540928 202294
rect 540608 202170 540678 202226
rect 540734 202170 540802 202226
rect 540858 202170 540928 202226
rect 540608 202102 540928 202170
rect 540608 202046 540678 202102
rect 540734 202046 540802 202102
rect 540858 202046 540928 202102
rect 540608 201978 540928 202046
rect 540608 201922 540678 201978
rect 540734 201922 540802 201978
rect 540858 201922 540928 201978
rect 540608 201888 540928 201922
rect 571328 202350 571648 202384
rect 571328 202294 571398 202350
rect 571454 202294 571522 202350
rect 571578 202294 571648 202350
rect 571328 202226 571648 202294
rect 571328 202170 571398 202226
rect 571454 202170 571522 202226
rect 571578 202170 571648 202226
rect 571328 202102 571648 202170
rect 571328 202046 571398 202102
rect 571454 202046 571522 202102
rect 571578 202046 571648 202102
rect 571328 201978 571648 202046
rect 571328 201922 571398 201978
rect 571454 201922 571522 201978
rect 571578 201922 571648 201978
rect 571328 201888 571648 201922
rect 463808 190350 464128 190384
rect 463808 190294 463878 190350
rect 463934 190294 464002 190350
rect 464058 190294 464128 190350
rect 463808 190226 464128 190294
rect 463808 190170 463878 190226
rect 463934 190170 464002 190226
rect 464058 190170 464128 190226
rect 463808 190102 464128 190170
rect 463808 190046 463878 190102
rect 463934 190046 464002 190102
rect 464058 190046 464128 190102
rect 463808 189978 464128 190046
rect 463808 189922 463878 189978
rect 463934 189922 464002 189978
rect 464058 189922 464128 189978
rect 463808 189888 464128 189922
rect 494528 190350 494848 190384
rect 494528 190294 494598 190350
rect 494654 190294 494722 190350
rect 494778 190294 494848 190350
rect 494528 190226 494848 190294
rect 494528 190170 494598 190226
rect 494654 190170 494722 190226
rect 494778 190170 494848 190226
rect 494528 190102 494848 190170
rect 494528 190046 494598 190102
rect 494654 190046 494722 190102
rect 494778 190046 494848 190102
rect 494528 189978 494848 190046
rect 494528 189922 494598 189978
rect 494654 189922 494722 189978
rect 494778 189922 494848 189978
rect 494528 189888 494848 189922
rect 525248 190350 525568 190384
rect 525248 190294 525318 190350
rect 525374 190294 525442 190350
rect 525498 190294 525568 190350
rect 525248 190226 525568 190294
rect 525248 190170 525318 190226
rect 525374 190170 525442 190226
rect 525498 190170 525568 190226
rect 525248 190102 525568 190170
rect 525248 190046 525318 190102
rect 525374 190046 525442 190102
rect 525498 190046 525568 190102
rect 525248 189978 525568 190046
rect 525248 189922 525318 189978
rect 525374 189922 525442 189978
rect 525498 189922 525568 189978
rect 525248 189888 525568 189922
rect 555968 190350 556288 190384
rect 555968 190294 556038 190350
rect 556094 190294 556162 190350
rect 556218 190294 556288 190350
rect 555968 190226 556288 190294
rect 555968 190170 556038 190226
rect 556094 190170 556162 190226
rect 556218 190170 556288 190226
rect 555968 190102 556288 190170
rect 555968 190046 556038 190102
rect 556094 190046 556162 190102
rect 556218 190046 556288 190102
rect 555968 189978 556288 190046
rect 555968 189922 556038 189978
rect 556094 189922 556162 189978
rect 556218 189922 556288 189978
rect 555968 189888 556288 189922
rect 448448 184350 448768 184384
rect 448448 184294 448518 184350
rect 448574 184294 448642 184350
rect 448698 184294 448768 184350
rect 448448 184226 448768 184294
rect 448448 184170 448518 184226
rect 448574 184170 448642 184226
rect 448698 184170 448768 184226
rect 448448 184102 448768 184170
rect 448448 184046 448518 184102
rect 448574 184046 448642 184102
rect 448698 184046 448768 184102
rect 448448 183978 448768 184046
rect 448448 183922 448518 183978
rect 448574 183922 448642 183978
rect 448698 183922 448768 183978
rect 448448 183888 448768 183922
rect 479168 184350 479488 184384
rect 479168 184294 479238 184350
rect 479294 184294 479362 184350
rect 479418 184294 479488 184350
rect 479168 184226 479488 184294
rect 479168 184170 479238 184226
rect 479294 184170 479362 184226
rect 479418 184170 479488 184226
rect 479168 184102 479488 184170
rect 479168 184046 479238 184102
rect 479294 184046 479362 184102
rect 479418 184046 479488 184102
rect 479168 183978 479488 184046
rect 479168 183922 479238 183978
rect 479294 183922 479362 183978
rect 479418 183922 479488 183978
rect 479168 183888 479488 183922
rect 509888 184350 510208 184384
rect 509888 184294 509958 184350
rect 510014 184294 510082 184350
rect 510138 184294 510208 184350
rect 509888 184226 510208 184294
rect 509888 184170 509958 184226
rect 510014 184170 510082 184226
rect 510138 184170 510208 184226
rect 509888 184102 510208 184170
rect 509888 184046 509958 184102
rect 510014 184046 510082 184102
rect 510138 184046 510208 184102
rect 509888 183978 510208 184046
rect 509888 183922 509958 183978
rect 510014 183922 510082 183978
rect 510138 183922 510208 183978
rect 509888 183888 510208 183922
rect 540608 184350 540928 184384
rect 540608 184294 540678 184350
rect 540734 184294 540802 184350
rect 540858 184294 540928 184350
rect 540608 184226 540928 184294
rect 540608 184170 540678 184226
rect 540734 184170 540802 184226
rect 540858 184170 540928 184226
rect 540608 184102 540928 184170
rect 540608 184046 540678 184102
rect 540734 184046 540802 184102
rect 540858 184046 540928 184102
rect 540608 183978 540928 184046
rect 540608 183922 540678 183978
rect 540734 183922 540802 183978
rect 540858 183922 540928 183978
rect 540608 183888 540928 183922
rect 571328 184350 571648 184384
rect 571328 184294 571398 184350
rect 571454 184294 571522 184350
rect 571578 184294 571648 184350
rect 571328 184226 571648 184294
rect 571328 184170 571398 184226
rect 571454 184170 571522 184226
rect 571578 184170 571648 184226
rect 571328 184102 571648 184170
rect 571328 184046 571398 184102
rect 571454 184046 571522 184102
rect 571578 184046 571648 184102
rect 571328 183978 571648 184046
rect 571328 183922 571398 183978
rect 571454 183922 571522 183978
rect 571578 183922 571648 183978
rect 571328 183888 571648 183922
rect 463808 172350 464128 172384
rect 463808 172294 463878 172350
rect 463934 172294 464002 172350
rect 464058 172294 464128 172350
rect 463808 172226 464128 172294
rect 463808 172170 463878 172226
rect 463934 172170 464002 172226
rect 464058 172170 464128 172226
rect 463808 172102 464128 172170
rect 463808 172046 463878 172102
rect 463934 172046 464002 172102
rect 464058 172046 464128 172102
rect 463808 171978 464128 172046
rect 463808 171922 463878 171978
rect 463934 171922 464002 171978
rect 464058 171922 464128 171978
rect 463808 171888 464128 171922
rect 494528 172350 494848 172384
rect 494528 172294 494598 172350
rect 494654 172294 494722 172350
rect 494778 172294 494848 172350
rect 494528 172226 494848 172294
rect 494528 172170 494598 172226
rect 494654 172170 494722 172226
rect 494778 172170 494848 172226
rect 494528 172102 494848 172170
rect 494528 172046 494598 172102
rect 494654 172046 494722 172102
rect 494778 172046 494848 172102
rect 494528 171978 494848 172046
rect 494528 171922 494598 171978
rect 494654 171922 494722 171978
rect 494778 171922 494848 171978
rect 494528 171888 494848 171922
rect 525248 172350 525568 172384
rect 525248 172294 525318 172350
rect 525374 172294 525442 172350
rect 525498 172294 525568 172350
rect 525248 172226 525568 172294
rect 525248 172170 525318 172226
rect 525374 172170 525442 172226
rect 525498 172170 525568 172226
rect 525248 172102 525568 172170
rect 525248 172046 525318 172102
rect 525374 172046 525442 172102
rect 525498 172046 525568 172102
rect 525248 171978 525568 172046
rect 525248 171922 525318 171978
rect 525374 171922 525442 171978
rect 525498 171922 525568 171978
rect 525248 171888 525568 171922
rect 555968 172350 556288 172384
rect 555968 172294 556038 172350
rect 556094 172294 556162 172350
rect 556218 172294 556288 172350
rect 555968 172226 556288 172294
rect 555968 172170 556038 172226
rect 556094 172170 556162 172226
rect 556218 172170 556288 172226
rect 555968 172102 556288 172170
rect 555968 172046 556038 172102
rect 556094 172046 556162 172102
rect 556218 172046 556288 172102
rect 555968 171978 556288 172046
rect 555968 171922 556038 171978
rect 556094 171922 556162 171978
rect 556218 171922 556288 171978
rect 555968 171888 556288 171922
rect 448448 166350 448768 166384
rect 448448 166294 448518 166350
rect 448574 166294 448642 166350
rect 448698 166294 448768 166350
rect 448448 166226 448768 166294
rect 448448 166170 448518 166226
rect 448574 166170 448642 166226
rect 448698 166170 448768 166226
rect 448448 166102 448768 166170
rect 448448 166046 448518 166102
rect 448574 166046 448642 166102
rect 448698 166046 448768 166102
rect 448448 165978 448768 166046
rect 448448 165922 448518 165978
rect 448574 165922 448642 165978
rect 448698 165922 448768 165978
rect 448448 165888 448768 165922
rect 479168 166350 479488 166384
rect 479168 166294 479238 166350
rect 479294 166294 479362 166350
rect 479418 166294 479488 166350
rect 479168 166226 479488 166294
rect 479168 166170 479238 166226
rect 479294 166170 479362 166226
rect 479418 166170 479488 166226
rect 479168 166102 479488 166170
rect 479168 166046 479238 166102
rect 479294 166046 479362 166102
rect 479418 166046 479488 166102
rect 479168 165978 479488 166046
rect 479168 165922 479238 165978
rect 479294 165922 479362 165978
rect 479418 165922 479488 165978
rect 479168 165888 479488 165922
rect 509888 166350 510208 166384
rect 509888 166294 509958 166350
rect 510014 166294 510082 166350
rect 510138 166294 510208 166350
rect 509888 166226 510208 166294
rect 509888 166170 509958 166226
rect 510014 166170 510082 166226
rect 510138 166170 510208 166226
rect 509888 166102 510208 166170
rect 509888 166046 509958 166102
rect 510014 166046 510082 166102
rect 510138 166046 510208 166102
rect 509888 165978 510208 166046
rect 509888 165922 509958 165978
rect 510014 165922 510082 165978
rect 510138 165922 510208 165978
rect 509888 165888 510208 165922
rect 540608 166350 540928 166384
rect 540608 166294 540678 166350
rect 540734 166294 540802 166350
rect 540858 166294 540928 166350
rect 540608 166226 540928 166294
rect 540608 166170 540678 166226
rect 540734 166170 540802 166226
rect 540858 166170 540928 166226
rect 540608 166102 540928 166170
rect 540608 166046 540678 166102
rect 540734 166046 540802 166102
rect 540858 166046 540928 166102
rect 540608 165978 540928 166046
rect 540608 165922 540678 165978
rect 540734 165922 540802 165978
rect 540858 165922 540928 165978
rect 540608 165888 540928 165922
rect 571328 166350 571648 166384
rect 571328 166294 571398 166350
rect 571454 166294 571522 166350
rect 571578 166294 571648 166350
rect 571328 166226 571648 166294
rect 571328 166170 571398 166226
rect 571454 166170 571522 166226
rect 571578 166170 571648 166226
rect 571328 166102 571648 166170
rect 571328 166046 571398 166102
rect 571454 166046 571522 166102
rect 571578 166046 571648 166102
rect 571328 165978 571648 166046
rect 571328 165922 571398 165978
rect 571454 165922 571522 165978
rect 571578 165922 571648 165978
rect 571328 165888 571648 165922
rect 463808 154350 464128 154384
rect 463808 154294 463878 154350
rect 463934 154294 464002 154350
rect 464058 154294 464128 154350
rect 463808 154226 464128 154294
rect 463808 154170 463878 154226
rect 463934 154170 464002 154226
rect 464058 154170 464128 154226
rect 463808 154102 464128 154170
rect 463808 154046 463878 154102
rect 463934 154046 464002 154102
rect 464058 154046 464128 154102
rect 463808 153978 464128 154046
rect 463808 153922 463878 153978
rect 463934 153922 464002 153978
rect 464058 153922 464128 153978
rect 463808 153888 464128 153922
rect 494528 154350 494848 154384
rect 494528 154294 494598 154350
rect 494654 154294 494722 154350
rect 494778 154294 494848 154350
rect 494528 154226 494848 154294
rect 494528 154170 494598 154226
rect 494654 154170 494722 154226
rect 494778 154170 494848 154226
rect 494528 154102 494848 154170
rect 494528 154046 494598 154102
rect 494654 154046 494722 154102
rect 494778 154046 494848 154102
rect 494528 153978 494848 154046
rect 494528 153922 494598 153978
rect 494654 153922 494722 153978
rect 494778 153922 494848 153978
rect 494528 153888 494848 153922
rect 525248 154350 525568 154384
rect 525248 154294 525318 154350
rect 525374 154294 525442 154350
rect 525498 154294 525568 154350
rect 525248 154226 525568 154294
rect 525248 154170 525318 154226
rect 525374 154170 525442 154226
rect 525498 154170 525568 154226
rect 525248 154102 525568 154170
rect 525248 154046 525318 154102
rect 525374 154046 525442 154102
rect 525498 154046 525568 154102
rect 525248 153978 525568 154046
rect 525248 153922 525318 153978
rect 525374 153922 525442 153978
rect 525498 153922 525568 153978
rect 525248 153888 525568 153922
rect 555968 154350 556288 154384
rect 555968 154294 556038 154350
rect 556094 154294 556162 154350
rect 556218 154294 556288 154350
rect 555968 154226 556288 154294
rect 555968 154170 556038 154226
rect 556094 154170 556162 154226
rect 556218 154170 556288 154226
rect 555968 154102 556288 154170
rect 555968 154046 556038 154102
rect 556094 154046 556162 154102
rect 556218 154046 556288 154102
rect 555968 153978 556288 154046
rect 555968 153922 556038 153978
rect 556094 153922 556162 153978
rect 556218 153922 556288 153978
rect 555968 153888 556288 153922
rect 448448 148350 448768 148384
rect 448448 148294 448518 148350
rect 448574 148294 448642 148350
rect 448698 148294 448768 148350
rect 448448 148226 448768 148294
rect 448448 148170 448518 148226
rect 448574 148170 448642 148226
rect 448698 148170 448768 148226
rect 448448 148102 448768 148170
rect 448448 148046 448518 148102
rect 448574 148046 448642 148102
rect 448698 148046 448768 148102
rect 448448 147978 448768 148046
rect 448448 147922 448518 147978
rect 448574 147922 448642 147978
rect 448698 147922 448768 147978
rect 448448 147888 448768 147922
rect 479168 148350 479488 148384
rect 479168 148294 479238 148350
rect 479294 148294 479362 148350
rect 479418 148294 479488 148350
rect 479168 148226 479488 148294
rect 479168 148170 479238 148226
rect 479294 148170 479362 148226
rect 479418 148170 479488 148226
rect 479168 148102 479488 148170
rect 479168 148046 479238 148102
rect 479294 148046 479362 148102
rect 479418 148046 479488 148102
rect 479168 147978 479488 148046
rect 479168 147922 479238 147978
rect 479294 147922 479362 147978
rect 479418 147922 479488 147978
rect 479168 147888 479488 147922
rect 509888 148350 510208 148384
rect 509888 148294 509958 148350
rect 510014 148294 510082 148350
rect 510138 148294 510208 148350
rect 509888 148226 510208 148294
rect 509888 148170 509958 148226
rect 510014 148170 510082 148226
rect 510138 148170 510208 148226
rect 509888 148102 510208 148170
rect 509888 148046 509958 148102
rect 510014 148046 510082 148102
rect 510138 148046 510208 148102
rect 509888 147978 510208 148046
rect 509888 147922 509958 147978
rect 510014 147922 510082 147978
rect 510138 147922 510208 147978
rect 509888 147888 510208 147922
rect 540608 148350 540928 148384
rect 540608 148294 540678 148350
rect 540734 148294 540802 148350
rect 540858 148294 540928 148350
rect 540608 148226 540928 148294
rect 540608 148170 540678 148226
rect 540734 148170 540802 148226
rect 540858 148170 540928 148226
rect 540608 148102 540928 148170
rect 540608 148046 540678 148102
rect 540734 148046 540802 148102
rect 540858 148046 540928 148102
rect 540608 147978 540928 148046
rect 540608 147922 540678 147978
rect 540734 147922 540802 147978
rect 540858 147922 540928 147978
rect 540608 147888 540928 147922
rect 571328 148350 571648 148384
rect 571328 148294 571398 148350
rect 571454 148294 571522 148350
rect 571578 148294 571648 148350
rect 571328 148226 571648 148294
rect 571328 148170 571398 148226
rect 571454 148170 571522 148226
rect 571578 148170 571648 148226
rect 571328 148102 571648 148170
rect 571328 148046 571398 148102
rect 571454 148046 571522 148102
rect 571578 148046 571648 148102
rect 571328 147978 571648 148046
rect 571328 147922 571398 147978
rect 571454 147922 571522 147978
rect 571578 147922 571648 147978
rect 571328 147888 571648 147922
rect 463808 136350 464128 136384
rect 463808 136294 463878 136350
rect 463934 136294 464002 136350
rect 464058 136294 464128 136350
rect 463808 136226 464128 136294
rect 463808 136170 463878 136226
rect 463934 136170 464002 136226
rect 464058 136170 464128 136226
rect 463808 136102 464128 136170
rect 463808 136046 463878 136102
rect 463934 136046 464002 136102
rect 464058 136046 464128 136102
rect 463808 135978 464128 136046
rect 463808 135922 463878 135978
rect 463934 135922 464002 135978
rect 464058 135922 464128 135978
rect 463808 135888 464128 135922
rect 494528 136350 494848 136384
rect 494528 136294 494598 136350
rect 494654 136294 494722 136350
rect 494778 136294 494848 136350
rect 494528 136226 494848 136294
rect 494528 136170 494598 136226
rect 494654 136170 494722 136226
rect 494778 136170 494848 136226
rect 494528 136102 494848 136170
rect 494528 136046 494598 136102
rect 494654 136046 494722 136102
rect 494778 136046 494848 136102
rect 494528 135978 494848 136046
rect 494528 135922 494598 135978
rect 494654 135922 494722 135978
rect 494778 135922 494848 135978
rect 494528 135888 494848 135922
rect 525248 136350 525568 136384
rect 525248 136294 525318 136350
rect 525374 136294 525442 136350
rect 525498 136294 525568 136350
rect 525248 136226 525568 136294
rect 525248 136170 525318 136226
rect 525374 136170 525442 136226
rect 525498 136170 525568 136226
rect 525248 136102 525568 136170
rect 525248 136046 525318 136102
rect 525374 136046 525442 136102
rect 525498 136046 525568 136102
rect 525248 135978 525568 136046
rect 525248 135922 525318 135978
rect 525374 135922 525442 135978
rect 525498 135922 525568 135978
rect 525248 135888 525568 135922
rect 555968 136350 556288 136384
rect 555968 136294 556038 136350
rect 556094 136294 556162 136350
rect 556218 136294 556288 136350
rect 555968 136226 556288 136294
rect 555968 136170 556038 136226
rect 556094 136170 556162 136226
rect 556218 136170 556288 136226
rect 555968 136102 556288 136170
rect 555968 136046 556038 136102
rect 556094 136046 556162 136102
rect 556218 136046 556288 136102
rect 555968 135978 556288 136046
rect 555968 135922 556038 135978
rect 556094 135922 556162 135978
rect 556218 135922 556288 135978
rect 555968 135888 556288 135922
rect 448448 130350 448768 130384
rect 448448 130294 448518 130350
rect 448574 130294 448642 130350
rect 448698 130294 448768 130350
rect 448448 130226 448768 130294
rect 448448 130170 448518 130226
rect 448574 130170 448642 130226
rect 448698 130170 448768 130226
rect 448448 130102 448768 130170
rect 448448 130046 448518 130102
rect 448574 130046 448642 130102
rect 448698 130046 448768 130102
rect 448448 129978 448768 130046
rect 448448 129922 448518 129978
rect 448574 129922 448642 129978
rect 448698 129922 448768 129978
rect 448448 129888 448768 129922
rect 479168 130350 479488 130384
rect 479168 130294 479238 130350
rect 479294 130294 479362 130350
rect 479418 130294 479488 130350
rect 479168 130226 479488 130294
rect 479168 130170 479238 130226
rect 479294 130170 479362 130226
rect 479418 130170 479488 130226
rect 479168 130102 479488 130170
rect 479168 130046 479238 130102
rect 479294 130046 479362 130102
rect 479418 130046 479488 130102
rect 479168 129978 479488 130046
rect 479168 129922 479238 129978
rect 479294 129922 479362 129978
rect 479418 129922 479488 129978
rect 479168 129888 479488 129922
rect 509888 130350 510208 130384
rect 509888 130294 509958 130350
rect 510014 130294 510082 130350
rect 510138 130294 510208 130350
rect 509888 130226 510208 130294
rect 509888 130170 509958 130226
rect 510014 130170 510082 130226
rect 510138 130170 510208 130226
rect 509888 130102 510208 130170
rect 509888 130046 509958 130102
rect 510014 130046 510082 130102
rect 510138 130046 510208 130102
rect 509888 129978 510208 130046
rect 509888 129922 509958 129978
rect 510014 129922 510082 129978
rect 510138 129922 510208 129978
rect 509888 129888 510208 129922
rect 540608 130350 540928 130384
rect 540608 130294 540678 130350
rect 540734 130294 540802 130350
rect 540858 130294 540928 130350
rect 540608 130226 540928 130294
rect 540608 130170 540678 130226
rect 540734 130170 540802 130226
rect 540858 130170 540928 130226
rect 540608 130102 540928 130170
rect 540608 130046 540678 130102
rect 540734 130046 540802 130102
rect 540858 130046 540928 130102
rect 540608 129978 540928 130046
rect 540608 129922 540678 129978
rect 540734 129922 540802 129978
rect 540858 129922 540928 129978
rect 540608 129888 540928 129922
rect 571328 130350 571648 130384
rect 571328 130294 571398 130350
rect 571454 130294 571522 130350
rect 571578 130294 571648 130350
rect 571328 130226 571648 130294
rect 571328 130170 571398 130226
rect 571454 130170 571522 130226
rect 571578 130170 571648 130226
rect 571328 130102 571648 130170
rect 571328 130046 571398 130102
rect 571454 130046 571522 130102
rect 571578 130046 571648 130102
rect 571328 129978 571648 130046
rect 571328 129922 571398 129978
rect 571454 129922 571522 129978
rect 571578 129922 571648 129978
rect 571328 129888 571648 129922
rect 463808 118350 464128 118384
rect 463808 118294 463878 118350
rect 463934 118294 464002 118350
rect 464058 118294 464128 118350
rect 463808 118226 464128 118294
rect 463808 118170 463878 118226
rect 463934 118170 464002 118226
rect 464058 118170 464128 118226
rect 463808 118102 464128 118170
rect 463808 118046 463878 118102
rect 463934 118046 464002 118102
rect 464058 118046 464128 118102
rect 463808 117978 464128 118046
rect 463808 117922 463878 117978
rect 463934 117922 464002 117978
rect 464058 117922 464128 117978
rect 463808 117888 464128 117922
rect 494528 118350 494848 118384
rect 494528 118294 494598 118350
rect 494654 118294 494722 118350
rect 494778 118294 494848 118350
rect 494528 118226 494848 118294
rect 494528 118170 494598 118226
rect 494654 118170 494722 118226
rect 494778 118170 494848 118226
rect 494528 118102 494848 118170
rect 494528 118046 494598 118102
rect 494654 118046 494722 118102
rect 494778 118046 494848 118102
rect 494528 117978 494848 118046
rect 494528 117922 494598 117978
rect 494654 117922 494722 117978
rect 494778 117922 494848 117978
rect 494528 117888 494848 117922
rect 525248 118350 525568 118384
rect 525248 118294 525318 118350
rect 525374 118294 525442 118350
rect 525498 118294 525568 118350
rect 525248 118226 525568 118294
rect 525248 118170 525318 118226
rect 525374 118170 525442 118226
rect 525498 118170 525568 118226
rect 525248 118102 525568 118170
rect 525248 118046 525318 118102
rect 525374 118046 525442 118102
rect 525498 118046 525568 118102
rect 525248 117978 525568 118046
rect 525248 117922 525318 117978
rect 525374 117922 525442 117978
rect 525498 117922 525568 117978
rect 525248 117888 525568 117922
rect 555968 118350 556288 118384
rect 555968 118294 556038 118350
rect 556094 118294 556162 118350
rect 556218 118294 556288 118350
rect 555968 118226 556288 118294
rect 555968 118170 556038 118226
rect 556094 118170 556162 118226
rect 556218 118170 556288 118226
rect 555968 118102 556288 118170
rect 555968 118046 556038 118102
rect 556094 118046 556162 118102
rect 556218 118046 556288 118102
rect 555968 117978 556288 118046
rect 555968 117922 556038 117978
rect 556094 117922 556162 117978
rect 556218 117922 556288 117978
rect 555968 117888 556288 117922
rect 448448 112350 448768 112384
rect 448448 112294 448518 112350
rect 448574 112294 448642 112350
rect 448698 112294 448768 112350
rect 448448 112226 448768 112294
rect 448448 112170 448518 112226
rect 448574 112170 448642 112226
rect 448698 112170 448768 112226
rect 448448 112102 448768 112170
rect 448448 112046 448518 112102
rect 448574 112046 448642 112102
rect 448698 112046 448768 112102
rect 448448 111978 448768 112046
rect 448448 111922 448518 111978
rect 448574 111922 448642 111978
rect 448698 111922 448768 111978
rect 448448 111888 448768 111922
rect 479168 112350 479488 112384
rect 479168 112294 479238 112350
rect 479294 112294 479362 112350
rect 479418 112294 479488 112350
rect 479168 112226 479488 112294
rect 479168 112170 479238 112226
rect 479294 112170 479362 112226
rect 479418 112170 479488 112226
rect 479168 112102 479488 112170
rect 479168 112046 479238 112102
rect 479294 112046 479362 112102
rect 479418 112046 479488 112102
rect 479168 111978 479488 112046
rect 479168 111922 479238 111978
rect 479294 111922 479362 111978
rect 479418 111922 479488 111978
rect 479168 111888 479488 111922
rect 509888 112350 510208 112384
rect 509888 112294 509958 112350
rect 510014 112294 510082 112350
rect 510138 112294 510208 112350
rect 509888 112226 510208 112294
rect 509888 112170 509958 112226
rect 510014 112170 510082 112226
rect 510138 112170 510208 112226
rect 509888 112102 510208 112170
rect 509888 112046 509958 112102
rect 510014 112046 510082 112102
rect 510138 112046 510208 112102
rect 509888 111978 510208 112046
rect 509888 111922 509958 111978
rect 510014 111922 510082 111978
rect 510138 111922 510208 111978
rect 509888 111888 510208 111922
rect 540608 112350 540928 112384
rect 540608 112294 540678 112350
rect 540734 112294 540802 112350
rect 540858 112294 540928 112350
rect 540608 112226 540928 112294
rect 540608 112170 540678 112226
rect 540734 112170 540802 112226
rect 540858 112170 540928 112226
rect 540608 112102 540928 112170
rect 540608 112046 540678 112102
rect 540734 112046 540802 112102
rect 540858 112046 540928 112102
rect 540608 111978 540928 112046
rect 540608 111922 540678 111978
rect 540734 111922 540802 111978
rect 540858 111922 540928 111978
rect 540608 111888 540928 111922
rect 571328 112350 571648 112384
rect 571328 112294 571398 112350
rect 571454 112294 571522 112350
rect 571578 112294 571648 112350
rect 571328 112226 571648 112294
rect 571328 112170 571398 112226
rect 571454 112170 571522 112226
rect 571578 112170 571648 112226
rect 571328 112102 571648 112170
rect 571328 112046 571398 112102
rect 571454 112046 571522 112102
rect 571578 112046 571648 112102
rect 571328 111978 571648 112046
rect 571328 111922 571398 111978
rect 571454 111922 571522 111978
rect 571578 111922 571648 111978
rect 571328 111888 571648 111922
rect 443436 101572 443492 101582
rect 463808 100350 464128 100384
rect 463808 100294 463878 100350
rect 463934 100294 464002 100350
rect 464058 100294 464128 100350
rect 463808 100226 464128 100294
rect 463808 100170 463878 100226
rect 463934 100170 464002 100226
rect 464058 100170 464128 100226
rect 463808 100102 464128 100170
rect 463808 100046 463878 100102
rect 463934 100046 464002 100102
rect 464058 100046 464128 100102
rect 463808 99978 464128 100046
rect 463808 99922 463878 99978
rect 463934 99922 464002 99978
rect 464058 99922 464128 99978
rect 463808 99888 464128 99922
rect 494528 100350 494848 100384
rect 494528 100294 494598 100350
rect 494654 100294 494722 100350
rect 494778 100294 494848 100350
rect 494528 100226 494848 100294
rect 494528 100170 494598 100226
rect 494654 100170 494722 100226
rect 494778 100170 494848 100226
rect 494528 100102 494848 100170
rect 494528 100046 494598 100102
rect 494654 100046 494722 100102
rect 494778 100046 494848 100102
rect 494528 99978 494848 100046
rect 494528 99922 494598 99978
rect 494654 99922 494722 99978
rect 494778 99922 494848 99978
rect 494528 99888 494848 99922
rect 525248 100350 525568 100384
rect 525248 100294 525318 100350
rect 525374 100294 525442 100350
rect 525498 100294 525568 100350
rect 525248 100226 525568 100294
rect 525248 100170 525318 100226
rect 525374 100170 525442 100226
rect 525498 100170 525568 100226
rect 525248 100102 525568 100170
rect 525248 100046 525318 100102
rect 525374 100046 525442 100102
rect 525498 100046 525568 100102
rect 525248 99978 525568 100046
rect 525248 99922 525318 99978
rect 525374 99922 525442 99978
rect 525498 99922 525568 99978
rect 525248 99888 525568 99922
rect 555968 100350 556288 100384
rect 555968 100294 556038 100350
rect 556094 100294 556162 100350
rect 556218 100294 556288 100350
rect 555968 100226 556288 100294
rect 555968 100170 556038 100226
rect 556094 100170 556162 100226
rect 556218 100170 556288 100226
rect 555968 100102 556288 100170
rect 555968 100046 556038 100102
rect 556094 100046 556162 100102
rect 556218 100046 556288 100102
rect 555968 99978 556288 100046
rect 555968 99922 556038 99978
rect 556094 99922 556162 99978
rect 556218 99922 556288 99978
rect 555968 99888 556288 99922
rect 443100 98152 443156 98162
rect 448448 94350 448768 94384
rect 448448 94294 448518 94350
rect 448574 94294 448642 94350
rect 448698 94294 448768 94350
rect 448448 94226 448768 94294
rect 448448 94170 448518 94226
rect 448574 94170 448642 94226
rect 448698 94170 448768 94226
rect 448448 94102 448768 94170
rect 448448 94046 448518 94102
rect 448574 94046 448642 94102
rect 448698 94046 448768 94102
rect 448448 93978 448768 94046
rect 448448 93922 448518 93978
rect 448574 93922 448642 93978
rect 448698 93922 448768 93978
rect 448448 93888 448768 93922
rect 479168 94350 479488 94384
rect 479168 94294 479238 94350
rect 479294 94294 479362 94350
rect 479418 94294 479488 94350
rect 479168 94226 479488 94294
rect 479168 94170 479238 94226
rect 479294 94170 479362 94226
rect 479418 94170 479488 94226
rect 479168 94102 479488 94170
rect 479168 94046 479238 94102
rect 479294 94046 479362 94102
rect 479418 94046 479488 94102
rect 479168 93978 479488 94046
rect 479168 93922 479238 93978
rect 479294 93922 479362 93978
rect 479418 93922 479488 93978
rect 479168 93888 479488 93922
rect 509888 94350 510208 94384
rect 509888 94294 509958 94350
rect 510014 94294 510082 94350
rect 510138 94294 510208 94350
rect 509888 94226 510208 94294
rect 509888 94170 509958 94226
rect 510014 94170 510082 94226
rect 510138 94170 510208 94226
rect 509888 94102 510208 94170
rect 509888 94046 509958 94102
rect 510014 94046 510082 94102
rect 510138 94046 510208 94102
rect 509888 93978 510208 94046
rect 509888 93922 509958 93978
rect 510014 93922 510082 93978
rect 510138 93922 510208 93978
rect 509888 93888 510208 93922
rect 540608 94350 540928 94384
rect 540608 94294 540678 94350
rect 540734 94294 540802 94350
rect 540858 94294 540928 94350
rect 540608 94226 540928 94294
rect 540608 94170 540678 94226
rect 540734 94170 540802 94226
rect 540858 94170 540928 94226
rect 540608 94102 540928 94170
rect 540608 94046 540678 94102
rect 540734 94046 540802 94102
rect 540858 94046 540928 94102
rect 540608 93978 540928 94046
rect 540608 93922 540678 93978
rect 540734 93922 540802 93978
rect 540858 93922 540928 93978
rect 540608 93888 540928 93922
rect 571328 94350 571648 94384
rect 571328 94294 571398 94350
rect 571454 94294 571522 94350
rect 571578 94294 571648 94350
rect 571328 94226 571648 94294
rect 571328 94170 571398 94226
rect 571454 94170 571522 94226
rect 571578 94170 571648 94226
rect 571328 94102 571648 94170
rect 571328 94046 571398 94102
rect 571454 94046 571522 94102
rect 571578 94046 571648 94102
rect 571328 93978 571648 94046
rect 571328 93922 571398 93978
rect 571454 93922 571522 93978
rect 571578 93922 571648 93978
rect 571328 93888 571648 93922
rect 443100 85798 443156 85808
rect 443100 16212 443156 85742
rect 463808 82350 464128 82384
rect 463808 82294 463878 82350
rect 463934 82294 464002 82350
rect 464058 82294 464128 82350
rect 463808 82226 464128 82294
rect 463808 82170 463878 82226
rect 463934 82170 464002 82226
rect 464058 82170 464128 82226
rect 463808 82102 464128 82170
rect 463808 82046 463878 82102
rect 463934 82046 464002 82102
rect 464058 82046 464128 82102
rect 463808 81978 464128 82046
rect 463808 81922 463878 81978
rect 463934 81922 464002 81978
rect 464058 81922 464128 81978
rect 463808 81888 464128 81922
rect 494528 82350 494848 82384
rect 494528 82294 494598 82350
rect 494654 82294 494722 82350
rect 494778 82294 494848 82350
rect 494528 82226 494848 82294
rect 494528 82170 494598 82226
rect 494654 82170 494722 82226
rect 494778 82170 494848 82226
rect 494528 82102 494848 82170
rect 494528 82046 494598 82102
rect 494654 82046 494722 82102
rect 494778 82046 494848 82102
rect 494528 81978 494848 82046
rect 494528 81922 494598 81978
rect 494654 81922 494722 81978
rect 494778 81922 494848 81978
rect 494528 81888 494848 81922
rect 525248 82350 525568 82384
rect 525248 82294 525318 82350
rect 525374 82294 525442 82350
rect 525498 82294 525568 82350
rect 525248 82226 525568 82294
rect 525248 82170 525318 82226
rect 525374 82170 525442 82226
rect 525498 82170 525568 82226
rect 525248 82102 525568 82170
rect 525248 82046 525318 82102
rect 525374 82046 525442 82102
rect 525498 82046 525568 82102
rect 525248 81978 525568 82046
rect 525248 81922 525318 81978
rect 525374 81922 525442 81978
rect 525498 81922 525568 81978
rect 525248 81888 525568 81922
rect 555968 82350 556288 82384
rect 555968 82294 556038 82350
rect 556094 82294 556162 82350
rect 556218 82294 556288 82350
rect 555968 82226 556288 82294
rect 555968 82170 556038 82226
rect 556094 82170 556162 82226
rect 556218 82170 556288 82226
rect 555968 82102 556288 82170
rect 555968 82046 556038 82102
rect 556094 82046 556162 82102
rect 556218 82046 556288 82102
rect 555968 81978 556288 82046
rect 555968 81922 556038 81978
rect 556094 81922 556162 81978
rect 556218 81922 556288 81978
rect 555968 81888 556288 81922
rect 443212 80758 443268 80768
rect 443212 20692 443268 80702
rect 448448 76350 448768 76384
rect 448448 76294 448518 76350
rect 448574 76294 448642 76350
rect 448698 76294 448768 76350
rect 448448 76226 448768 76294
rect 448448 76170 448518 76226
rect 448574 76170 448642 76226
rect 448698 76170 448768 76226
rect 448448 76102 448768 76170
rect 448448 76046 448518 76102
rect 448574 76046 448642 76102
rect 448698 76046 448768 76102
rect 448448 75978 448768 76046
rect 448448 75922 448518 75978
rect 448574 75922 448642 75978
rect 448698 75922 448768 75978
rect 448448 75888 448768 75922
rect 479168 76350 479488 76384
rect 479168 76294 479238 76350
rect 479294 76294 479362 76350
rect 479418 76294 479488 76350
rect 479168 76226 479488 76294
rect 479168 76170 479238 76226
rect 479294 76170 479362 76226
rect 479418 76170 479488 76226
rect 479168 76102 479488 76170
rect 479168 76046 479238 76102
rect 479294 76046 479362 76102
rect 479418 76046 479488 76102
rect 479168 75978 479488 76046
rect 479168 75922 479238 75978
rect 479294 75922 479362 75978
rect 479418 75922 479488 75978
rect 479168 75888 479488 75922
rect 509888 76350 510208 76384
rect 509888 76294 509958 76350
rect 510014 76294 510082 76350
rect 510138 76294 510208 76350
rect 509888 76226 510208 76294
rect 509888 76170 509958 76226
rect 510014 76170 510082 76226
rect 510138 76170 510208 76226
rect 509888 76102 510208 76170
rect 509888 76046 509958 76102
rect 510014 76046 510082 76102
rect 510138 76046 510208 76102
rect 509888 75978 510208 76046
rect 509888 75922 509958 75978
rect 510014 75922 510082 75978
rect 510138 75922 510208 75978
rect 509888 75888 510208 75922
rect 540608 76350 540928 76384
rect 540608 76294 540678 76350
rect 540734 76294 540802 76350
rect 540858 76294 540928 76350
rect 540608 76226 540928 76294
rect 540608 76170 540678 76226
rect 540734 76170 540802 76226
rect 540858 76170 540928 76226
rect 540608 76102 540928 76170
rect 540608 76046 540678 76102
rect 540734 76046 540802 76102
rect 540858 76046 540928 76102
rect 540608 75978 540928 76046
rect 540608 75922 540678 75978
rect 540734 75922 540802 75978
rect 540858 75922 540928 75978
rect 540608 75888 540928 75922
rect 571328 76350 571648 76384
rect 571328 76294 571398 76350
rect 571454 76294 571522 76350
rect 571578 76294 571648 76350
rect 571328 76226 571648 76294
rect 571328 76170 571398 76226
rect 571454 76170 571522 76226
rect 571578 76170 571648 76226
rect 571328 76102 571648 76170
rect 571328 76046 571398 76102
rect 571454 76046 571522 76102
rect 571578 76046 571648 76102
rect 571328 75978 571648 76046
rect 571328 75922 571398 75978
rect 571454 75922 571522 75978
rect 571578 75922 571648 75978
rect 571328 75888 571648 75922
rect 463808 64350 464128 64384
rect 463808 64294 463878 64350
rect 463934 64294 464002 64350
rect 464058 64294 464128 64350
rect 463808 64226 464128 64294
rect 463808 64170 463878 64226
rect 463934 64170 464002 64226
rect 464058 64170 464128 64226
rect 463808 64102 464128 64170
rect 463808 64046 463878 64102
rect 463934 64046 464002 64102
rect 464058 64046 464128 64102
rect 463808 63978 464128 64046
rect 463808 63922 463878 63978
rect 463934 63922 464002 63978
rect 464058 63922 464128 63978
rect 463808 63888 464128 63922
rect 494528 64350 494848 64384
rect 494528 64294 494598 64350
rect 494654 64294 494722 64350
rect 494778 64294 494848 64350
rect 494528 64226 494848 64294
rect 494528 64170 494598 64226
rect 494654 64170 494722 64226
rect 494778 64170 494848 64226
rect 494528 64102 494848 64170
rect 494528 64046 494598 64102
rect 494654 64046 494722 64102
rect 494778 64046 494848 64102
rect 494528 63978 494848 64046
rect 494528 63922 494598 63978
rect 494654 63922 494722 63978
rect 494778 63922 494848 63978
rect 494528 63888 494848 63922
rect 525248 64350 525568 64384
rect 525248 64294 525318 64350
rect 525374 64294 525442 64350
rect 525498 64294 525568 64350
rect 525248 64226 525568 64294
rect 525248 64170 525318 64226
rect 525374 64170 525442 64226
rect 525498 64170 525568 64226
rect 525248 64102 525568 64170
rect 525248 64046 525318 64102
rect 525374 64046 525442 64102
rect 525498 64046 525568 64102
rect 525248 63978 525568 64046
rect 525248 63922 525318 63978
rect 525374 63922 525442 63978
rect 525498 63922 525568 63978
rect 525248 63888 525568 63922
rect 555968 64350 556288 64384
rect 555968 64294 556038 64350
rect 556094 64294 556162 64350
rect 556218 64294 556288 64350
rect 555968 64226 556288 64294
rect 555968 64170 556038 64226
rect 556094 64170 556162 64226
rect 556218 64170 556288 64226
rect 555968 64102 556288 64170
rect 555968 64046 556038 64102
rect 556094 64046 556162 64102
rect 556218 64046 556288 64102
rect 555968 63978 556288 64046
rect 555968 63922 556038 63978
rect 556094 63922 556162 63978
rect 556218 63922 556288 63978
rect 555968 63888 556288 63922
rect 448448 58350 448768 58384
rect 448448 58294 448518 58350
rect 448574 58294 448642 58350
rect 448698 58294 448768 58350
rect 448448 58226 448768 58294
rect 448448 58170 448518 58226
rect 448574 58170 448642 58226
rect 448698 58170 448768 58226
rect 448448 58102 448768 58170
rect 448448 58046 448518 58102
rect 448574 58046 448642 58102
rect 448698 58046 448768 58102
rect 448448 57978 448768 58046
rect 448448 57922 448518 57978
rect 448574 57922 448642 57978
rect 448698 57922 448768 57978
rect 448448 57888 448768 57922
rect 479168 58350 479488 58384
rect 479168 58294 479238 58350
rect 479294 58294 479362 58350
rect 479418 58294 479488 58350
rect 479168 58226 479488 58294
rect 479168 58170 479238 58226
rect 479294 58170 479362 58226
rect 479418 58170 479488 58226
rect 479168 58102 479488 58170
rect 479168 58046 479238 58102
rect 479294 58046 479362 58102
rect 479418 58046 479488 58102
rect 479168 57978 479488 58046
rect 479168 57922 479238 57978
rect 479294 57922 479362 57978
rect 479418 57922 479488 57978
rect 479168 57888 479488 57922
rect 509888 58350 510208 58384
rect 509888 58294 509958 58350
rect 510014 58294 510082 58350
rect 510138 58294 510208 58350
rect 509888 58226 510208 58294
rect 509888 58170 509958 58226
rect 510014 58170 510082 58226
rect 510138 58170 510208 58226
rect 509888 58102 510208 58170
rect 509888 58046 509958 58102
rect 510014 58046 510082 58102
rect 510138 58046 510208 58102
rect 509888 57978 510208 58046
rect 509888 57922 509958 57978
rect 510014 57922 510082 57978
rect 510138 57922 510208 57978
rect 509888 57888 510208 57922
rect 540608 58350 540928 58384
rect 540608 58294 540678 58350
rect 540734 58294 540802 58350
rect 540858 58294 540928 58350
rect 540608 58226 540928 58294
rect 540608 58170 540678 58226
rect 540734 58170 540802 58226
rect 540858 58170 540928 58226
rect 540608 58102 540928 58170
rect 540608 58046 540678 58102
rect 540734 58046 540802 58102
rect 540858 58046 540928 58102
rect 540608 57978 540928 58046
rect 540608 57922 540678 57978
rect 540734 57922 540802 57978
rect 540858 57922 540928 57978
rect 540608 57888 540928 57922
rect 571328 58350 571648 58384
rect 571328 58294 571398 58350
rect 571454 58294 571522 58350
rect 571578 58294 571648 58350
rect 571328 58226 571648 58294
rect 571328 58170 571398 58226
rect 571454 58170 571522 58226
rect 571578 58170 571648 58226
rect 571328 58102 571648 58170
rect 571328 58046 571398 58102
rect 571454 58046 571522 58102
rect 571578 58046 571648 58102
rect 571328 57978 571648 58046
rect 571328 57922 571398 57978
rect 571454 57922 571522 57978
rect 571578 57922 571648 57978
rect 571328 57888 571648 57922
rect 463808 46350 464128 46384
rect 463808 46294 463878 46350
rect 463934 46294 464002 46350
rect 464058 46294 464128 46350
rect 463808 46226 464128 46294
rect 463808 46170 463878 46226
rect 463934 46170 464002 46226
rect 464058 46170 464128 46226
rect 463808 46102 464128 46170
rect 463808 46046 463878 46102
rect 463934 46046 464002 46102
rect 464058 46046 464128 46102
rect 463808 45978 464128 46046
rect 463808 45922 463878 45978
rect 463934 45922 464002 45978
rect 464058 45922 464128 45978
rect 463808 45888 464128 45922
rect 494528 46350 494848 46384
rect 494528 46294 494598 46350
rect 494654 46294 494722 46350
rect 494778 46294 494848 46350
rect 494528 46226 494848 46294
rect 494528 46170 494598 46226
rect 494654 46170 494722 46226
rect 494778 46170 494848 46226
rect 494528 46102 494848 46170
rect 494528 46046 494598 46102
rect 494654 46046 494722 46102
rect 494778 46046 494848 46102
rect 494528 45978 494848 46046
rect 494528 45922 494598 45978
rect 494654 45922 494722 45978
rect 494778 45922 494848 45978
rect 494528 45888 494848 45922
rect 525248 46350 525568 46384
rect 525248 46294 525318 46350
rect 525374 46294 525442 46350
rect 525498 46294 525568 46350
rect 525248 46226 525568 46294
rect 525248 46170 525318 46226
rect 525374 46170 525442 46226
rect 525498 46170 525568 46226
rect 525248 46102 525568 46170
rect 525248 46046 525318 46102
rect 525374 46046 525442 46102
rect 525498 46046 525568 46102
rect 525248 45978 525568 46046
rect 525248 45922 525318 45978
rect 525374 45922 525442 45978
rect 525498 45922 525568 45978
rect 525248 45888 525568 45922
rect 555968 46350 556288 46384
rect 555968 46294 556038 46350
rect 556094 46294 556162 46350
rect 556218 46294 556288 46350
rect 555968 46226 556288 46294
rect 555968 46170 556038 46226
rect 556094 46170 556162 46226
rect 556218 46170 556288 46226
rect 555968 46102 556288 46170
rect 555968 46046 556038 46102
rect 556094 46046 556162 46102
rect 556218 46046 556288 46102
rect 555968 45978 556288 46046
rect 555968 45922 556038 45978
rect 556094 45922 556162 45978
rect 556218 45922 556288 45978
rect 555968 45888 556288 45922
rect 448448 40350 448768 40384
rect 448448 40294 448518 40350
rect 448574 40294 448642 40350
rect 448698 40294 448768 40350
rect 448448 40226 448768 40294
rect 448448 40170 448518 40226
rect 448574 40170 448642 40226
rect 448698 40170 448768 40226
rect 448448 40102 448768 40170
rect 448448 40046 448518 40102
rect 448574 40046 448642 40102
rect 448698 40046 448768 40102
rect 448448 39978 448768 40046
rect 448448 39922 448518 39978
rect 448574 39922 448642 39978
rect 448698 39922 448768 39978
rect 448448 39888 448768 39922
rect 479168 40350 479488 40384
rect 479168 40294 479238 40350
rect 479294 40294 479362 40350
rect 479418 40294 479488 40350
rect 479168 40226 479488 40294
rect 479168 40170 479238 40226
rect 479294 40170 479362 40226
rect 479418 40170 479488 40226
rect 479168 40102 479488 40170
rect 479168 40046 479238 40102
rect 479294 40046 479362 40102
rect 479418 40046 479488 40102
rect 479168 39978 479488 40046
rect 479168 39922 479238 39978
rect 479294 39922 479362 39978
rect 479418 39922 479488 39978
rect 479168 39888 479488 39922
rect 509888 40350 510208 40384
rect 509888 40294 509958 40350
rect 510014 40294 510082 40350
rect 510138 40294 510208 40350
rect 509888 40226 510208 40294
rect 509888 40170 509958 40226
rect 510014 40170 510082 40226
rect 510138 40170 510208 40226
rect 509888 40102 510208 40170
rect 509888 40046 509958 40102
rect 510014 40046 510082 40102
rect 510138 40046 510208 40102
rect 509888 39978 510208 40046
rect 509888 39922 509958 39978
rect 510014 39922 510082 39978
rect 510138 39922 510208 39978
rect 509888 39888 510208 39922
rect 540608 40350 540928 40384
rect 540608 40294 540678 40350
rect 540734 40294 540802 40350
rect 540858 40294 540928 40350
rect 540608 40226 540928 40294
rect 540608 40170 540678 40226
rect 540734 40170 540802 40226
rect 540858 40170 540928 40226
rect 540608 40102 540928 40170
rect 540608 40046 540678 40102
rect 540734 40046 540802 40102
rect 540858 40046 540928 40102
rect 540608 39978 540928 40046
rect 540608 39922 540678 39978
rect 540734 39922 540802 39978
rect 540858 39922 540928 39978
rect 540608 39888 540928 39922
rect 571328 40350 571648 40384
rect 571328 40294 571398 40350
rect 571454 40294 571522 40350
rect 571578 40294 571648 40350
rect 571328 40226 571648 40294
rect 571328 40170 571398 40226
rect 571454 40170 571522 40226
rect 571578 40170 571648 40226
rect 571328 40102 571648 40170
rect 571328 40046 571398 40102
rect 571454 40046 571522 40102
rect 571578 40046 571648 40102
rect 571328 39978 571648 40046
rect 571328 39922 571398 39978
rect 571454 39922 571522 39978
rect 571578 39922 571648 39978
rect 571328 39888 571648 39922
rect 463808 28350 464128 28384
rect 463808 28294 463878 28350
rect 463934 28294 464002 28350
rect 464058 28294 464128 28350
rect 463808 28226 464128 28294
rect 463808 28170 463878 28226
rect 463934 28170 464002 28226
rect 464058 28170 464128 28226
rect 463808 28102 464128 28170
rect 463808 28046 463878 28102
rect 463934 28046 464002 28102
rect 464058 28046 464128 28102
rect 463808 27978 464128 28046
rect 463808 27922 463878 27978
rect 463934 27922 464002 27978
rect 464058 27922 464128 27978
rect 463808 27888 464128 27922
rect 494528 28350 494848 28384
rect 494528 28294 494598 28350
rect 494654 28294 494722 28350
rect 494778 28294 494848 28350
rect 494528 28226 494848 28294
rect 494528 28170 494598 28226
rect 494654 28170 494722 28226
rect 494778 28170 494848 28226
rect 494528 28102 494848 28170
rect 494528 28046 494598 28102
rect 494654 28046 494722 28102
rect 494778 28046 494848 28102
rect 494528 27978 494848 28046
rect 494528 27922 494598 27978
rect 494654 27922 494722 27978
rect 494778 27922 494848 27978
rect 494528 27888 494848 27922
rect 525248 28350 525568 28384
rect 525248 28294 525318 28350
rect 525374 28294 525442 28350
rect 525498 28294 525568 28350
rect 525248 28226 525568 28294
rect 525248 28170 525318 28226
rect 525374 28170 525442 28226
rect 525498 28170 525568 28226
rect 525248 28102 525568 28170
rect 525248 28046 525318 28102
rect 525374 28046 525442 28102
rect 525498 28046 525568 28102
rect 525248 27978 525568 28046
rect 525248 27922 525318 27978
rect 525374 27922 525442 27978
rect 525498 27922 525568 27978
rect 525248 27888 525568 27922
rect 555968 28350 556288 28384
rect 555968 28294 556038 28350
rect 556094 28294 556162 28350
rect 556218 28294 556288 28350
rect 555968 28226 556288 28294
rect 555968 28170 556038 28226
rect 556094 28170 556162 28226
rect 556218 28170 556288 28226
rect 555968 28102 556288 28170
rect 555968 28046 556038 28102
rect 556094 28046 556162 28102
rect 556218 28046 556288 28102
rect 555968 27978 556288 28046
rect 555968 27922 556038 27978
rect 556094 27922 556162 27978
rect 556218 27922 556288 27978
rect 555968 27888 556288 27922
rect 443212 20626 443268 20636
rect 587132 20098 587188 258188
rect 587132 20032 587188 20042
rect 589098 256350 589718 273922
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 589098 58350 589718 75922
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 443100 16146 443156 16156
rect 442988 4722 443044 4732
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 4350 466838 19026
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 10350 470558 19026
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 479724 8038 479780 8048
rect 479724 4116 479780 7982
rect 479724 4050 479780 4060
rect 496938 4350 497558 19026
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 475916 2818 475972 2828
rect 475916 1764 475972 2762
rect 475916 1698 475972 1708
rect 474012 838 474068 848
rect 474012 644 474068 782
rect 474012 578 474068 588
rect 485548 658 485604 682
rect 485548 578 485604 588
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 10350 501278 19026
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 500658 -1120 501278 9922
rect 523516 8578 523572 8588
rect 506380 6418 506436 6428
rect 506380 3444 506436 6362
rect 506380 3378 506436 3388
rect 512092 6238 512148 6248
rect 512092 3444 512148 6182
rect 512092 3378 512148 3388
rect 517804 6058 517860 6068
rect 517804 3444 517860 6002
rect 523516 4340 523572 8522
rect 523516 4274 523572 4284
rect 527658 4350 528278 19026
rect 531378 10350 531998 19026
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 517804 3378 517860 3388
rect 527658 4226 528278 4294
rect 531132 9478 531188 9488
rect 531132 4340 531188 9422
rect 531132 4274 531188 4284
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 515900 3178 515956 3188
rect 515900 1764 515956 3122
rect 515900 1698 515956 1708
rect 527324 644 527380 654
rect 527324 298 527380 588
rect 527324 232 527380 242
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 -1120 531998 9922
rect 540652 7858 540708 7868
rect 534940 5878 534996 5888
rect 534940 3444 534996 5822
rect 540652 4004 540708 7802
rect 540652 3938 540708 3948
rect 546364 7678 546420 7688
rect 546364 3892 546420 7622
rect 546364 3826 546420 3836
rect 557788 7498 557844 7508
rect 557788 3780 557844 7442
rect 557788 3714 557844 3724
rect 558378 4350 558998 19026
rect 562098 10350 562718 19026
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 534940 3378 534996 3388
rect 552636 3444 552692 3454
rect 552636 3358 552692 3388
rect 552636 3292 552692 3302
rect 542668 2998 542724 3008
rect 542668 1764 542724 2942
rect 542668 1698 542724 1708
rect 533036 644 533092 654
rect 533036 118 533092 588
rect 553980 644 554036 654
rect 553980 478 554036 588
rect 553980 412 554036 422
rect 533036 52 533092 62
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 -160 558998 3922
rect 559692 4798 559748 4808
rect 559692 3444 559748 4742
rect 559692 3378 559748 3388
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 -1120 562718 9922
rect 581308 15958 581364 15968
rect 571228 9298 571284 9308
rect 571228 6804 571284 9242
rect 571228 6738 571284 6748
rect 571228 4978 571284 4988
rect 571228 3444 571284 4922
rect 581308 4228 581364 15902
rect 581308 4162 581364 4172
rect 589098 4350 589718 21922
rect 590492 245028 590548 245038
rect 590492 19348 590548 244972
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 590716 231924 590772 231934
rect 590604 205380 590660 205390
rect 590604 20804 590660 205324
rect 590604 20738 590660 20748
rect 590716 19796 590772 231868
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 590716 19730 590772 19740
rect 590828 192164 590884 192174
rect 590492 19282 590548 19292
rect 590828 18340 590884 192108
rect 590828 18274 590884 18284
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 571228 3378 571284 3388
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 22518 562294 22574 562350
rect 22642 562294 22698 562350
rect 22518 562170 22574 562226
rect 22642 562170 22698 562226
rect 22518 562046 22574 562102
rect 22642 562046 22698 562102
rect 22518 561922 22574 561978
rect 22642 561922 22698 561978
rect 22518 544294 22574 544350
rect 22642 544294 22698 544350
rect 22518 544170 22574 544226
rect 22642 544170 22698 544226
rect 22518 544046 22574 544102
rect 22642 544046 22698 544102
rect 22518 543922 22574 543978
rect 22642 543922 22698 543978
rect 22518 526294 22574 526350
rect 22642 526294 22698 526350
rect 22518 526170 22574 526226
rect 22642 526170 22698 526226
rect 22518 526046 22574 526102
rect 22642 526046 22698 526102
rect 22518 525922 22574 525978
rect 22642 525922 22698 525978
rect 22518 508294 22574 508350
rect 22642 508294 22698 508350
rect 22518 508170 22574 508226
rect 22642 508170 22698 508226
rect 22518 508046 22574 508102
rect 22642 508046 22698 508102
rect 22518 507922 22574 507978
rect 22642 507922 22698 507978
rect 22518 490294 22574 490350
rect 22642 490294 22698 490350
rect 22518 490170 22574 490226
rect 22642 490170 22698 490226
rect 22518 490046 22574 490102
rect 22642 490046 22698 490102
rect 22518 489922 22574 489978
rect 22642 489922 22698 489978
rect 22518 472294 22574 472350
rect 22642 472294 22698 472350
rect 22518 472170 22574 472226
rect 22642 472170 22698 472226
rect 22518 472046 22574 472102
rect 22642 472046 22698 472102
rect 22518 471922 22574 471978
rect 22642 471922 22698 471978
rect 22518 454294 22574 454350
rect 22642 454294 22698 454350
rect 22518 454170 22574 454226
rect 22642 454170 22698 454226
rect 22518 454046 22574 454102
rect 22642 454046 22698 454102
rect 22518 453922 22574 453978
rect 22642 453922 22698 453978
rect 22518 436294 22574 436350
rect 22642 436294 22698 436350
rect 22518 436170 22574 436226
rect 22642 436170 22698 436226
rect 22518 436046 22574 436102
rect 22642 436046 22698 436102
rect 22518 435922 22574 435978
rect 22642 435922 22698 435978
rect 22518 418294 22574 418350
rect 22642 418294 22698 418350
rect 22518 418170 22574 418226
rect 22642 418170 22698 418226
rect 22518 418046 22574 418102
rect 22642 418046 22698 418102
rect 22518 417922 22574 417978
rect 22642 417922 22698 417978
rect 22518 400294 22574 400350
rect 22642 400294 22698 400350
rect 22518 400170 22574 400226
rect 22642 400170 22698 400226
rect 22518 400046 22574 400102
rect 22642 400046 22698 400102
rect 22518 399922 22574 399978
rect 22642 399922 22698 399978
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 37878 568294 37934 568350
rect 38002 568294 38058 568350
rect 37878 568170 37934 568226
rect 38002 568170 38058 568226
rect 37878 568046 37934 568102
rect 38002 568046 38058 568102
rect 37878 567922 37934 567978
rect 38002 567922 38058 567978
rect 68598 568294 68654 568350
rect 68722 568294 68778 568350
rect 68598 568170 68654 568226
rect 68722 568170 68778 568226
rect 68598 568046 68654 568102
rect 68722 568046 68778 568102
rect 68598 567922 68654 567978
rect 68722 567922 68778 567978
rect 99318 568294 99374 568350
rect 99442 568294 99498 568350
rect 99318 568170 99374 568226
rect 99442 568170 99498 568226
rect 99318 568046 99374 568102
rect 99442 568046 99498 568102
rect 99318 567922 99374 567978
rect 99442 567922 99498 567978
rect 130038 568294 130094 568350
rect 130162 568294 130218 568350
rect 130038 568170 130094 568226
rect 130162 568170 130218 568226
rect 130038 568046 130094 568102
rect 130162 568046 130218 568102
rect 130038 567922 130094 567978
rect 130162 567922 130218 567978
rect 160758 568294 160814 568350
rect 160882 568294 160938 568350
rect 160758 568170 160814 568226
rect 160882 568170 160938 568226
rect 160758 568046 160814 568102
rect 160882 568046 160938 568102
rect 160758 567922 160814 567978
rect 160882 567922 160938 567978
rect 191478 568294 191534 568350
rect 191602 568294 191658 568350
rect 191478 568170 191534 568226
rect 191602 568170 191658 568226
rect 191478 568046 191534 568102
rect 191602 568046 191658 568102
rect 191478 567922 191534 567978
rect 191602 567922 191658 567978
rect 222198 568294 222254 568350
rect 222322 568294 222378 568350
rect 222198 568170 222254 568226
rect 222322 568170 222378 568226
rect 222198 568046 222254 568102
rect 222322 568046 222378 568102
rect 222198 567922 222254 567978
rect 222322 567922 222378 567978
rect 252918 568294 252974 568350
rect 253042 568294 253098 568350
rect 252918 568170 252974 568226
rect 253042 568170 253098 568226
rect 252918 568046 252974 568102
rect 253042 568046 253098 568102
rect 252918 567922 252974 567978
rect 253042 567922 253098 567978
rect 283638 568294 283694 568350
rect 283762 568294 283818 568350
rect 283638 568170 283694 568226
rect 283762 568170 283818 568226
rect 283638 568046 283694 568102
rect 283762 568046 283818 568102
rect 283638 567922 283694 567978
rect 283762 567922 283818 567978
rect 314358 568294 314414 568350
rect 314482 568294 314538 568350
rect 314358 568170 314414 568226
rect 314482 568170 314538 568226
rect 314358 568046 314414 568102
rect 314482 568046 314538 568102
rect 314358 567922 314414 567978
rect 314482 567922 314538 567978
rect 345078 568294 345134 568350
rect 345202 568294 345258 568350
rect 345078 568170 345134 568226
rect 345202 568170 345258 568226
rect 345078 568046 345134 568102
rect 345202 568046 345258 568102
rect 345078 567922 345134 567978
rect 345202 567922 345258 567978
rect 375798 568294 375854 568350
rect 375922 568294 375978 568350
rect 375798 568170 375854 568226
rect 375922 568170 375978 568226
rect 375798 568046 375854 568102
rect 375922 568046 375978 568102
rect 375798 567922 375854 567978
rect 375922 567922 375978 567978
rect 406518 568294 406574 568350
rect 406642 568294 406698 568350
rect 406518 568170 406574 568226
rect 406642 568170 406698 568226
rect 406518 568046 406574 568102
rect 406642 568046 406698 568102
rect 406518 567922 406574 567978
rect 406642 567922 406698 567978
rect 437238 568294 437294 568350
rect 437362 568294 437418 568350
rect 437238 568170 437294 568226
rect 437362 568170 437418 568226
rect 437238 568046 437294 568102
rect 437362 568046 437418 568102
rect 437238 567922 437294 567978
rect 437362 567922 437418 567978
rect 467958 568294 468014 568350
rect 468082 568294 468138 568350
rect 467958 568170 468014 568226
rect 468082 568170 468138 568226
rect 467958 568046 468014 568102
rect 468082 568046 468138 568102
rect 467958 567922 468014 567978
rect 468082 567922 468138 567978
rect 498678 568294 498734 568350
rect 498802 568294 498858 568350
rect 498678 568170 498734 568226
rect 498802 568170 498858 568226
rect 498678 568046 498734 568102
rect 498802 568046 498858 568102
rect 498678 567922 498734 567978
rect 498802 567922 498858 567978
rect 529398 568294 529454 568350
rect 529522 568294 529578 568350
rect 529398 568170 529454 568226
rect 529522 568170 529578 568226
rect 529398 568046 529454 568102
rect 529522 568046 529578 568102
rect 529398 567922 529454 567978
rect 529522 567922 529578 567978
rect 53238 562294 53294 562350
rect 53362 562294 53418 562350
rect 53238 562170 53294 562226
rect 53362 562170 53418 562226
rect 53238 562046 53294 562102
rect 53362 562046 53418 562102
rect 53238 561922 53294 561978
rect 53362 561922 53418 561978
rect 83958 562294 84014 562350
rect 84082 562294 84138 562350
rect 83958 562170 84014 562226
rect 84082 562170 84138 562226
rect 83958 562046 84014 562102
rect 84082 562046 84138 562102
rect 83958 561922 84014 561978
rect 84082 561922 84138 561978
rect 114678 562294 114734 562350
rect 114802 562294 114858 562350
rect 114678 562170 114734 562226
rect 114802 562170 114858 562226
rect 114678 562046 114734 562102
rect 114802 562046 114858 562102
rect 114678 561922 114734 561978
rect 114802 561922 114858 561978
rect 145398 562294 145454 562350
rect 145522 562294 145578 562350
rect 145398 562170 145454 562226
rect 145522 562170 145578 562226
rect 145398 562046 145454 562102
rect 145522 562046 145578 562102
rect 145398 561922 145454 561978
rect 145522 561922 145578 561978
rect 176118 562294 176174 562350
rect 176242 562294 176298 562350
rect 176118 562170 176174 562226
rect 176242 562170 176298 562226
rect 176118 562046 176174 562102
rect 176242 562046 176298 562102
rect 176118 561922 176174 561978
rect 176242 561922 176298 561978
rect 206838 562294 206894 562350
rect 206962 562294 207018 562350
rect 206838 562170 206894 562226
rect 206962 562170 207018 562226
rect 206838 562046 206894 562102
rect 206962 562046 207018 562102
rect 206838 561922 206894 561978
rect 206962 561922 207018 561978
rect 237558 562294 237614 562350
rect 237682 562294 237738 562350
rect 237558 562170 237614 562226
rect 237682 562170 237738 562226
rect 237558 562046 237614 562102
rect 237682 562046 237738 562102
rect 237558 561922 237614 561978
rect 237682 561922 237738 561978
rect 268278 562294 268334 562350
rect 268402 562294 268458 562350
rect 268278 562170 268334 562226
rect 268402 562170 268458 562226
rect 268278 562046 268334 562102
rect 268402 562046 268458 562102
rect 268278 561922 268334 561978
rect 268402 561922 268458 561978
rect 298998 562294 299054 562350
rect 299122 562294 299178 562350
rect 298998 562170 299054 562226
rect 299122 562170 299178 562226
rect 298998 562046 299054 562102
rect 299122 562046 299178 562102
rect 298998 561922 299054 561978
rect 299122 561922 299178 561978
rect 329718 562294 329774 562350
rect 329842 562294 329898 562350
rect 329718 562170 329774 562226
rect 329842 562170 329898 562226
rect 329718 562046 329774 562102
rect 329842 562046 329898 562102
rect 329718 561922 329774 561978
rect 329842 561922 329898 561978
rect 360438 562294 360494 562350
rect 360562 562294 360618 562350
rect 360438 562170 360494 562226
rect 360562 562170 360618 562226
rect 360438 562046 360494 562102
rect 360562 562046 360618 562102
rect 360438 561922 360494 561978
rect 360562 561922 360618 561978
rect 391158 562294 391214 562350
rect 391282 562294 391338 562350
rect 391158 562170 391214 562226
rect 391282 562170 391338 562226
rect 391158 562046 391214 562102
rect 391282 562046 391338 562102
rect 391158 561922 391214 561978
rect 391282 561922 391338 561978
rect 421878 562294 421934 562350
rect 422002 562294 422058 562350
rect 421878 562170 421934 562226
rect 422002 562170 422058 562226
rect 421878 562046 421934 562102
rect 422002 562046 422058 562102
rect 421878 561922 421934 561978
rect 422002 561922 422058 561978
rect 452598 562294 452654 562350
rect 452722 562294 452778 562350
rect 452598 562170 452654 562226
rect 452722 562170 452778 562226
rect 452598 562046 452654 562102
rect 452722 562046 452778 562102
rect 452598 561922 452654 561978
rect 452722 561922 452778 561978
rect 483318 562294 483374 562350
rect 483442 562294 483498 562350
rect 483318 562170 483374 562226
rect 483442 562170 483498 562226
rect 483318 562046 483374 562102
rect 483442 562046 483498 562102
rect 483318 561922 483374 561978
rect 483442 561922 483498 561978
rect 514038 562294 514094 562350
rect 514162 562294 514218 562350
rect 514038 562170 514094 562226
rect 514162 562170 514218 562226
rect 514038 562046 514094 562102
rect 514162 562046 514218 562102
rect 514038 561922 514094 561978
rect 514162 561922 514218 561978
rect 544758 562294 544814 562350
rect 544882 562294 544938 562350
rect 544758 562170 544814 562226
rect 544882 562170 544938 562226
rect 544758 562046 544814 562102
rect 544882 562046 544938 562102
rect 544758 561922 544814 561978
rect 544882 561922 544938 561978
rect 37878 550294 37934 550350
rect 38002 550294 38058 550350
rect 37878 550170 37934 550226
rect 38002 550170 38058 550226
rect 37878 550046 37934 550102
rect 38002 550046 38058 550102
rect 37878 549922 37934 549978
rect 38002 549922 38058 549978
rect 68598 550294 68654 550350
rect 68722 550294 68778 550350
rect 68598 550170 68654 550226
rect 68722 550170 68778 550226
rect 68598 550046 68654 550102
rect 68722 550046 68778 550102
rect 68598 549922 68654 549978
rect 68722 549922 68778 549978
rect 99318 550294 99374 550350
rect 99442 550294 99498 550350
rect 99318 550170 99374 550226
rect 99442 550170 99498 550226
rect 99318 550046 99374 550102
rect 99442 550046 99498 550102
rect 99318 549922 99374 549978
rect 99442 549922 99498 549978
rect 130038 550294 130094 550350
rect 130162 550294 130218 550350
rect 130038 550170 130094 550226
rect 130162 550170 130218 550226
rect 130038 550046 130094 550102
rect 130162 550046 130218 550102
rect 130038 549922 130094 549978
rect 130162 549922 130218 549978
rect 160758 550294 160814 550350
rect 160882 550294 160938 550350
rect 160758 550170 160814 550226
rect 160882 550170 160938 550226
rect 160758 550046 160814 550102
rect 160882 550046 160938 550102
rect 160758 549922 160814 549978
rect 160882 549922 160938 549978
rect 191478 550294 191534 550350
rect 191602 550294 191658 550350
rect 191478 550170 191534 550226
rect 191602 550170 191658 550226
rect 191478 550046 191534 550102
rect 191602 550046 191658 550102
rect 191478 549922 191534 549978
rect 191602 549922 191658 549978
rect 222198 550294 222254 550350
rect 222322 550294 222378 550350
rect 222198 550170 222254 550226
rect 222322 550170 222378 550226
rect 222198 550046 222254 550102
rect 222322 550046 222378 550102
rect 222198 549922 222254 549978
rect 222322 549922 222378 549978
rect 252918 550294 252974 550350
rect 253042 550294 253098 550350
rect 252918 550170 252974 550226
rect 253042 550170 253098 550226
rect 252918 550046 252974 550102
rect 253042 550046 253098 550102
rect 252918 549922 252974 549978
rect 253042 549922 253098 549978
rect 283638 550294 283694 550350
rect 283762 550294 283818 550350
rect 283638 550170 283694 550226
rect 283762 550170 283818 550226
rect 283638 550046 283694 550102
rect 283762 550046 283818 550102
rect 283638 549922 283694 549978
rect 283762 549922 283818 549978
rect 314358 550294 314414 550350
rect 314482 550294 314538 550350
rect 314358 550170 314414 550226
rect 314482 550170 314538 550226
rect 314358 550046 314414 550102
rect 314482 550046 314538 550102
rect 314358 549922 314414 549978
rect 314482 549922 314538 549978
rect 345078 550294 345134 550350
rect 345202 550294 345258 550350
rect 345078 550170 345134 550226
rect 345202 550170 345258 550226
rect 345078 550046 345134 550102
rect 345202 550046 345258 550102
rect 345078 549922 345134 549978
rect 345202 549922 345258 549978
rect 375798 550294 375854 550350
rect 375922 550294 375978 550350
rect 375798 550170 375854 550226
rect 375922 550170 375978 550226
rect 375798 550046 375854 550102
rect 375922 550046 375978 550102
rect 375798 549922 375854 549978
rect 375922 549922 375978 549978
rect 406518 550294 406574 550350
rect 406642 550294 406698 550350
rect 406518 550170 406574 550226
rect 406642 550170 406698 550226
rect 406518 550046 406574 550102
rect 406642 550046 406698 550102
rect 406518 549922 406574 549978
rect 406642 549922 406698 549978
rect 437238 550294 437294 550350
rect 437362 550294 437418 550350
rect 437238 550170 437294 550226
rect 437362 550170 437418 550226
rect 437238 550046 437294 550102
rect 437362 550046 437418 550102
rect 437238 549922 437294 549978
rect 437362 549922 437418 549978
rect 467958 550294 468014 550350
rect 468082 550294 468138 550350
rect 467958 550170 468014 550226
rect 468082 550170 468138 550226
rect 467958 550046 468014 550102
rect 468082 550046 468138 550102
rect 467958 549922 468014 549978
rect 468082 549922 468138 549978
rect 498678 550294 498734 550350
rect 498802 550294 498858 550350
rect 498678 550170 498734 550226
rect 498802 550170 498858 550226
rect 498678 550046 498734 550102
rect 498802 550046 498858 550102
rect 498678 549922 498734 549978
rect 498802 549922 498858 549978
rect 529398 550294 529454 550350
rect 529522 550294 529578 550350
rect 529398 550170 529454 550226
rect 529522 550170 529578 550226
rect 529398 550046 529454 550102
rect 529522 550046 529578 550102
rect 529398 549922 529454 549978
rect 529522 549922 529578 549978
rect 53238 544294 53294 544350
rect 53362 544294 53418 544350
rect 53238 544170 53294 544226
rect 53362 544170 53418 544226
rect 53238 544046 53294 544102
rect 53362 544046 53418 544102
rect 53238 543922 53294 543978
rect 53362 543922 53418 543978
rect 83958 544294 84014 544350
rect 84082 544294 84138 544350
rect 83958 544170 84014 544226
rect 84082 544170 84138 544226
rect 83958 544046 84014 544102
rect 84082 544046 84138 544102
rect 83958 543922 84014 543978
rect 84082 543922 84138 543978
rect 114678 544294 114734 544350
rect 114802 544294 114858 544350
rect 114678 544170 114734 544226
rect 114802 544170 114858 544226
rect 114678 544046 114734 544102
rect 114802 544046 114858 544102
rect 114678 543922 114734 543978
rect 114802 543922 114858 543978
rect 145398 544294 145454 544350
rect 145522 544294 145578 544350
rect 145398 544170 145454 544226
rect 145522 544170 145578 544226
rect 145398 544046 145454 544102
rect 145522 544046 145578 544102
rect 145398 543922 145454 543978
rect 145522 543922 145578 543978
rect 176118 544294 176174 544350
rect 176242 544294 176298 544350
rect 176118 544170 176174 544226
rect 176242 544170 176298 544226
rect 176118 544046 176174 544102
rect 176242 544046 176298 544102
rect 176118 543922 176174 543978
rect 176242 543922 176298 543978
rect 206838 544294 206894 544350
rect 206962 544294 207018 544350
rect 206838 544170 206894 544226
rect 206962 544170 207018 544226
rect 206838 544046 206894 544102
rect 206962 544046 207018 544102
rect 206838 543922 206894 543978
rect 206962 543922 207018 543978
rect 237558 544294 237614 544350
rect 237682 544294 237738 544350
rect 237558 544170 237614 544226
rect 237682 544170 237738 544226
rect 237558 544046 237614 544102
rect 237682 544046 237738 544102
rect 237558 543922 237614 543978
rect 237682 543922 237738 543978
rect 268278 544294 268334 544350
rect 268402 544294 268458 544350
rect 268278 544170 268334 544226
rect 268402 544170 268458 544226
rect 268278 544046 268334 544102
rect 268402 544046 268458 544102
rect 268278 543922 268334 543978
rect 268402 543922 268458 543978
rect 298998 544294 299054 544350
rect 299122 544294 299178 544350
rect 298998 544170 299054 544226
rect 299122 544170 299178 544226
rect 298998 544046 299054 544102
rect 299122 544046 299178 544102
rect 298998 543922 299054 543978
rect 299122 543922 299178 543978
rect 329718 544294 329774 544350
rect 329842 544294 329898 544350
rect 329718 544170 329774 544226
rect 329842 544170 329898 544226
rect 329718 544046 329774 544102
rect 329842 544046 329898 544102
rect 329718 543922 329774 543978
rect 329842 543922 329898 543978
rect 360438 544294 360494 544350
rect 360562 544294 360618 544350
rect 360438 544170 360494 544226
rect 360562 544170 360618 544226
rect 360438 544046 360494 544102
rect 360562 544046 360618 544102
rect 360438 543922 360494 543978
rect 360562 543922 360618 543978
rect 391158 544294 391214 544350
rect 391282 544294 391338 544350
rect 391158 544170 391214 544226
rect 391282 544170 391338 544226
rect 391158 544046 391214 544102
rect 391282 544046 391338 544102
rect 391158 543922 391214 543978
rect 391282 543922 391338 543978
rect 421878 544294 421934 544350
rect 422002 544294 422058 544350
rect 421878 544170 421934 544226
rect 422002 544170 422058 544226
rect 421878 544046 421934 544102
rect 422002 544046 422058 544102
rect 421878 543922 421934 543978
rect 422002 543922 422058 543978
rect 452598 544294 452654 544350
rect 452722 544294 452778 544350
rect 452598 544170 452654 544226
rect 452722 544170 452778 544226
rect 452598 544046 452654 544102
rect 452722 544046 452778 544102
rect 452598 543922 452654 543978
rect 452722 543922 452778 543978
rect 483318 544294 483374 544350
rect 483442 544294 483498 544350
rect 483318 544170 483374 544226
rect 483442 544170 483498 544226
rect 483318 544046 483374 544102
rect 483442 544046 483498 544102
rect 483318 543922 483374 543978
rect 483442 543922 483498 543978
rect 514038 544294 514094 544350
rect 514162 544294 514218 544350
rect 514038 544170 514094 544226
rect 514162 544170 514218 544226
rect 514038 544046 514094 544102
rect 514162 544046 514218 544102
rect 514038 543922 514094 543978
rect 514162 543922 514218 543978
rect 544758 544294 544814 544350
rect 544882 544294 544938 544350
rect 544758 544170 544814 544226
rect 544882 544170 544938 544226
rect 544758 544046 544814 544102
rect 544882 544046 544938 544102
rect 544758 543922 544814 543978
rect 544882 543922 544938 543978
rect 37878 532294 37934 532350
rect 38002 532294 38058 532350
rect 37878 532170 37934 532226
rect 38002 532170 38058 532226
rect 37878 532046 37934 532102
rect 38002 532046 38058 532102
rect 37878 531922 37934 531978
rect 38002 531922 38058 531978
rect 68598 532294 68654 532350
rect 68722 532294 68778 532350
rect 68598 532170 68654 532226
rect 68722 532170 68778 532226
rect 68598 532046 68654 532102
rect 68722 532046 68778 532102
rect 68598 531922 68654 531978
rect 68722 531922 68778 531978
rect 99318 532294 99374 532350
rect 99442 532294 99498 532350
rect 99318 532170 99374 532226
rect 99442 532170 99498 532226
rect 99318 532046 99374 532102
rect 99442 532046 99498 532102
rect 99318 531922 99374 531978
rect 99442 531922 99498 531978
rect 130038 532294 130094 532350
rect 130162 532294 130218 532350
rect 130038 532170 130094 532226
rect 130162 532170 130218 532226
rect 130038 532046 130094 532102
rect 130162 532046 130218 532102
rect 130038 531922 130094 531978
rect 130162 531922 130218 531978
rect 160758 532294 160814 532350
rect 160882 532294 160938 532350
rect 160758 532170 160814 532226
rect 160882 532170 160938 532226
rect 160758 532046 160814 532102
rect 160882 532046 160938 532102
rect 160758 531922 160814 531978
rect 160882 531922 160938 531978
rect 191478 532294 191534 532350
rect 191602 532294 191658 532350
rect 191478 532170 191534 532226
rect 191602 532170 191658 532226
rect 191478 532046 191534 532102
rect 191602 532046 191658 532102
rect 191478 531922 191534 531978
rect 191602 531922 191658 531978
rect 222198 532294 222254 532350
rect 222322 532294 222378 532350
rect 222198 532170 222254 532226
rect 222322 532170 222378 532226
rect 222198 532046 222254 532102
rect 222322 532046 222378 532102
rect 222198 531922 222254 531978
rect 222322 531922 222378 531978
rect 252918 532294 252974 532350
rect 253042 532294 253098 532350
rect 252918 532170 252974 532226
rect 253042 532170 253098 532226
rect 252918 532046 252974 532102
rect 253042 532046 253098 532102
rect 252918 531922 252974 531978
rect 253042 531922 253098 531978
rect 283638 532294 283694 532350
rect 283762 532294 283818 532350
rect 283638 532170 283694 532226
rect 283762 532170 283818 532226
rect 283638 532046 283694 532102
rect 283762 532046 283818 532102
rect 283638 531922 283694 531978
rect 283762 531922 283818 531978
rect 314358 532294 314414 532350
rect 314482 532294 314538 532350
rect 314358 532170 314414 532226
rect 314482 532170 314538 532226
rect 314358 532046 314414 532102
rect 314482 532046 314538 532102
rect 314358 531922 314414 531978
rect 314482 531922 314538 531978
rect 345078 532294 345134 532350
rect 345202 532294 345258 532350
rect 345078 532170 345134 532226
rect 345202 532170 345258 532226
rect 345078 532046 345134 532102
rect 345202 532046 345258 532102
rect 345078 531922 345134 531978
rect 345202 531922 345258 531978
rect 375798 532294 375854 532350
rect 375922 532294 375978 532350
rect 375798 532170 375854 532226
rect 375922 532170 375978 532226
rect 375798 532046 375854 532102
rect 375922 532046 375978 532102
rect 375798 531922 375854 531978
rect 375922 531922 375978 531978
rect 406518 532294 406574 532350
rect 406642 532294 406698 532350
rect 406518 532170 406574 532226
rect 406642 532170 406698 532226
rect 406518 532046 406574 532102
rect 406642 532046 406698 532102
rect 406518 531922 406574 531978
rect 406642 531922 406698 531978
rect 437238 532294 437294 532350
rect 437362 532294 437418 532350
rect 437238 532170 437294 532226
rect 437362 532170 437418 532226
rect 437238 532046 437294 532102
rect 437362 532046 437418 532102
rect 437238 531922 437294 531978
rect 437362 531922 437418 531978
rect 467958 532294 468014 532350
rect 468082 532294 468138 532350
rect 467958 532170 468014 532226
rect 468082 532170 468138 532226
rect 467958 532046 468014 532102
rect 468082 532046 468138 532102
rect 467958 531922 468014 531978
rect 468082 531922 468138 531978
rect 498678 532294 498734 532350
rect 498802 532294 498858 532350
rect 498678 532170 498734 532226
rect 498802 532170 498858 532226
rect 498678 532046 498734 532102
rect 498802 532046 498858 532102
rect 498678 531922 498734 531978
rect 498802 531922 498858 531978
rect 529398 532294 529454 532350
rect 529522 532294 529578 532350
rect 529398 532170 529454 532226
rect 529522 532170 529578 532226
rect 529398 532046 529454 532102
rect 529522 532046 529578 532102
rect 529398 531922 529454 531978
rect 529522 531922 529578 531978
rect 53238 526294 53294 526350
rect 53362 526294 53418 526350
rect 53238 526170 53294 526226
rect 53362 526170 53418 526226
rect 53238 526046 53294 526102
rect 53362 526046 53418 526102
rect 53238 525922 53294 525978
rect 53362 525922 53418 525978
rect 83958 526294 84014 526350
rect 84082 526294 84138 526350
rect 83958 526170 84014 526226
rect 84082 526170 84138 526226
rect 83958 526046 84014 526102
rect 84082 526046 84138 526102
rect 83958 525922 84014 525978
rect 84082 525922 84138 525978
rect 114678 526294 114734 526350
rect 114802 526294 114858 526350
rect 114678 526170 114734 526226
rect 114802 526170 114858 526226
rect 114678 526046 114734 526102
rect 114802 526046 114858 526102
rect 114678 525922 114734 525978
rect 114802 525922 114858 525978
rect 145398 526294 145454 526350
rect 145522 526294 145578 526350
rect 145398 526170 145454 526226
rect 145522 526170 145578 526226
rect 145398 526046 145454 526102
rect 145522 526046 145578 526102
rect 145398 525922 145454 525978
rect 145522 525922 145578 525978
rect 176118 526294 176174 526350
rect 176242 526294 176298 526350
rect 176118 526170 176174 526226
rect 176242 526170 176298 526226
rect 176118 526046 176174 526102
rect 176242 526046 176298 526102
rect 176118 525922 176174 525978
rect 176242 525922 176298 525978
rect 206838 526294 206894 526350
rect 206962 526294 207018 526350
rect 206838 526170 206894 526226
rect 206962 526170 207018 526226
rect 206838 526046 206894 526102
rect 206962 526046 207018 526102
rect 206838 525922 206894 525978
rect 206962 525922 207018 525978
rect 237558 526294 237614 526350
rect 237682 526294 237738 526350
rect 237558 526170 237614 526226
rect 237682 526170 237738 526226
rect 237558 526046 237614 526102
rect 237682 526046 237738 526102
rect 237558 525922 237614 525978
rect 237682 525922 237738 525978
rect 268278 526294 268334 526350
rect 268402 526294 268458 526350
rect 268278 526170 268334 526226
rect 268402 526170 268458 526226
rect 268278 526046 268334 526102
rect 268402 526046 268458 526102
rect 268278 525922 268334 525978
rect 268402 525922 268458 525978
rect 298998 526294 299054 526350
rect 299122 526294 299178 526350
rect 298998 526170 299054 526226
rect 299122 526170 299178 526226
rect 298998 526046 299054 526102
rect 299122 526046 299178 526102
rect 298998 525922 299054 525978
rect 299122 525922 299178 525978
rect 329718 526294 329774 526350
rect 329842 526294 329898 526350
rect 329718 526170 329774 526226
rect 329842 526170 329898 526226
rect 329718 526046 329774 526102
rect 329842 526046 329898 526102
rect 329718 525922 329774 525978
rect 329842 525922 329898 525978
rect 360438 526294 360494 526350
rect 360562 526294 360618 526350
rect 360438 526170 360494 526226
rect 360562 526170 360618 526226
rect 360438 526046 360494 526102
rect 360562 526046 360618 526102
rect 360438 525922 360494 525978
rect 360562 525922 360618 525978
rect 391158 526294 391214 526350
rect 391282 526294 391338 526350
rect 391158 526170 391214 526226
rect 391282 526170 391338 526226
rect 391158 526046 391214 526102
rect 391282 526046 391338 526102
rect 391158 525922 391214 525978
rect 391282 525922 391338 525978
rect 421878 526294 421934 526350
rect 422002 526294 422058 526350
rect 421878 526170 421934 526226
rect 422002 526170 422058 526226
rect 421878 526046 421934 526102
rect 422002 526046 422058 526102
rect 421878 525922 421934 525978
rect 422002 525922 422058 525978
rect 452598 526294 452654 526350
rect 452722 526294 452778 526350
rect 452598 526170 452654 526226
rect 452722 526170 452778 526226
rect 452598 526046 452654 526102
rect 452722 526046 452778 526102
rect 452598 525922 452654 525978
rect 452722 525922 452778 525978
rect 483318 526294 483374 526350
rect 483442 526294 483498 526350
rect 483318 526170 483374 526226
rect 483442 526170 483498 526226
rect 483318 526046 483374 526102
rect 483442 526046 483498 526102
rect 483318 525922 483374 525978
rect 483442 525922 483498 525978
rect 514038 526294 514094 526350
rect 514162 526294 514218 526350
rect 514038 526170 514094 526226
rect 514162 526170 514218 526226
rect 514038 526046 514094 526102
rect 514162 526046 514218 526102
rect 514038 525922 514094 525978
rect 514162 525922 514218 525978
rect 544758 526294 544814 526350
rect 544882 526294 544938 526350
rect 544758 526170 544814 526226
rect 544882 526170 544938 526226
rect 544758 526046 544814 526102
rect 544882 526046 544938 526102
rect 544758 525922 544814 525978
rect 544882 525922 544938 525978
rect 37878 514294 37934 514350
rect 38002 514294 38058 514350
rect 37878 514170 37934 514226
rect 38002 514170 38058 514226
rect 37878 514046 37934 514102
rect 38002 514046 38058 514102
rect 37878 513922 37934 513978
rect 38002 513922 38058 513978
rect 68598 514294 68654 514350
rect 68722 514294 68778 514350
rect 68598 514170 68654 514226
rect 68722 514170 68778 514226
rect 68598 514046 68654 514102
rect 68722 514046 68778 514102
rect 68598 513922 68654 513978
rect 68722 513922 68778 513978
rect 99318 514294 99374 514350
rect 99442 514294 99498 514350
rect 99318 514170 99374 514226
rect 99442 514170 99498 514226
rect 99318 514046 99374 514102
rect 99442 514046 99498 514102
rect 99318 513922 99374 513978
rect 99442 513922 99498 513978
rect 130038 514294 130094 514350
rect 130162 514294 130218 514350
rect 130038 514170 130094 514226
rect 130162 514170 130218 514226
rect 130038 514046 130094 514102
rect 130162 514046 130218 514102
rect 130038 513922 130094 513978
rect 130162 513922 130218 513978
rect 160758 514294 160814 514350
rect 160882 514294 160938 514350
rect 160758 514170 160814 514226
rect 160882 514170 160938 514226
rect 160758 514046 160814 514102
rect 160882 514046 160938 514102
rect 160758 513922 160814 513978
rect 160882 513922 160938 513978
rect 191478 514294 191534 514350
rect 191602 514294 191658 514350
rect 191478 514170 191534 514226
rect 191602 514170 191658 514226
rect 191478 514046 191534 514102
rect 191602 514046 191658 514102
rect 191478 513922 191534 513978
rect 191602 513922 191658 513978
rect 222198 514294 222254 514350
rect 222322 514294 222378 514350
rect 222198 514170 222254 514226
rect 222322 514170 222378 514226
rect 222198 514046 222254 514102
rect 222322 514046 222378 514102
rect 222198 513922 222254 513978
rect 222322 513922 222378 513978
rect 252918 514294 252974 514350
rect 253042 514294 253098 514350
rect 252918 514170 252974 514226
rect 253042 514170 253098 514226
rect 252918 514046 252974 514102
rect 253042 514046 253098 514102
rect 252918 513922 252974 513978
rect 253042 513922 253098 513978
rect 283638 514294 283694 514350
rect 283762 514294 283818 514350
rect 283638 514170 283694 514226
rect 283762 514170 283818 514226
rect 283638 514046 283694 514102
rect 283762 514046 283818 514102
rect 283638 513922 283694 513978
rect 283762 513922 283818 513978
rect 314358 514294 314414 514350
rect 314482 514294 314538 514350
rect 314358 514170 314414 514226
rect 314482 514170 314538 514226
rect 314358 514046 314414 514102
rect 314482 514046 314538 514102
rect 314358 513922 314414 513978
rect 314482 513922 314538 513978
rect 345078 514294 345134 514350
rect 345202 514294 345258 514350
rect 345078 514170 345134 514226
rect 345202 514170 345258 514226
rect 345078 514046 345134 514102
rect 345202 514046 345258 514102
rect 345078 513922 345134 513978
rect 345202 513922 345258 513978
rect 375798 514294 375854 514350
rect 375922 514294 375978 514350
rect 375798 514170 375854 514226
rect 375922 514170 375978 514226
rect 375798 514046 375854 514102
rect 375922 514046 375978 514102
rect 375798 513922 375854 513978
rect 375922 513922 375978 513978
rect 406518 514294 406574 514350
rect 406642 514294 406698 514350
rect 406518 514170 406574 514226
rect 406642 514170 406698 514226
rect 406518 514046 406574 514102
rect 406642 514046 406698 514102
rect 406518 513922 406574 513978
rect 406642 513922 406698 513978
rect 437238 514294 437294 514350
rect 437362 514294 437418 514350
rect 437238 514170 437294 514226
rect 437362 514170 437418 514226
rect 437238 514046 437294 514102
rect 437362 514046 437418 514102
rect 437238 513922 437294 513978
rect 437362 513922 437418 513978
rect 467958 514294 468014 514350
rect 468082 514294 468138 514350
rect 467958 514170 468014 514226
rect 468082 514170 468138 514226
rect 467958 514046 468014 514102
rect 468082 514046 468138 514102
rect 467958 513922 468014 513978
rect 468082 513922 468138 513978
rect 498678 514294 498734 514350
rect 498802 514294 498858 514350
rect 498678 514170 498734 514226
rect 498802 514170 498858 514226
rect 498678 514046 498734 514102
rect 498802 514046 498858 514102
rect 498678 513922 498734 513978
rect 498802 513922 498858 513978
rect 529398 514294 529454 514350
rect 529522 514294 529578 514350
rect 529398 514170 529454 514226
rect 529522 514170 529578 514226
rect 529398 514046 529454 514102
rect 529522 514046 529578 514102
rect 529398 513922 529454 513978
rect 529522 513922 529578 513978
rect 53238 508294 53294 508350
rect 53362 508294 53418 508350
rect 53238 508170 53294 508226
rect 53362 508170 53418 508226
rect 53238 508046 53294 508102
rect 53362 508046 53418 508102
rect 53238 507922 53294 507978
rect 53362 507922 53418 507978
rect 83958 508294 84014 508350
rect 84082 508294 84138 508350
rect 83958 508170 84014 508226
rect 84082 508170 84138 508226
rect 83958 508046 84014 508102
rect 84082 508046 84138 508102
rect 83958 507922 84014 507978
rect 84082 507922 84138 507978
rect 114678 508294 114734 508350
rect 114802 508294 114858 508350
rect 114678 508170 114734 508226
rect 114802 508170 114858 508226
rect 114678 508046 114734 508102
rect 114802 508046 114858 508102
rect 114678 507922 114734 507978
rect 114802 507922 114858 507978
rect 145398 508294 145454 508350
rect 145522 508294 145578 508350
rect 145398 508170 145454 508226
rect 145522 508170 145578 508226
rect 145398 508046 145454 508102
rect 145522 508046 145578 508102
rect 145398 507922 145454 507978
rect 145522 507922 145578 507978
rect 176118 508294 176174 508350
rect 176242 508294 176298 508350
rect 176118 508170 176174 508226
rect 176242 508170 176298 508226
rect 176118 508046 176174 508102
rect 176242 508046 176298 508102
rect 176118 507922 176174 507978
rect 176242 507922 176298 507978
rect 206838 508294 206894 508350
rect 206962 508294 207018 508350
rect 206838 508170 206894 508226
rect 206962 508170 207018 508226
rect 206838 508046 206894 508102
rect 206962 508046 207018 508102
rect 206838 507922 206894 507978
rect 206962 507922 207018 507978
rect 237558 508294 237614 508350
rect 237682 508294 237738 508350
rect 237558 508170 237614 508226
rect 237682 508170 237738 508226
rect 237558 508046 237614 508102
rect 237682 508046 237738 508102
rect 237558 507922 237614 507978
rect 237682 507922 237738 507978
rect 268278 508294 268334 508350
rect 268402 508294 268458 508350
rect 268278 508170 268334 508226
rect 268402 508170 268458 508226
rect 268278 508046 268334 508102
rect 268402 508046 268458 508102
rect 268278 507922 268334 507978
rect 268402 507922 268458 507978
rect 298998 508294 299054 508350
rect 299122 508294 299178 508350
rect 298998 508170 299054 508226
rect 299122 508170 299178 508226
rect 298998 508046 299054 508102
rect 299122 508046 299178 508102
rect 298998 507922 299054 507978
rect 299122 507922 299178 507978
rect 329718 508294 329774 508350
rect 329842 508294 329898 508350
rect 329718 508170 329774 508226
rect 329842 508170 329898 508226
rect 329718 508046 329774 508102
rect 329842 508046 329898 508102
rect 329718 507922 329774 507978
rect 329842 507922 329898 507978
rect 360438 508294 360494 508350
rect 360562 508294 360618 508350
rect 360438 508170 360494 508226
rect 360562 508170 360618 508226
rect 360438 508046 360494 508102
rect 360562 508046 360618 508102
rect 360438 507922 360494 507978
rect 360562 507922 360618 507978
rect 391158 508294 391214 508350
rect 391282 508294 391338 508350
rect 391158 508170 391214 508226
rect 391282 508170 391338 508226
rect 391158 508046 391214 508102
rect 391282 508046 391338 508102
rect 391158 507922 391214 507978
rect 391282 507922 391338 507978
rect 421878 508294 421934 508350
rect 422002 508294 422058 508350
rect 421878 508170 421934 508226
rect 422002 508170 422058 508226
rect 421878 508046 421934 508102
rect 422002 508046 422058 508102
rect 421878 507922 421934 507978
rect 422002 507922 422058 507978
rect 452598 508294 452654 508350
rect 452722 508294 452778 508350
rect 452598 508170 452654 508226
rect 452722 508170 452778 508226
rect 452598 508046 452654 508102
rect 452722 508046 452778 508102
rect 452598 507922 452654 507978
rect 452722 507922 452778 507978
rect 483318 508294 483374 508350
rect 483442 508294 483498 508350
rect 483318 508170 483374 508226
rect 483442 508170 483498 508226
rect 483318 508046 483374 508102
rect 483442 508046 483498 508102
rect 483318 507922 483374 507978
rect 483442 507922 483498 507978
rect 514038 508294 514094 508350
rect 514162 508294 514218 508350
rect 514038 508170 514094 508226
rect 514162 508170 514218 508226
rect 514038 508046 514094 508102
rect 514162 508046 514218 508102
rect 514038 507922 514094 507978
rect 514162 507922 514218 507978
rect 544758 508294 544814 508350
rect 544882 508294 544938 508350
rect 544758 508170 544814 508226
rect 544882 508170 544938 508226
rect 544758 508046 544814 508102
rect 544882 508046 544938 508102
rect 544758 507922 544814 507978
rect 544882 507922 544938 507978
rect 37878 496294 37934 496350
rect 38002 496294 38058 496350
rect 37878 496170 37934 496226
rect 38002 496170 38058 496226
rect 37878 496046 37934 496102
rect 38002 496046 38058 496102
rect 37878 495922 37934 495978
rect 38002 495922 38058 495978
rect 68598 496294 68654 496350
rect 68722 496294 68778 496350
rect 68598 496170 68654 496226
rect 68722 496170 68778 496226
rect 68598 496046 68654 496102
rect 68722 496046 68778 496102
rect 68598 495922 68654 495978
rect 68722 495922 68778 495978
rect 99318 496294 99374 496350
rect 99442 496294 99498 496350
rect 99318 496170 99374 496226
rect 99442 496170 99498 496226
rect 99318 496046 99374 496102
rect 99442 496046 99498 496102
rect 99318 495922 99374 495978
rect 99442 495922 99498 495978
rect 130038 496294 130094 496350
rect 130162 496294 130218 496350
rect 130038 496170 130094 496226
rect 130162 496170 130218 496226
rect 130038 496046 130094 496102
rect 130162 496046 130218 496102
rect 130038 495922 130094 495978
rect 130162 495922 130218 495978
rect 160758 496294 160814 496350
rect 160882 496294 160938 496350
rect 160758 496170 160814 496226
rect 160882 496170 160938 496226
rect 160758 496046 160814 496102
rect 160882 496046 160938 496102
rect 160758 495922 160814 495978
rect 160882 495922 160938 495978
rect 191478 496294 191534 496350
rect 191602 496294 191658 496350
rect 191478 496170 191534 496226
rect 191602 496170 191658 496226
rect 191478 496046 191534 496102
rect 191602 496046 191658 496102
rect 191478 495922 191534 495978
rect 191602 495922 191658 495978
rect 222198 496294 222254 496350
rect 222322 496294 222378 496350
rect 222198 496170 222254 496226
rect 222322 496170 222378 496226
rect 222198 496046 222254 496102
rect 222322 496046 222378 496102
rect 222198 495922 222254 495978
rect 222322 495922 222378 495978
rect 252918 496294 252974 496350
rect 253042 496294 253098 496350
rect 252918 496170 252974 496226
rect 253042 496170 253098 496226
rect 252918 496046 252974 496102
rect 253042 496046 253098 496102
rect 252918 495922 252974 495978
rect 253042 495922 253098 495978
rect 283638 496294 283694 496350
rect 283762 496294 283818 496350
rect 283638 496170 283694 496226
rect 283762 496170 283818 496226
rect 283638 496046 283694 496102
rect 283762 496046 283818 496102
rect 283638 495922 283694 495978
rect 283762 495922 283818 495978
rect 314358 496294 314414 496350
rect 314482 496294 314538 496350
rect 314358 496170 314414 496226
rect 314482 496170 314538 496226
rect 314358 496046 314414 496102
rect 314482 496046 314538 496102
rect 314358 495922 314414 495978
rect 314482 495922 314538 495978
rect 345078 496294 345134 496350
rect 345202 496294 345258 496350
rect 345078 496170 345134 496226
rect 345202 496170 345258 496226
rect 345078 496046 345134 496102
rect 345202 496046 345258 496102
rect 345078 495922 345134 495978
rect 345202 495922 345258 495978
rect 375798 496294 375854 496350
rect 375922 496294 375978 496350
rect 375798 496170 375854 496226
rect 375922 496170 375978 496226
rect 375798 496046 375854 496102
rect 375922 496046 375978 496102
rect 375798 495922 375854 495978
rect 375922 495922 375978 495978
rect 406518 496294 406574 496350
rect 406642 496294 406698 496350
rect 406518 496170 406574 496226
rect 406642 496170 406698 496226
rect 406518 496046 406574 496102
rect 406642 496046 406698 496102
rect 406518 495922 406574 495978
rect 406642 495922 406698 495978
rect 437238 496294 437294 496350
rect 437362 496294 437418 496350
rect 437238 496170 437294 496226
rect 437362 496170 437418 496226
rect 437238 496046 437294 496102
rect 437362 496046 437418 496102
rect 437238 495922 437294 495978
rect 437362 495922 437418 495978
rect 467958 496294 468014 496350
rect 468082 496294 468138 496350
rect 467958 496170 468014 496226
rect 468082 496170 468138 496226
rect 467958 496046 468014 496102
rect 468082 496046 468138 496102
rect 467958 495922 468014 495978
rect 468082 495922 468138 495978
rect 498678 496294 498734 496350
rect 498802 496294 498858 496350
rect 498678 496170 498734 496226
rect 498802 496170 498858 496226
rect 498678 496046 498734 496102
rect 498802 496046 498858 496102
rect 498678 495922 498734 495978
rect 498802 495922 498858 495978
rect 529398 496294 529454 496350
rect 529522 496294 529578 496350
rect 529398 496170 529454 496226
rect 529522 496170 529578 496226
rect 529398 496046 529454 496102
rect 529522 496046 529578 496102
rect 529398 495922 529454 495978
rect 529522 495922 529578 495978
rect 53238 490294 53294 490350
rect 53362 490294 53418 490350
rect 53238 490170 53294 490226
rect 53362 490170 53418 490226
rect 53238 490046 53294 490102
rect 53362 490046 53418 490102
rect 53238 489922 53294 489978
rect 53362 489922 53418 489978
rect 83958 490294 84014 490350
rect 84082 490294 84138 490350
rect 83958 490170 84014 490226
rect 84082 490170 84138 490226
rect 83958 490046 84014 490102
rect 84082 490046 84138 490102
rect 83958 489922 84014 489978
rect 84082 489922 84138 489978
rect 114678 490294 114734 490350
rect 114802 490294 114858 490350
rect 114678 490170 114734 490226
rect 114802 490170 114858 490226
rect 114678 490046 114734 490102
rect 114802 490046 114858 490102
rect 114678 489922 114734 489978
rect 114802 489922 114858 489978
rect 145398 490294 145454 490350
rect 145522 490294 145578 490350
rect 145398 490170 145454 490226
rect 145522 490170 145578 490226
rect 145398 490046 145454 490102
rect 145522 490046 145578 490102
rect 145398 489922 145454 489978
rect 145522 489922 145578 489978
rect 176118 490294 176174 490350
rect 176242 490294 176298 490350
rect 176118 490170 176174 490226
rect 176242 490170 176298 490226
rect 176118 490046 176174 490102
rect 176242 490046 176298 490102
rect 176118 489922 176174 489978
rect 176242 489922 176298 489978
rect 206838 490294 206894 490350
rect 206962 490294 207018 490350
rect 206838 490170 206894 490226
rect 206962 490170 207018 490226
rect 206838 490046 206894 490102
rect 206962 490046 207018 490102
rect 206838 489922 206894 489978
rect 206962 489922 207018 489978
rect 237558 490294 237614 490350
rect 237682 490294 237738 490350
rect 237558 490170 237614 490226
rect 237682 490170 237738 490226
rect 237558 490046 237614 490102
rect 237682 490046 237738 490102
rect 237558 489922 237614 489978
rect 237682 489922 237738 489978
rect 268278 490294 268334 490350
rect 268402 490294 268458 490350
rect 268278 490170 268334 490226
rect 268402 490170 268458 490226
rect 268278 490046 268334 490102
rect 268402 490046 268458 490102
rect 268278 489922 268334 489978
rect 268402 489922 268458 489978
rect 298998 490294 299054 490350
rect 299122 490294 299178 490350
rect 298998 490170 299054 490226
rect 299122 490170 299178 490226
rect 298998 490046 299054 490102
rect 299122 490046 299178 490102
rect 298998 489922 299054 489978
rect 299122 489922 299178 489978
rect 329718 490294 329774 490350
rect 329842 490294 329898 490350
rect 329718 490170 329774 490226
rect 329842 490170 329898 490226
rect 329718 490046 329774 490102
rect 329842 490046 329898 490102
rect 329718 489922 329774 489978
rect 329842 489922 329898 489978
rect 360438 490294 360494 490350
rect 360562 490294 360618 490350
rect 360438 490170 360494 490226
rect 360562 490170 360618 490226
rect 360438 490046 360494 490102
rect 360562 490046 360618 490102
rect 360438 489922 360494 489978
rect 360562 489922 360618 489978
rect 391158 490294 391214 490350
rect 391282 490294 391338 490350
rect 391158 490170 391214 490226
rect 391282 490170 391338 490226
rect 391158 490046 391214 490102
rect 391282 490046 391338 490102
rect 391158 489922 391214 489978
rect 391282 489922 391338 489978
rect 421878 490294 421934 490350
rect 422002 490294 422058 490350
rect 421878 490170 421934 490226
rect 422002 490170 422058 490226
rect 421878 490046 421934 490102
rect 422002 490046 422058 490102
rect 421878 489922 421934 489978
rect 422002 489922 422058 489978
rect 452598 490294 452654 490350
rect 452722 490294 452778 490350
rect 452598 490170 452654 490226
rect 452722 490170 452778 490226
rect 452598 490046 452654 490102
rect 452722 490046 452778 490102
rect 452598 489922 452654 489978
rect 452722 489922 452778 489978
rect 483318 490294 483374 490350
rect 483442 490294 483498 490350
rect 483318 490170 483374 490226
rect 483442 490170 483498 490226
rect 483318 490046 483374 490102
rect 483442 490046 483498 490102
rect 483318 489922 483374 489978
rect 483442 489922 483498 489978
rect 514038 490294 514094 490350
rect 514162 490294 514218 490350
rect 514038 490170 514094 490226
rect 514162 490170 514218 490226
rect 514038 490046 514094 490102
rect 514162 490046 514218 490102
rect 514038 489922 514094 489978
rect 514162 489922 514218 489978
rect 544758 490294 544814 490350
rect 544882 490294 544938 490350
rect 544758 490170 544814 490226
rect 544882 490170 544938 490226
rect 544758 490046 544814 490102
rect 544882 490046 544938 490102
rect 544758 489922 544814 489978
rect 544882 489922 544938 489978
rect 37878 478294 37934 478350
rect 38002 478294 38058 478350
rect 37878 478170 37934 478226
rect 38002 478170 38058 478226
rect 37878 478046 37934 478102
rect 38002 478046 38058 478102
rect 37878 477922 37934 477978
rect 38002 477922 38058 477978
rect 68598 478294 68654 478350
rect 68722 478294 68778 478350
rect 68598 478170 68654 478226
rect 68722 478170 68778 478226
rect 68598 478046 68654 478102
rect 68722 478046 68778 478102
rect 68598 477922 68654 477978
rect 68722 477922 68778 477978
rect 99318 478294 99374 478350
rect 99442 478294 99498 478350
rect 99318 478170 99374 478226
rect 99442 478170 99498 478226
rect 99318 478046 99374 478102
rect 99442 478046 99498 478102
rect 99318 477922 99374 477978
rect 99442 477922 99498 477978
rect 130038 478294 130094 478350
rect 130162 478294 130218 478350
rect 130038 478170 130094 478226
rect 130162 478170 130218 478226
rect 130038 478046 130094 478102
rect 130162 478046 130218 478102
rect 130038 477922 130094 477978
rect 130162 477922 130218 477978
rect 160758 478294 160814 478350
rect 160882 478294 160938 478350
rect 160758 478170 160814 478226
rect 160882 478170 160938 478226
rect 160758 478046 160814 478102
rect 160882 478046 160938 478102
rect 160758 477922 160814 477978
rect 160882 477922 160938 477978
rect 191478 478294 191534 478350
rect 191602 478294 191658 478350
rect 191478 478170 191534 478226
rect 191602 478170 191658 478226
rect 191478 478046 191534 478102
rect 191602 478046 191658 478102
rect 191478 477922 191534 477978
rect 191602 477922 191658 477978
rect 222198 478294 222254 478350
rect 222322 478294 222378 478350
rect 222198 478170 222254 478226
rect 222322 478170 222378 478226
rect 222198 478046 222254 478102
rect 222322 478046 222378 478102
rect 222198 477922 222254 477978
rect 222322 477922 222378 477978
rect 252918 478294 252974 478350
rect 253042 478294 253098 478350
rect 252918 478170 252974 478226
rect 253042 478170 253098 478226
rect 252918 478046 252974 478102
rect 253042 478046 253098 478102
rect 252918 477922 252974 477978
rect 253042 477922 253098 477978
rect 283638 478294 283694 478350
rect 283762 478294 283818 478350
rect 283638 478170 283694 478226
rect 283762 478170 283818 478226
rect 283638 478046 283694 478102
rect 283762 478046 283818 478102
rect 283638 477922 283694 477978
rect 283762 477922 283818 477978
rect 314358 478294 314414 478350
rect 314482 478294 314538 478350
rect 314358 478170 314414 478226
rect 314482 478170 314538 478226
rect 314358 478046 314414 478102
rect 314482 478046 314538 478102
rect 314358 477922 314414 477978
rect 314482 477922 314538 477978
rect 345078 478294 345134 478350
rect 345202 478294 345258 478350
rect 345078 478170 345134 478226
rect 345202 478170 345258 478226
rect 345078 478046 345134 478102
rect 345202 478046 345258 478102
rect 345078 477922 345134 477978
rect 345202 477922 345258 477978
rect 375798 478294 375854 478350
rect 375922 478294 375978 478350
rect 375798 478170 375854 478226
rect 375922 478170 375978 478226
rect 375798 478046 375854 478102
rect 375922 478046 375978 478102
rect 375798 477922 375854 477978
rect 375922 477922 375978 477978
rect 406518 478294 406574 478350
rect 406642 478294 406698 478350
rect 406518 478170 406574 478226
rect 406642 478170 406698 478226
rect 406518 478046 406574 478102
rect 406642 478046 406698 478102
rect 406518 477922 406574 477978
rect 406642 477922 406698 477978
rect 437238 478294 437294 478350
rect 437362 478294 437418 478350
rect 437238 478170 437294 478226
rect 437362 478170 437418 478226
rect 437238 478046 437294 478102
rect 437362 478046 437418 478102
rect 437238 477922 437294 477978
rect 437362 477922 437418 477978
rect 467958 478294 468014 478350
rect 468082 478294 468138 478350
rect 467958 478170 468014 478226
rect 468082 478170 468138 478226
rect 467958 478046 468014 478102
rect 468082 478046 468138 478102
rect 467958 477922 468014 477978
rect 468082 477922 468138 477978
rect 498678 478294 498734 478350
rect 498802 478294 498858 478350
rect 498678 478170 498734 478226
rect 498802 478170 498858 478226
rect 498678 478046 498734 478102
rect 498802 478046 498858 478102
rect 498678 477922 498734 477978
rect 498802 477922 498858 477978
rect 529398 478294 529454 478350
rect 529522 478294 529578 478350
rect 529398 478170 529454 478226
rect 529522 478170 529578 478226
rect 529398 478046 529454 478102
rect 529522 478046 529578 478102
rect 529398 477922 529454 477978
rect 529522 477922 529578 477978
rect 53238 472294 53294 472350
rect 53362 472294 53418 472350
rect 53238 472170 53294 472226
rect 53362 472170 53418 472226
rect 53238 472046 53294 472102
rect 53362 472046 53418 472102
rect 53238 471922 53294 471978
rect 53362 471922 53418 471978
rect 83958 472294 84014 472350
rect 84082 472294 84138 472350
rect 83958 472170 84014 472226
rect 84082 472170 84138 472226
rect 83958 472046 84014 472102
rect 84082 472046 84138 472102
rect 83958 471922 84014 471978
rect 84082 471922 84138 471978
rect 114678 472294 114734 472350
rect 114802 472294 114858 472350
rect 114678 472170 114734 472226
rect 114802 472170 114858 472226
rect 114678 472046 114734 472102
rect 114802 472046 114858 472102
rect 114678 471922 114734 471978
rect 114802 471922 114858 471978
rect 145398 472294 145454 472350
rect 145522 472294 145578 472350
rect 145398 472170 145454 472226
rect 145522 472170 145578 472226
rect 145398 472046 145454 472102
rect 145522 472046 145578 472102
rect 145398 471922 145454 471978
rect 145522 471922 145578 471978
rect 176118 472294 176174 472350
rect 176242 472294 176298 472350
rect 176118 472170 176174 472226
rect 176242 472170 176298 472226
rect 176118 472046 176174 472102
rect 176242 472046 176298 472102
rect 176118 471922 176174 471978
rect 176242 471922 176298 471978
rect 206838 472294 206894 472350
rect 206962 472294 207018 472350
rect 206838 472170 206894 472226
rect 206962 472170 207018 472226
rect 206838 472046 206894 472102
rect 206962 472046 207018 472102
rect 206838 471922 206894 471978
rect 206962 471922 207018 471978
rect 237558 472294 237614 472350
rect 237682 472294 237738 472350
rect 237558 472170 237614 472226
rect 237682 472170 237738 472226
rect 237558 472046 237614 472102
rect 237682 472046 237738 472102
rect 237558 471922 237614 471978
rect 237682 471922 237738 471978
rect 268278 472294 268334 472350
rect 268402 472294 268458 472350
rect 268278 472170 268334 472226
rect 268402 472170 268458 472226
rect 268278 472046 268334 472102
rect 268402 472046 268458 472102
rect 268278 471922 268334 471978
rect 268402 471922 268458 471978
rect 298998 472294 299054 472350
rect 299122 472294 299178 472350
rect 298998 472170 299054 472226
rect 299122 472170 299178 472226
rect 298998 472046 299054 472102
rect 299122 472046 299178 472102
rect 298998 471922 299054 471978
rect 299122 471922 299178 471978
rect 329718 472294 329774 472350
rect 329842 472294 329898 472350
rect 329718 472170 329774 472226
rect 329842 472170 329898 472226
rect 329718 472046 329774 472102
rect 329842 472046 329898 472102
rect 329718 471922 329774 471978
rect 329842 471922 329898 471978
rect 360438 472294 360494 472350
rect 360562 472294 360618 472350
rect 360438 472170 360494 472226
rect 360562 472170 360618 472226
rect 360438 472046 360494 472102
rect 360562 472046 360618 472102
rect 360438 471922 360494 471978
rect 360562 471922 360618 471978
rect 391158 472294 391214 472350
rect 391282 472294 391338 472350
rect 391158 472170 391214 472226
rect 391282 472170 391338 472226
rect 391158 472046 391214 472102
rect 391282 472046 391338 472102
rect 391158 471922 391214 471978
rect 391282 471922 391338 471978
rect 421878 472294 421934 472350
rect 422002 472294 422058 472350
rect 421878 472170 421934 472226
rect 422002 472170 422058 472226
rect 421878 472046 421934 472102
rect 422002 472046 422058 472102
rect 421878 471922 421934 471978
rect 422002 471922 422058 471978
rect 452598 472294 452654 472350
rect 452722 472294 452778 472350
rect 452598 472170 452654 472226
rect 452722 472170 452778 472226
rect 452598 472046 452654 472102
rect 452722 472046 452778 472102
rect 452598 471922 452654 471978
rect 452722 471922 452778 471978
rect 483318 472294 483374 472350
rect 483442 472294 483498 472350
rect 483318 472170 483374 472226
rect 483442 472170 483498 472226
rect 483318 472046 483374 472102
rect 483442 472046 483498 472102
rect 483318 471922 483374 471978
rect 483442 471922 483498 471978
rect 514038 472294 514094 472350
rect 514162 472294 514218 472350
rect 514038 472170 514094 472226
rect 514162 472170 514218 472226
rect 514038 472046 514094 472102
rect 514162 472046 514218 472102
rect 514038 471922 514094 471978
rect 514162 471922 514218 471978
rect 544758 472294 544814 472350
rect 544882 472294 544938 472350
rect 544758 472170 544814 472226
rect 544882 472170 544938 472226
rect 544758 472046 544814 472102
rect 544882 472046 544938 472102
rect 544758 471922 544814 471978
rect 544882 471922 544938 471978
rect 37878 460294 37934 460350
rect 38002 460294 38058 460350
rect 37878 460170 37934 460226
rect 38002 460170 38058 460226
rect 37878 460046 37934 460102
rect 38002 460046 38058 460102
rect 37878 459922 37934 459978
rect 38002 459922 38058 459978
rect 68598 460294 68654 460350
rect 68722 460294 68778 460350
rect 68598 460170 68654 460226
rect 68722 460170 68778 460226
rect 68598 460046 68654 460102
rect 68722 460046 68778 460102
rect 68598 459922 68654 459978
rect 68722 459922 68778 459978
rect 99318 460294 99374 460350
rect 99442 460294 99498 460350
rect 99318 460170 99374 460226
rect 99442 460170 99498 460226
rect 99318 460046 99374 460102
rect 99442 460046 99498 460102
rect 99318 459922 99374 459978
rect 99442 459922 99498 459978
rect 130038 460294 130094 460350
rect 130162 460294 130218 460350
rect 130038 460170 130094 460226
rect 130162 460170 130218 460226
rect 130038 460046 130094 460102
rect 130162 460046 130218 460102
rect 130038 459922 130094 459978
rect 130162 459922 130218 459978
rect 160758 460294 160814 460350
rect 160882 460294 160938 460350
rect 160758 460170 160814 460226
rect 160882 460170 160938 460226
rect 160758 460046 160814 460102
rect 160882 460046 160938 460102
rect 160758 459922 160814 459978
rect 160882 459922 160938 459978
rect 191478 460294 191534 460350
rect 191602 460294 191658 460350
rect 191478 460170 191534 460226
rect 191602 460170 191658 460226
rect 191478 460046 191534 460102
rect 191602 460046 191658 460102
rect 191478 459922 191534 459978
rect 191602 459922 191658 459978
rect 222198 460294 222254 460350
rect 222322 460294 222378 460350
rect 222198 460170 222254 460226
rect 222322 460170 222378 460226
rect 222198 460046 222254 460102
rect 222322 460046 222378 460102
rect 222198 459922 222254 459978
rect 222322 459922 222378 459978
rect 252918 460294 252974 460350
rect 253042 460294 253098 460350
rect 252918 460170 252974 460226
rect 253042 460170 253098 460226
rect 252918 460046 252974 460102
rect 253042 460046 253098 460102
rect 252918 459922 252974 459978
rect 253042 459922 253098 459978
rect 283638 460294 283694 460350
rect 283762 460294 283818 460350
rect 283638 460170 283694 460226
rect 283762 460170 283818 460226
rect 283638 460046 283694 460102
rect 283762 460046 283818 460102
rect 283638 459922 283694 459978
rect 283762 459922 283818 459978
rect 314358 460294 314414 460350
rect 314482 460294 314538 460350
rect 314358 460170 314414 460226
rect 314482 460170 314538 460226
rect 314358 460046 314414 460102
rect 314482 460046 314538 460102
rect 314358 459922 314414 459978
rect 314482 459922 314538 459978
rect 345078 460294 345134 460350
rect 345202 460294 345258 460350
rect 345078 460170 345134 460226
rect 345202 460170 345258 460226
rect 345078 460046 345134 460102
rect 345202 460046 345258 460102
rect 345078 459922 345134 459978
rect 345202 459922 345258 459978
rect 375798 460294 375854 460350
rect 375922 460294 375978 460350
rect 375798 460170 375854 460226
rect 375922 460170 375978 460226
rect 375798 460046 375854 460102
rect 375922 460046 375978 460102
rect 375798 459922 375854 459978
rect 375922 459922 375978 459978
rect 406518 460294 406574 460350
rect 406642 460294 406698 460350
rect 406518 460170 406574 460226
rect 406642 460170 406698 460226
rect 406518 460046 406574 460102
rect 406642 460046 406698 460102
rect 406518 459922 406574 459978
rect 406642 459922 406698 459978
rect 437238 460294 437294 460350
rect 437362 460294 437418 460350
rect 437238 460170 437294 460226
rect 437362 460170 437418 460226
rect 437238 460046 437294 460102
rect 437362 460046 437418 460102
rect 437238 459922 437294 459978
rect 437362 459922 437418 459978
rect 467958 460294 468014 460350
rect 468082 460294 468138 460350
rect 467958 460170 468014 460226
rect 468082 460170 468138 460226
rect 467958 460046 468014 460102
rect 468082 460046 468138 460102
rect 467958 459922 468014 459978
rect 468082 459922 468138 459978
rect 498678 460294 498734 460350
rect 498802 460294 498858 460350
rect 498678 460170 498734 460226
rect 498802 460170 498858 460226
rect 498678 460046 498734 460102
rect 498802 460046 498858 460102
rect 498678 459922 498734 459978
rect 498802 459922 498858 459978
rect 529398 460294 529454 460350
rect 529522 460294 529578 460350
rect 529398 460170 529454 460226
rect 529522 460170 529578 460226
rect 529398 460046 529454 460102
rect 529522 460046 529578 460102
rect 529398 459922 529454 459978
rect 529522 459922 529578 459978
rect 53238 454294 53294 454350
rect 53362 454294 53418 454350
rect 53238 454170 53294 454226
rect 53362 454170 53418 454226
rect 53238 454046 53294 454102
rect 53362 454046 53418 454102
rect 53238 453922 53294 453978
rect 53362 453922 53418 453978
rect 83958 454294 84014 454350
rect 84082 454294 84138 454350
rect 83958 454170 84014 454226
rect 84082 454170 84138 454226
rect 83958 454046 84014 454102
rect 84082 454046 84138 454102
rect 83958 453922 84014 453978
rect 84082 453922 84138 453978
rect 114678 454294 114734 454350
rect 114802 454294 114858 454350
rect 114678 454170 114734 454226
rect 114802 454170 114858 454226
rect 114678 454046 114734 454102
rect 114802 454046 114858 454102
rect 114678 453922 114734 453978
rect 114802 453922 114858 453978
rect 145398 454294 145454 454350
rect 145522 454294 145578 454350
rect 145398 454170 145454 454226
rect 145522 454170 145578 454226
rect 145398 454046 145454 454102
rect 145522 454046 145578 454102
rect 145398 453922 145454 453978
rect 145522 453922 145578 453978
rect 176118 454294 176174 454350
rect 176242 454294 176298 454350
rect 176118 454170 176174 454226
rect 176242 454170 176298 454226
rect 176118 454046 176174 454102
rect 176242 454046 176298 454102
rect 176118 453922 176174 453978
rect 176242 453922 176298 453978
rect 206838 454294 206894 454350
rect 206962 454294 207018 454350
rect 206838 454170 206894 454226
rect 206962 454170 207018 454226
rect 206838 454046 206894 454102
rect 206962 454046 207018 454102
rect 206838 453922 206894 453978
rect 206962 453922 207018 453978
rect 237558 454294 237614 454350
rect 237682 454294 237738 454350
rect 237558 454170 237614 454226
rect 237682 454170 237738 454226
rect 237558 454046 237614 454102
rect 237682 454046 237738 454102
rect 237558 453922 237614 453978
rect 237682 453922 237738 453978
rect 268278 454294 268334 454350
rect 268402 454294 268458 454350
rect 268278 454170 268334 454226
rect 268402 454170 268458 454226
rect 268278 454046 268334 454102
rect 268402 454046 268458 454102
rect 268278 453922 268334 453978
rect 268402 453922 268458 453978
rect 298998 454294 299054 454350
rect 299122 454294 299178 454350
rect 298998 454170 299054 454226
rect 299122 454170 299178 454226
rect 298998 454046 299054 454102
rect 299122 454046 299178 454102
rect 298998 453922 299054 453978
rect 299122 453922 299178 453978
rect 329718 454294 329774 454350
rect 329842 454294 329898 454350
rect 329718 454170 329774 454226
rect 329842 454170 329898 454226
rect 329718 454046 329774 454102
rect 329842 454046 329898 454102
rect 329718 453922 329774 453978
rect 329842 453922 329898 453978
rect 360438 454294 360494 454350
rect 360562 454294 360618 454350
rect 360438 454170 360494 454226
rect 360562 454170 360618 454226
rect 360438 454046 360494 454102
rect 360562 454046 360618 454102
rect 360438 453922 360494 453978
rect 360562 453922 360618 453978
rect 391158 454294 391214 454350
rect 391282 454294 391338 454350
rect 391158 454170 391214 454226
rect 391282 454170 391338 454226
rect 391158 454046 391214 454102
rect 391282 454046 391338 454102
rect 391158 453922 391214 453978
rect 391282 453922 391338 453978
rect 421878 454294 421934 454350
rect 422002 454294 422058 454350
rect 421878 454170 421934 454226
rect 422002 454170 422058 454226
rect 421878 454046 421934 454102
rect 422002 454046 422058 454102
rect 421878 453922 421934 453978
rect 422002 453922 422058 453978
rect 452598 454294 452654 454350
rect 452722 454294 452778 454350
rect 452598 454170 452654 454226
rect 452722 454170 452778 454226
rect 452598 454046 452654 454102
rect 452722 454046 452778 454102
rect 452598 453922 452654 453978
rect 452722 453922 452778 453978
rect 483318 454294 483374 454350
rect 483442 454294 483498 454350
rect 483318 454170 483374 454226
rect 483442 454170 483498 454226
rect 483318 454046 483374 454102
rect 483442 454046 483498 454102
rect 483318 453922 483374 453978
rect 483442 453922 483498 453978
rect 514038 454294 514094 454350
rect 514162 454294 514218 454350
rect 514038 454170 514094 454226
rect 514162 454170 514218 454226
rect 514038 454046 514094 454102
rect 514162 454046 514218 454102
rect 514038 453922 514094 453978
rect 514162 453922 514218 453978
rect 544758 454294 544814 454350
rect 544882 454294 544938 454350
rect 544758 454170 544814 454226
rect 544882 454170 544938 454226
rect 544758 454046 544814 454102
rect 544882 454046 544938 454102
rect 544758 453922 544814 453978
rect 544882 453922 544938 453978
rect 37878 442294 37934 442350
rect 38002 442294 38058 442350
rect 37878 442170 37934 442226
rect 38002 442170 38058 442226
rect 37878 442046 37934 442102
rect 38002 442046 38058 442102
rect 37878 441922 37934 441978
rect 38002 441922 38058 441978
rect 68598 442294 68654 442350
rect 68722 442294 68778 442350
rect 68598 442170 68654 442226
rect 68722 442170 68778 442226
rect 68598 442046 68654 442102
rect 68722 442046 68778 442102
rect 68598 441922 68654 441978
rect 68722 441922 68778 441978
rect 99318 442294 99374 442350
rect 99442 442294 99498 442350
rect 99318 442170 99374 442226
rect 99442 442170 99498 442226
rect 99318 442046 99374 442102
rect 99442 442046 99498 442102
rect 99318 441922 99374 441978
rect 99442 441922 99498 441978
rect 130038 442294 130094 442350
rect 130162 442294 130218 442350
rect 130038 442170 130094 442226
rect 130162 442170 130218 442226
rect 130038 442046 130094 442102
rect 130162 442046 130218 442102
rect 130038 441922 130094 441978
rect 130162 441922 130218 441978
rect 160758 442294 160814 442350
rect 160882 442294 160938 442350
rect 160758 442170 160814 442226
rect 160882 442170 160938 442226
rect 160758 442046 160814 442102
rect 160882 442046 160938 442102
rect 160758 441922 160814 441978
rect 160882 441922 160938 441978
rect 191478 442294 191534 442350
rect 191602 442294 191658 442350
rect 191478 442170 191534 442226
rect 191602 442170 191658 442226
rect 191478 442046 191534 442102
rect 191602 442046 191658 442102
rect 191478 441922 191534 441978
rect 191602 441922 191658 441978
rect 222198 442294 222254 442350
rect 222322 442294 222378 442350
rect 222198 442170 222254 442226
rect 222322 442170 222378 442226
rect 222198 442046 222254 442102
rect 222322 442046 222378 442102
rect 222198 441922 222254 441978
rect 222322 441922 222378 441978
rect 252918 442294 252974 442350
rect 253042 442294 253098 442350
rect 252918 442170 252974 442226
rect 253042 442170 253098 442226
rect 252918 442046 252974 442102
rect 253042 442046 253098 442102
rect 252918 441922 252974 441978
rect 253042 441922 253098 441978
rect 283638 442294 283694 442350
rect 283762 442294 283818 442350
rect 283638 442170 283694 442226
rect 283762 442170 283818 442226
rect 283638 442046 283694 442102
rect 283762 442046 283818 442102
rect 283638 441922 283694 441978
rect 283762 441922 283818 441978
rect 314358 442294 314414 442350
rect 314482 442294 314538 442350
rect 314358 442170 314414 442226
rect 314482 442170 314538 442226
rect 314358 442046 314414 442102
rect 314482 442046 314538 442102
rect 314358 441922 314414 441978
rect 314482 441922 314538 441978
rect 345078 442294 345134 442350
rect 345202 442294 345258 442350
rect 345078 442170 345134 442226
rect 345202 442170 345258 442226
rect 345078 442046 345134 442102
rect 345202 442046 345258 442102
rect 345078 441922 345134 441978
rect 345202 441922 345258 441978
rect 375798 442294 375854 442350
rect 375922 442294 375978 442350
rect 375798 442170 375854 442226
rect 375922 442170 375978 442226
rect 375798 442046 375854 442102
rect 375922 442046 375978 442102
rect 375798 441922 375854 441978
rect 375922 441922 375978 441978
rect 406518 442294 406574 442350
rect 406642 442294 406698 442350
rect 406518 442170 406574 442226
rect 406642 442170 406698 442226
rect 406518 442046 406574 442102
rect 406642 442046 406698 442102
rect 406518 441922 406574 441978
rect 406642 441922 406698 441978
rect 437238 442294 437294 442350
rect 437362 442294 437418 442350
rect 437238 442170 437294 442226
rect 437362 442170 437418 442226
rect 437238 442046 437294 442102
rect 437362 442046 437418 442102
rect 437238 441922 437294 441978
rect 437362 441922 437418 441978
rect 467958 442294 468014 442350
rect 468082 442294 468138 442350
rect 467958 442170 468014 442226
rect 468082 442170 468138 442226
rect 467958 442046 468014 442102
rect 468082 442046 468138 442102
rect 467958 441922 468014 441978
rect 468082 441922 468138 441978
rect 498678 442294 498734 442350
rect 498802 442294 498858 442350
rect 498678 442170 498734 442226
rect 498802 442170 498858 442226
rect 498678 442046 498734 442102
rect 498802 442046 498858 442102
rect 498678 441922 498734 441978
rect 498802 441922 498858 441978
rect 529398 442294 529454 442350
rect 529522 442294 529578 442350
rect 529398 442170 529454 442226
rect 529522 442170 529578 442226
rect 529398 442046 529454 442102
rect 529522 442046 529578 442102
rect 529398 441922 529454 441978
rect 529522 441922 529578 441978
rect 53238 436294 53294 436350
rect 53362 436294 53418 436350
rect 53238 436170 53294 436226
rect 53362 436170 53418 436226
rect 53238 436046 53294 436102
rect 53362 436046 53418 436102
rect 53238 435922 53294 435978
rect 53362 435922 53418 435978
rect 83958 436294 84014 436350
rect 84082 436294 84138 436350
rect 83958 436170 84014 436226
rect 84082 436170 84138 436226
rect 83958 436046 84014 436102
rect 84082 436046 84138 436102
rect 83958 435922 84014 435978
rect 84082 435922 84138 435978
rect 114678 436294 114734 436350
rect 114802 436294 114858 436350
rect 114678 436170 114734 436226
rect 114802 436170 114858 436226
rect 114678 436046 114734 436102
rect 114802 436046 114858 436102
rect 114678 435922 114734 435978
rect 114802 435922 114858 435978
rect 145398 436294 145454 436350
rect 145522 436294 145578 436350
rect 145398 436170 145454 436226
rect 145522 436170 145578 436226
rect 145398 436046 145454 436102
rect 145522 436046 145578 436102
rect 145398 435922 145454 435978
rect 145522 435922 145578 435978
rect 176118 436294 176174 436350
rect 176242 436294 176298 436350
rect 176118 436170 176174 436226
rect 176242 436170 176298 436226
rect 176118 436046 176174 436102
rect 176242 436046 176298 436102
rect 176118 435922 176174 435978
rect 176242 435922 176298 435978
rect 206838 436294 206894 436350
rect 206962 436294 207018 436350
rect 206838 436170 206894 436226
rect 206962 436170 207018 436226
rect 206838 436046 206894 436102
rect 206962 436046 207018 436102
rect 206838 435922 206894 435978
rect 206962 435922 207018 435978
rect 237558 436294 237614 436350
rect 237682 436294 237738 436350
rect 237558 436170 237614 436226
rect 237682 436170 237738 436226
rect 237558 436046 237614 436102
rect 237682 436046 237738 436102
rect 237558 435922 237614 435978
rect 237682 435922 237738 435978
rect 268278 436294 268334 436350
rect 268402 436294 268458 436350
rect 268278 436170 268334 436226
rect 268402 436170 268458 436226
rect 268278 436046 268334 436102
rect 268402 436046 268458 436102
rect 268278 435922 268334 435978
rect 268402 435922 268458 435978
rect 298998 436294 299054 436350
rect 299122 436294 299178 436350
rect 298998 436170 299054 436226
rect 299122 436170 299178 436226
rect 298998 436046 299054 436102
rect 299122 436046 299178 436102
rect 298998 435922 299054 435978
rect 299122 435922 299178 435978
rect 329718 436294 329774 436350
rect 329842 436294 329898 436350
rect 329718 436170 329774 436226
rect 329842 436170 329898 436226
rect 329718 436046 329774 436102
rect 329842 436046 329898 436102
rect 329718 435922 329774 435978
rect 329842 435922 329898 435978
rect 360438 436294 360494 436350
rect 360562 436294 360618 436350
rect 360438 436170 360494 436226
rect 360562 436170 360618 436226
rect 360438 436046 360494 436102
rect 360562 436046 360618 436102
rect 360438 435922 360494 435978
rect 360562 435922 360618 435978
rect 391158 436294 391214 436350
rect 391282 436294 391338 436350
rect 391158 436170 391214 436226
rect 391282 436170 391338 436226
rect 391158 436046 391214 436102
rect 391282 436046 391338 436102
rect 391158 435922 391214 435978
rect 391282 435922 391338 435978
rect 421878 436294 421934 436350
rect 422002 436294 422058 436350
rect 421878 436170 421934 436226
rect 422002 436170 422058 436226
rect 421878 436046 421934 436102
rect 422002 436046 422058 436102
rect 421878 435922 421934 435978
rect 422002 435922 422058 435978
rect 452598 436294 452654 436350
rect 452722 436294 452778 436350
rect 452598 436170 452654 436226
rect 452722 436170 452778 436226
rect 452598 436046 452654 436102
rect 452722 436046 452778 436102
rect 452598 435922 452654 435978
rect 452722 435922 452778 435978
rect 483318 436294 483374 436350
rect 483442 436294 483498 436350
rect 483318 436170 483374 436226
rect 483442 436170 483498 436226
rect 483318 436046 483374 436102
rect 483442 436046 483498 436102
rect 483318 435922 483374 435978
rect 483442 435922 483498 435978
rect 514038 436294 514094 436350
rect 514162 436294 514218 436350
rect 514038 436170 514094 436226
rect 514162 436170 514218 436226
rect 514038 436046 514094 436102
rect 514162 436046 514218 436102
rect 514038 435922 514094 435978
rect 514162 435922 514218 435978
rect 544758 436294 544814 436350
rect 544882 436294 544938 436350
rect 544758 436170 544814 436226
rect 544882 436170 544938 436226
rect 544758 436046 544814 436102
rect 544882 436046 544938 436102
rect 544758 435922 544814 435978
rect 544882 435922 544938 435978
rect 37878 424294 37934 424350
rect 38002 424294 38058 424350
rect 37878 424170 37934 424226
rect 38002 424170 38058 424226
rect 37878 424046 37934 424102
rect 38002 424046 38058 424102
rect 37878 423922 37934 423978
rect 38002 423922 38058 423978
rect 68598 424294 68654 424350
rect 68722 424294 68778 424350
rect 68598 424170 68654 424226
rect 68722 424170 68778 424226
rect 68598 424046 68654 424102
rect 68722 424046 68778 424102
rect 68598 423922 68654 423978
rect 68722 423922 68778 423978
rect 99318 424294 99374 424350
rect 99442 424294 99498 424350
rect 99318 424170 99374 424226
rect 99442 424170 99498 424226
rect 99318 424046 99374 424102
rect 99442 424046 99498 424102
rect 99318 423922 99374 423978
rect 99442 423922 99498 423978
rect 130038 424294 130094 424350
rect 130162 424294 130218 424350
rect 130038 424170 130094 424226
rect 130162 424170 130218 424226
rect 130038 424046 130094 424102
rect 130162 424046 130218 424102
rect 130038 423922 130094 423978
rect 130162 423922 130218 423978
rect 160758 424294 160814 424350
rect 160882 424294 160938 424350
rect 160758 424170 160814 424226
rect 160882 424170 160938 424226
rect 160758 424046 160814 424102
rect 160882 424046 160938 424102
rect 160758 423922 160814 423978
rect 160882 423922 160938 423978
rect 191478 424294 191534 424350
rect 191602 424294 191658 424350
rect 191478 424170 191534 424226
rect 191602 424170 191658 424226
rect 191478 424046 191534 424102
rect 191602 424046 191658 424102
rect 191478 423922 191534 423978
rect 191602 423922 191658 423978
rect 222198 424294 222254 424350
rect 222322 424294 222378 424350
rect 222198 424170 222254 424226
rect 222322 424170 222378 424226
rect 222198 424046 222254 424102
rect 222322 424046 222378 424102
rect 222198 423922 222254 423978
rect 222322 423922 222378 423978
rect 252918 424294 252974 424350
rect 253042 424294 253098 424350
rect 252918 424170 252974 424226
rect 253042 424170 253098 424226
rect 252918 424046 252974 424102
rect 253042 424046 253098 424102
rect 252918 423922 252974 423978
rect 253042 423922 253098 423978
rect 283638 424294 283694 424350
rect 283762 424294 283818 424350
rect 283638 424170 283694 424226
rect 283762 424170 283818 424226
rect 283638 424046 283694 424102
rect 283762 424046 283818 424102
rect 283638 423922 283694 423978
rect 283762 423922 283818 423978
rect 314358 424294 314414 424350
rect 314482 424294 314538 424350
rect 314358 424170 314414 424226
rect 314482 424170 314538 424226
rect 314358 424046 314414 424102
rect 314482 424046 314538 424102
rect 314358 423922 314414 423978
rect 314482 423922 314538 423978
rect 345078 424294 345134 424350
rect 345202 424294 345258 424350
rect 345078 424170 345134 424226
rect 345202 424170 345258 424226
rect 345078 424046 345134 424102
rect 345202 424046 345258 424102
rect 345078 423922 345134 423978
rect 345202 423922 345258 423978
rect 375798 424294 375854 424350
rect 375922 424294 375978 424350
rect 375798 424170 375854 424226
rect 375922 424170 375978 424226
rect 375798 424046 375854 424102
rect 375922 424046 375978 424102
rect 375798 423922 375854 423978
rect 375922 423922 375978 423978
rect 406518 424294 406574 424350
rect 406642 424294 406698 424350
rect 406518 424170 406574 424226
rect 406642 424170 406698 424226
rect 406518 424046 406574 424102
rect 406642 424046 406698 424102
rect 406518 423922 406574 423978
rect 406642 423922 406698 423978
rect 437238 424294 437294 424350
rect 437362 424294 437418 424350
rect 437238 424170 437294 424226
rect 437362 424170 437418 424226
rect 437238 424046 437294 424102
rect 437362 424046 437418 424102
rect 437238 423922 437294 423978
rect 437362 423922 437418 423978
rect 467958 424294 468014 424350
rect 468082 424294 468138 424350
rect 467958 424170 468014 424226
rect 468082 424170 468138 424226
rect 467958 424046 468014 424102
rect 468082 424046 468138 424102
rect 467958 423922 468014 423978
rect 468082 423922 468138 423978
rect 498678 424294 498734 424350
rect 498802 424294 498858 424350
rect 498678 424170 498734 424226
rect 498802 424170 498858 424226
rect 498678 424046 498734 424102
rect 498802 424046 498858 424102
rect 498678 423922 498734 423978
rect 498802 423922 498858 423978
rect 529398 424294 529454 424350
rect 529522 424294 529578 424350
rect 529398 424170 529454 424226
rect 529522 424170 529578 424226
rect 529398 424046 529454 424102
rect 529522 424046 529578 424102
rect 529398 423922 529454 423978
rect 529522 423922 529578 423978
rect 53238 418294 53294 418350
rect 53362 418294 53418 418350
rect 53238 418170 53294 418226
rect 53362 418170 53418 418226
rect 53238 418046 53294 418102
rect 53362 418046 53418 418102
rect 53238 417922 53294 417978
rect 53362 417922 53418 417978
rect 83958 418294 84014 418350
rect 84082 418294 84138 418350
rect 83958 418170 84014 418226
rect 84082 418170 84138 418226
rect 83958 418046 84014 418102
rect 84082 418046 84138 418102
rect 83958 417922 84014 417978
rect 84082 417922 84138 417978
rect 114678 418294 114734 418350
rect 114802 418294 114858 418350
rect 114678 418170 114734 418226
rect 114802 418170 114858 418226
rect 114678 418046 114734 418102
rect 114802 418046 114858 418102
rect 114678 417922 114734 417978
rect 114802 417922 114858 417978
rect 145398 418294 145454 418350
rect 145522 418294 145578 418350
rect 145398 418170 145454 418226
rect 145522 418170 145578 418226
rect 145398 418046 145454 418102
rect 145522 418046 145578 418102
rect 145398 417922 145454 417978
rect 145522 417922 145578 417978
rect 176118 418294 176174 418350
rect 176242 418294 176298 418350
rect 176118 418170 176174 418226
rect 176242 418170 176298 418226
rect 176118 418046 176174 418102
rect 176242 418046 176298 418102
rect 176118 417922 176174 417978
rect 176242 417922 176298 417978
rect 206838 418294 206894 418350
rect 206962 418294 207018 418350
rect 206838 418170 206894 418226
rect 206962 418170 207018 418226
rect 206838 418046 206894 418102
rect 206962 418046 207018 418102
rect 206838 417922 206894 417978
rect 206962 417922 207018 417978
rect 237558 418294 237614 418350
rect 237682 418294 237738 418350
rect 237558 418170 237614 418226
rect 237682 418170 237738 418226
rect 237558 418046 237614 418102
rect 237682 418046 237738 418102
rect 237558 417922 237614 417978
rect 237682 417922 237738 417978
rect 268278 418294 268334 418350
rect 268402 418294 268458 418350
rect 268278 418170 268334 418226
rect 268402 418170 268458 418226
rect 268278 418046 268334 418102
rect 268402 418046 268458 418102
rect 268278 417922 268334 417978
rect 268402 417922 268458 417978
rect 298998 418294 299054 418350
rect 299122 418294 299178 418350
rect 298998 418170 299054 418226
rect 299122 418170 299178 418226
rect 298998 418046 299054 418102
rect 299122 418046 299178 418102
rect 298998 417922 299054 417978
rect 299122 417922 299178 417978
rect 329718 418294 329774 418350
rect 329842 418294 329898 418350
rect 329718 418170 329774 418226
rect 329842 418170 329898 418226
rect 329718 418046 329774 418102
rect 329842 418046 329898 418102
rect 329718 417922 329774 417978
rect 329842 417922 329898 417978
rect 360438 418294 360494 418350
rect 360562 418294 360618 418350
rect 360438 418170 360494 418226
rect 360562 418170 360618 418226
rect 360438 418046 360494 418102
rect 360562 418046 360618 418102
rect 360438 417922 360494 417978
rect 360562 417922 360618 417978
rect 391158 418294 391214 418350
rect 391282 418294 391338 418350
rect 391158 418170 391214 418226
rect 391282 418170 391338 418226
rect 391158 418046 391214 418102
rect 391282 418046 391338 418102
rect 391158 417922 391214 417978
rect 391282 417922 391338 417978
rect 421878 418294 421934 418350
rect 422002 418294 422058 418350
rect 421878 418170 421934 418226
rect 422002 418170 422058 418226
rect 421878 418046 421934 418102
rect 422002 418046 422058 418102
rect 421878 417922 421934 417978
rect 422002 417922 422058 417978
rect 452598 418294 452654 418350
rect 452722 418294 452778 418350
rect 452598 418170 452654 418226
rect 452722 418170 452778 418226
rect 452598 418046 452654 418102
rect 452722 418046 452778 418102
rect 452598 417922 452654 417978
rect 452722 417922 452778 417978
rect 483318 418294 483374 418350
rect 483442 418294 483498 418350
rect 483318 418170 483374 418226
rect 483442 418170 483498 418226
rect 483318 418046 483374 418102
rect 483442 418046 483498 418102
rect 483318 417922 483374 417978
rect 483442 417922 483498 417978
rect 514038 418294 514094 418350
rect 514162 418294 514218 418350
rect 514038 418170 514094 418226
rect 514162 418170 514218 418226
rect 514038 418046 514094 418102
rect 514162 418046 514218 418102
rect 514038 417922 514094 417978
rect 514162 417922 514218 417978
rect 544758 418294 544814 418350
rect 544882 418294 544938 418350
rect 544758 418170 544814 418226
rect 544882 418170 544938 418226
rect 544758 418046 544814 418102
rect 544882 418046 544938 418102
rect 544758 417922 544814 417978
rect 544882 417922 544938 417978
rect 37878 406294 37934 406350
rect 38002 406294 38058 406350
rect 37878 406170 37934 406226
rect 38002 406170 38058 406226
rect 37878 406046 37934 406102
rect 38002 406046 38058 406102
rect 37878 405922 37934 405978
rect 38002 405922 38058 405978
rect 68598 406294 68654 406350
rect 68722 406294 68778 406350
rect 68598 406170 68654 406226
rect 68722 406170 68778 406226
rect 68598 406046 68654 406102
rect 68722 406046 68778 406102
rect 68598 405922 68654 405978
rect 68722 405922 68778 405978
rect 99318 406294 99374 406350
rect 99442 406294 99498 406350
rect 99318 406170 99374 406226
rect 99442 406170 99498 406226
rect 99318 406046 99374 406102
rect 99442 406046 99498 406102
rect 99318 405922 99374 405978
rect 99442 405922 99498 405978
rect 130038 406294 130094 406350
rect 130162 406294 130218 406350
rect 130038 406170 130094 406226
rect 130162 406170 130218 406226
rect 130038 406046 130094 406102
rect 130162 406046 130218 406102
rect 130038 405922 130094 405978
rect 130162 405922 130218 405978
rect 160758 406294 160814 406350
rect 160882 406294 160938 406350
rect 160758 406170 160814 406226
rect 160882 406170 160938 406226
rect 160758 406046 160814 406102
rect 160882 406046 160938 406102
rect 160758 405922 160814 405978
rect 160882 405922 160938 405978
rect 191478 406294 191534 406350
rect 191602 406294 191658 406350
rect 191478 406170 191534 406226
rect 191602 406170 191658 406226
rect 191478 406046 191534 406102
rect 191602 406046 191658 406102
rect 191478 405922 191534 405978
rect 191602 405922 191658 405978
rect 222198 406294 222254 406350
rect 222322 406294 222378 406350
rect 222198 406170 222254 406226
rect 222322 406170 222378 406226
rect 222198 406046 222254 406102
rect 222322 406046 222378 406102
rect 222198 405922 222254 405978
rect 222322 405922 222378 405978
rect 252918 406294 252974 406350
rect 253042 406294 253098 406350
rect 252918 406170 252974 406226
rect 253042 406170 253098 406226
rect 252918 406046 252974 406102
rect 253042 406046 253098 406102
rect 252918 405922 252974 405978
rect 253042 405922 253098 405978
rect 283638 406294 283694 406350
rect 283762 406294 283818 406350
rect 283638 406170 283694 406226
rect 283762 406170 283818 406226
rect 283638 406046 283694 406102
rect 283762 406046 283818 406102
rect 283638 405922 283694 405978
rect 283762 405922 283818 405978
rect 314358 406294 314414 406350
rect 314482 406294 314538 406350
rect 314358 406170 314414 406226
rect 314482 406170 314538 406226
rect 314358 406046 314414 406102
rect 314482 406046 314538 406102
rect 314358 405922 314414 405978
rect 314482 405922 314538 405978
rect 345078 406294 345134 406350
rect 345202 406294 345258 406350
rect 345078 406170 345134 406226
rect 345202 406170 345258 406226
rect 345078 406046 345134 406102
rect 345202 406046 345258 406102
rect 345078 405922 345134 405978
rect 345202 405922 345258 405978
rect 375798 406294 375854 406350
rect 375922 406294 375978 406350
rect 375798 406170 375854 406226
rect 375922 406170 375978 406226
rect 375798 406046 375854 406102
rect 375922 406046 375978 406102
rect 375798 405922 375854 405978
rect 375922 405922 375978 405978
rect 406518 406294 406574 406350
rect 406642 406294 406698 406350
rect 406518 406170 406574 406226
rect 406642 406170 406698 406226
rect 406518 406046 406574 406102
rect 406642 406046 406698 406102
rect 406518 405922 406574 405978
rect 406642 405922 406698 405978
rect 437238 406294 437294 406350
rect 437362 406294 437418 406350
rect 437238 406170 437294 406226
rect 437362 406170 437418 406226
rect 437238 406046 437294 406102
rect 437362 406046 437418 406102
rect 437238 405922 437294 405978
rect 437362 405922 437418 405978
rect 467958 406294 468014 406350
rect 468082 406294 468138 406350
rect 467958 406170 468014 406226
rect 468082 406170 468138 406226
rect 467958 406046 468014 406102
rect 468082 406046 468138 406102
rect 467958 405922 468014 405978
rect 468082 405922 468138 405978
rect 498678 406294 498734 406350
rect 498802 406294 498858 406350
rect 498678 406170 498734 406226
rect 498802 406170 498858 406226
rect 498678 406046 498734 406102
rect 498802 406046 498858 406102
rect 498678 405922 498734 405978
rect 498802 405922 498858 405978
rect 529398 406294 529454 406350
rect 529522 406294 529578 406350
rect 529398 406170 529454 406226
rect 529522 406170 529578 406226
rect 529398 406046 529454 406102
rect 529522 406046 529578 406102
rect 529398 405922 529454 405978
rect 529522 405922 529578 405978
rect 53238 400294 53294 400350
rect 53362 400294 53418 400350
rect 53238 400170 53294 400226
rect 53362 400170 53418 400226
rect 53238 400046 53294 400102
rect 53362 400046 53418 400102
rect 53238 399922 53294 399978
rect 53362 399922 53418 399978
rect 83958 400294 84014 400350
rect 84082 400294 84138 400350
rect 83958 400170 84014 400226
rect 84082 400170 84138 400226
rect 83958 400046 84014 400102
rect 84082 400046 84138 400102
rect 83958 399922 84014 399978
rect 84082 399922 84138 399978
rect 114678 400294 114734 400350
rect 114802 400294 114858 400350
rect 114678 400170 114734 400226
rect 114802 400170 114858 400226
rect 114678 400046 114734 400102
rect 114802 400046 114858 400102
rect 114678 399922 114734 399978
rect 114802 399922 114858 399978
rect 145398 400294 145454 400350
rect 145522 400294 145578 400350
rect 145398 400170 145454 400226
rect 145522 400170 145578 400226
rect 145398 400046 145454 400102
rect 145522 400046 145578 400102
rect 145398 399922 145454 399978
rect 145522 399922 145578 399978
rect 176118 400294 176174 400350
rect 176242 400294 176298 400350
rect 176118 400170 176174 400226
rect 176242 400170 176298 400226
rect 176118 400046 176174 400102
rect 176242 400046 176298 400102
rect 176118 399922 176174 399978
rect 176242 399922 176298 399978
rect 206838 400294 206894 400350
rect 206962 400294 207018 400350
rect 206838 400170 206894 400226
rect 206962 400170 207018 400226
rect 206838 400046 206894 400102
rect 206962 400046 207018 400102
rect 206838 399922 206894 399978
rect 206962 399922 207018 399978
rect 237558 400294 237614 400350
rect 237682 400294 237738 400350
rect 237558 400170 237614 400226
rect 237682 400170 237738 400226
rect 237558 400046 237614 400102
rect 237682 400046 237738 400102
rect 237558 399922 237614 399978
rect 237682 399922 237738 399978
rect 268278 400294 268334 400350
rect 268402 400294 268458 400350
rect 268278 400170 268334 400226
rect 268402 400170 268458 400226
rect 268278 400046 268334 400102
rect 268402 400046 268458 400102
rect 268278 399922 268334 399978
rect 268402 399922 268458 399978
rect 298998 400294 299054 400350
rect 299122 400294 299178 400350
rect 298998 400170 299054 400226
rect 299122 400170 299178 400226
rect 298998 400046 299054 400102
rect 299122 400046 299178 400102
rect 298998 399922 299054 399978
rect 299122 399922 299178 399978
rect 329718 400294 329774 400350
rect 329842 400294 329898 400350
rect 329718 400170 329774 400226
rect 329842 400170 329898 400226
rect 329718 400046 329774 400102
rect 329842 400046 329898 400102
rect 329718 399922 329774 399978
rect 329842 399922 329898 399978
rect 360438 400294 360494 400350
rect 360562 400294 360618 400350
rect 360438 400170 360494 400226
rect 360562 400170 360618 400226
rect 360438 400046 360494 400102
rect 360562 400046 360618 400102
rect 360438 399922 360494 399978
rect 360562 399922 360618 399978
rect 391158 400294 391214 400350
rect 391282 400294 391338 400350
rect 391158 400170 391214 400226
rect 391282 400170 391338 400226
rect 391158 400046 391214 400102
rect 391282 400046 391338 400102
rect 391158 399922 391214 399978
rect 391282 399922 391338 399978
rect 421878 400294 421934 400350
rect 422002 400294 422058 400350
rect 421878 400170 421934 400226
rect 422002 400170 422058 400226
rect 421878 400046 421934 400102
rect 422002 400046 422058 400102
rect 421878 399922 421934 399978
rect 422002 399922 422058 399978
rect 452598 400294 452654 400350
rect 452722 400294 452778 400350
rect 452598 400170 452654 400226
rect 452722 400170 452778 400226
rect 452598 400046 452654 400102
rect 452722 400046 452778 400102
rect 452598 399922 452654 399978
rect 452722 399922 452778 399978
rect 483318 400294 483374 400350
rect 483442 400294 483498 400350
rect 483318 400170 483374 400226
rect 483442 400170 483498 400226
rect 483318 400046 483374 400102
rect 483442 400046 483498 400102
rect 483318 399922 483374 399978
rect 483442 399922 483498 399978
rect 514038 400294 514094 400350
rect 514162 400294 514218 400350
rect 514038 400170 514094 400226
rect 514162 400170 514218 400226
rect 514038 400046 514094 400102
rect 514162 400046 514218 400102
rect 514038 399922 514094 399978
rect 514162 399922 514218 399978
rect 544758 400294 544814 400350
rect 544882 400294 544938 400350
rect 544758 400170 544814 400226
rect 544882 400170 544938 400226
rect 544758 400046 544814 400102
rect 544882 400046 544938 400102
rect 544758 399922 544814 399978
rect 544882 399922 544938 399978
rect 37782 370294 37838 370350
rect 37906 370294 37962 370350
rect 37782 370170 37838 370226
rect 37906 370170 37962 370226
rect 37782 370046 37838 370102
rect 37906 370046 37962 370102
rect 37782 369922 37838 369978
rect 37906 369922 37962 369978
rect 68502 370294 68558 370350
rect 68626 370294 68682 370350
rect 68502 370170 68558 370226
rect 68626 370170 68682 370226
rect 68502 370046 68558 370102
rect 68626 370046 68682 370102
rect 68502 369922 68558 369978
rect 68626 369922 68682 369978
rect 99222 370294 99278 370350
rect 99346 370294 99402 370350
rect 99222 370170 99278 370226
rect 99346 370170 99402 370226
rect 99222 370046 99278 370102
rect 99346 370046 99402 370102
rect 99222 369922 99278 369978
rect 99346 369922 99402 369978
rect 129942 370294 129998 370350
rect 130066 370294 130122 370350
rect 129942 370170 129998 370226
rect 130066 370170 130122 370226
rect 129942 370046 129998 370102
rect 130066 370046 130122 370102
rect 129942 369922 129998 369978
rect 130066 369922 130122 369978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect 22422 364294 22478 364350
rect 22546 364294 22602 364350
rect 22422 364170 22478 364226
rect 22546 364170 22602 364226
rect 22422 364046 22478 364102
rect 22546 364046 22602 364102
rect 22422 363922 22478 363978
rect 22546 363922 22602 363978
rect 53142 364294 53198 364350
rect 53266 364294 53322 364350
rect 53142 364170 53198 364226
rect 53266 364170 53322 364226
rect 53142 364046 53198 364102
rect 53266 364046 53322 364102
rect 53142 363922 53198 363978
rect 53266 363922 53322 363978
rect 83862 364294 83918 364350
rect 83986 364294 84042 364350
rect 83862 364170 83918 364226
rect 83986 364170 84042 364226
rect 83862 364046 83918 364102
rect 83986 364046 84042 364102
rect 83862 363922 83918 363978
rect 83986 363922 84042 363978
rect 114582 364294 114638 364350
rect 114706 364294 114762 364350
rect 114582 364170 114638 364226
rect 114706 364170 114762 364226
rect 114582 364046 114638 364102
rect 114706 364046 114762 364102
rect 114582 363922 114638 363978
rect 114706 363922 114762 363978
rect 145302 364294 145358 364350
rect 145426 364294 145482 364350
rect 145302 364170 145358 364226
rect 145426 364170 145482 364226
rect 145302 364046 145358 364102
rect 145426 364046 145482 364102
rect 145302 363922 145358 363978
rect 145426 363922 145482 363978
rect 37782 352294 37838 352350
rect 37906 352294 37962 352350
rect 37782 352170 37838 352226
rect 37906 352170 37962 352226
rect 37782 352046 37838 352102
rect 37906 352046 37962 352102
rect 37782 351922 37838 351978
rect 37906 351922 37962 351978
rect 68502 352294 68558 352350
rect 68626 352294 68682 352350
rect 68502 352170 68558 352226
rect 68626 352170 68682 352226
rect 68502 352046 68558 352102
rect 68626 352046 68682 352102
rect 68502 351922 68558 351978
rect 68626 351922 68682 351978
rect 99222 352294 99278 352350
rect 99346 352294 99402 352350
rect 99222 352170 99278 352226
rect 99346 352170 99402 352226
rect 99222 352046 99278 352102
rect 99346 352046 99402 352102
rect 99222 351922 99278 351978
rect 99346 351922 99402 351978
rect 129942 352294 129998 352350
rect 130066 352294 130122 352350
rect 129942 352170 129998 352226
rect 130066 352170 130122 352226
rect 129942 352046 129998 352102
rect 130066 352046 130122 352102
rect 129942 351922 129998 351978
rect 130066 351922 130122 351978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 22422 346294 22478 346350
rect 22546 346294 22602 346350
rect 22422 346170 22478 346226
rect 22546 346170 22602 346226
rect 22422 346046 22478 346102
rect 22546 346046 22602 346102
rect 22422 345922 22478 345978
rect 22546 345922 22602 345978
rect 53142 346294 53198 346350
rect 53266 346294 53322 346350
rect 53142 346170 53198 346226
rect 53266 346170 53322 346226
rect 53142 346046 53198 346102
rect 53266 346046 53322 346102
rect 53142 345922 53198 345978
rect 53266 345922 53322 345978
rect 83862 346294 83918 346350
rect 83986 346294 84042 346350
rect 83862 346170 83918 346226
rect 83986 346170 84042 346226
rect 83862 346046 83918 346102
rect 83986 346046 84042 346102
rect 83862 345922 83918 345978
rect 83986 345922 84042 345978
rect 114582 346294 114638 346350
rect 114706 346294 114762 346350
rect 114582 346170 114638 346226
rect 114706 346170 114762 346226
rect 114582 346046 114638 346102
rect 114706 346046 114762 346102
rect 114582 345922 114638 345978
rect 114706 345922 114762 345978
rect 145302 346294 145358 346350
rect 145426 346294 145482 346350
rect 145302 346170 145358 346226
rect 145426 346170 145482 346226
rect 145302 346046 145358 346102
rect 145426 346046 145482 346102
rect 145302 345922 145358 345978
rect 145426 345922 145482 345978
rect 37782 334294 37838 334350
rect 37906 334294 37962 334350
rect 37782 334170 37838 334226
rect 37906 334170 37962 334226
rect 37782 334046 37838 334102
rect 37906 334046 37962 334102
rect 37782 333922 37838 333978
rect 37906 333922 37962 333978
rect 68502 334294 68558 334350
rect 68626 334294 68682 334350
rect 68502 334170 68558 334226
rect 68626 334170 68682 334226
rect 68502 334046 68558 334102
rect 68626 334046 68682 334102
rect 68502 333922 68558 333978
rect 68626 333922 68682 333978
rect 99222 334294 99278 334350
rect 99346 334294 99402 334350
rect 99222 334170 99278 334226
rect 99346 334170 99402 334226
rect 99222 334046 99278 334102
rect 99346 334046 99402 334102
rect 99222 333922 99278 333978
rect 99346 333922 99402 333978
rect 129942 334294 129998 334350
rect 130066 334294 130122 334350
rect 129942 334170 129998 334226
rect 130066 334170 130122 334226
rect 129942 334046 129998 334102
rect 130066 334046 130122 334102
rect 129942 333922 129998 333978
rect 130066 333922 130122 333978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 4172 16622 4228 16678
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 22422 328294 22478 328350
rect 22546 328294 22602 328350
rect 22422 328170 22478 328226
rect 22546 328170 22602 328226
rect 22422 328046 22478 328102
rect 22546 328046 22602 328102
rect 22422 327922 22478 327978
rect 22546 327922 22602 327978
rect 53142 328294 53198 328350
rect 53266 328294 53322 328350
rect 53142 328170 53198 328226
rect 53266 328170 53322 328226
rect 53142 328046 53198 328102
rect 53266 328046 53322 328102
rect 53142 327922 53198 327978
rect 53266 327922 53322 327978
rect 83862 328294 83918 328350
rect 83986 328294 84042 328350
rect 83862 328170 83918 328226
rect 83986 328170 84042 328226
rect 83862 328046 83918 328102
rect 83986 328046 84042 328102
rect 83862 327922 83918 327978
rect 83986 327922 84042 327978
rect 114582 328294 114638 328350
rect 114706 328294 114762 328350
rect 114582 328170 114638 328226
rect 114706 328170 114762 328226
rect 114582 328046 114638 328102
rect 114706 328046 114762 328102
rect 114582 327922 114638 327978
rect 114706 327922 114762 327978
rect 145302 328294 145358 328350
rect 145426 328294 145482 328350
rect 145302 328170 145358 328226
rect 145426 328170 145482 328226
rect 145302 328046 145358 328102
rect 145426 328046 145482 328102
rect 145302 327922 145358 327978
rect 145426 327922 145482 327978
rect 37782 316294 37838 316350
rect 37906 316294 37962 316350
rect 37782 316170 37838 316226
rect 37906 316170 37962 316226
rect 37782 316046 37838 316102
rect 37906 316046 37962 316102
rect 37782 315922 37838 315978
rect 37906 315922 37962 315978
rect 68502 316294 68558 316350
rect 68626 316294 68682 316350
rect 68502 316170 68558 316226
rect 68626 316170 68682 316226
rect 68502 316046 68558 316102
rect 68626 316046 68682 316102
rect 68502 315922 68558 315978
rect 68626 315922 68682 315978
rect 99222 316294 99278 316350
rect 99346 316294 99402 316350
rect 99222 316170 99278 316226
rect 99346 316170 99402 316226
rect 99222 316046 99278 316102
rect 99346 316046 99402 316102
rect 99222 315922 99278 315978
rect 99346 315922 99402 315978
rect 129942 316294 129998 316350
rect 130066 316294 130122 316350
rect 129942 316170 129998 316226
rect 130066 316170 130122 316226
rect 129942 316046 129998 316102
rect 130066 316046 130122 316102
rect 129942 315922 129998 315978
rect 130066 315922 130122 315978
rect 22422 310294 22478 310350
rect 22546 310294 22602 310350
rect 22422 310170 22478 310226
rect 22546 310170 22602 310226
rect 22422 310046 22478 310102
rect 22546 310046 22602 310102
rect 22422 309922 22478 309978
rect 22546 309922 22602 309978
rect 53142 310294 53198 310350
rect 53266 310294 53322 310350
rect 53142 310170 53198 310226
rect 53266 310170 53322 310226
rect 53142 310046 53198 310102
rect 53266 310046 53322 310102
rect 53142 309922 53198 309978
rect 53266 309922 53322 309978
rect 83862 310294 83918 310350
rect 83986 310294 84042 310350
rect 83862 310170 83918 310226
rect 83986 310170 84042 310226
rect 83862 310046 83918 310102
rect 83986 310046 84042 310102
rect 83862 309922 83918 309978
rect 83986 309922 84042 309978
rect 114582 310294 114638 310350
rect 114706 310294 114762 310350
rect 114582 310170 114638 310226
rect 114706 310170 114762 310226
rect 114582 310046 114638 310102
rect 114706 310046 114762 310102
rect 114582 309922 114638 309978
rect 114706 309922 114762 309978
rect 145302 310294 145358 310350
rect 145426 310294 145482 310350
rect 145302 310170 145358 310226
rect 145426 310170 145482 310226
rect 145302 310046 145358 310102
rect 145426 310046 145482 310102
rect 145302 309922 145358 309978
rect 145426 309922 145482 309978
rect 37782 298294 37838 298350
rect 37906 298294 37962 298350
rect 37782 298170 37838 298226
rect 37906 298170 37962 298226
rect 37782 298046 37838 298102
rect 37906 298046 37962 298102
rect 37782 297922 37838 297978
rect 37906 297922 37962 297978
rect 68502 298294 68558 298350
rect 68626 298294 68682 298350
rect 68502 298170 68558 298226
rect 68626 298170 68682 298226
rect 68502 298046 68558 298102
rect 68626 298046 68682 298102
rect 68502 297922 68558 297978
rect 68626 297922 68682 297978
rect 99222 298294 99278 298350
rect 99346 298294 99402 298350
rect 99222 298170 99278 298226
rect 99346 298170 99402 298226
rect 99222 298046 99278 298102
rect 99346 298046 99402 298102
rect 99222 297922 99278 297978
rect 99346 297922 99402 297978
rect 129942 298294 129998 298350
rect 130066 298294 130122 298350
rect 129942 298170 129998 298226
rect 130066 298170 130122 298226
rect 129942 298046 129998 298102
rect 130066 298046 130122 298102
rect 129942 297922 129998 297978
rect 130066 297922 130122 297978
rect 22422 292294 22478 292350
rect 22546 292294 22602 292350
rect 22422 292170 22478 292226
rect 22546 292170 22602 292226
rect 22422 292046 22478 292102
rect 22546 292046 22602 292102
rect 22422 291922 22478 291978
rect 22546 291922 22602 291978
rect 53142 292294 53198 292350
rect 53266 292294 53322 292350
rect 53142 292170 53198 292226
rect 53266 292170 53322 292226
rect 53142 292046 53198 292102
rect 53266 292046 53322 292102
rect 53142 291922 53198 291978
rect 53266 291922 53322 291978
rect 83862 292294 83918 292350
rect 83986 292294 84042 292350
rect 83862 292170 83918 292226
rect 83986 292170 84042 292226
rect 83862 292046 83918 292102
rect 83986 292046 84042 292102
rect 83862 291922 83918 291978
rect 83986 291922 84042 291978
rect 114582 292294 114638 292350
rect 114706 292294 114762 292350
rect 114582 292170 114638 292226
rect 114706 292170 114762 292226
rect 114582 292046 114638 292102
rect 114706 292046 114762 292102
rect 114582 291922 114638 291978
rect 114706 291922 114762 291978
rect 145302 292294 145358 292350
rect 145426 292294 145482 292350
rect 145302 292170 145358 292226
rect 145426 292170 145482 292226
rect 145302 292046 145358 292102
rect 145426 292046 145482 292102
rect 145302 291922 145358 291978
rect 145426 291922 145482 291978
rect 37782 280294 37838 280350
rect 37906 280294 37962 280350
rect 37782 280170 37838 280226
rect 37906 280170 37962 280226
rect 37782 280046 37838 280102
rect 37906 280046 37962 280102
rect 37782 279922 37838 279978
rect 37906 279922 37962 279978
rect 68502 280294 68558 280350
rect 68626 280294 68682 280350
rect 68502 280170 68558 280226
rect 68626 280170 68682 280226
rect 68502 280046 68558 280102
rect 68626 280046 68682 280102
rect 68502 279922 68558 279978
rect 68626 279922 68682 279978
rect 99222 280294 99278 280350
rect 99346 280294 99402 280350
rect 99222 280170 99278 280226
rect 99346 280170 99402 280226
rect 99222 280046 99278 280102
rect 99346 280046 99402 280102
rect 99222 279922 99278 279978
rect 99346 279922 99402 279978
rect 129942 280294 129998 280350
rect 130066 280294 130122 280350
rect 129942 280170 129998 280226
rect 130066 280170 130122 280226
rect 129942 280046 129998 280102
rect 130066 280046 130122 280102
rect 129942 279922 129998 279978
rect 130066 279922 130122 279978
rect 22422 274294 22478 274350
rect 22546 274294 22602 274350
rect 22422 274170 22478 274226
rect 22546 274170 22602 274226
rect 22422 274046 22478 274102
rect 22546 274046 22602 274102
rect 22422 273922 22478 273978
rect 22546 273922 22602 273978
rect 53142 274294 53198 274350
rect 53266 274294 53322 274350
rect 53142 274170 53198 274226
rect 53266 274170 53322 274226
rect 53142 274046 53198 274102
rect 53266 274046 53322 274102
rect 53142 273922 53198 273978
rect 53266 273922 53322 273978
rect 83862 274294 83918 274350
rect 83986 274294 84042 274350
rect 83862 274170 83918 274226
rect 83986 274170 84042 274226
rect 83862 274046 83918 274102
rect 83986 274046 84042 274102
rect 83862 273922 83918 273978
rect 83986 273922 84042 273978
rect 114582 274294 114638 274350
rect 114706 274294 114762 274350
rect 114582 274170 114638 274226
rect 114706 274170 114762 274226
rect 114582 274046 114638 274102
rect 114706 274046 114762 274102
rect 114582 273922 114638 273978
rect 114706 273922 114762 273978
rect 145302 274294 145358 274350
rect 145426 274294 145482 274350
rect 145302 274170 145358 274226
rect 145426 274170 145482 274226
rect 145302 274046 145358 274102
rect 145426 274046 145482 274102
rect 145302 273922 145358 273978
rect 145426 273922 145482 273978
rect 37782 262294 37838 262350
rect 37906 262294 37962 262350
rect 37782 262170 37838 262226
rect 37906 262170 37962 262226
rect 37782 262046 37838 262102
rect 37906 262046 37962 262102
rect 37782 261922 37838 261978
rect 37906 261922 37962 261978
rect 68502 262294 68558 262350
rect 68626 262294 68682 262350
rect 68502 262170 68558 262226
rect 68626 262170 68682 262226
rect 68502 262046 68558 262102
rect 68626 262046 68682 262102
rect 68502 261922 68558 261978
rect 68626 261922 68682 261978
rect 99222 262294 99278 262350
rect 99346 262294 99402 262350
rect 99222 262170 99278 262226
rect 99346 262170 99402 262226
rect 99222 262046 99278 262102
rect 99346 262046 99402 262102
rect 99222 261922 99278 261978
rect 99346 261922 99402 261978
rect 129942 262294 129998 262350
rect 130066 262294 130122 262350
rect 129942 262170 129998 262226
rect 130066 262170 130122 262226
rect 129942 262046 129998 262102
rect 130066 262046 130122 262102
rect 129942 261922 129998 261978
rect 130066 261922 130122 261978
rect 22422 256294 22478 256350
rect 22546 256294 22602 256350
rect 22422 256170 22478 256226
rect 22546 256170 22602 256226
rect 22422 256046 22478 256102
rect 22546 256046 22602 256102
rect 22422 255922 22478 255978
rect 22546 255922 22602 255978
rect 53142 256294 53198 256350
rect 53266 256294 53322 256350
rect 53142 256170 53198 256226
rect 53266 256170 53322 256226
rect 53142 256046 53198 256102
rect 53266 256046 53322 256102
rect 53142 255922 53198 255978
rect 53266 255922 53322 255978
rect 83862 256294 83918 256350
rect 83986 256294 84042 256350
rect 83862 256170 83918 256226
rect 83986 256170 84042 256226
rect 83862 256046 83918 256102
rect 83986 256046 84042 256102
rect 83862 255922 83918 255978
rect 83986 255922 84042 255978
rect 114582 256294 114638 256350
rect 114706 256294 114762 256350
rect 114582 256170 114638 256226
rect 114706 256170 114762 256226
rect 114582 256046 114638 256102
rect 114706 256046 114762 256102
rect 114582 255922 114638 255978
rect 114706 255922 114762 255978
rect 145302 256294 145358 256350
rect 145426 256294 145482 256350
rect 145302 256170 145358 256226
rect 145426 256170 145482 256226
rect 145302 256046 145358 256102
rect 145426 256046 145482 256102
rect 145302 255922 145358 255978
rect 145426 255922 145482 255978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 37782 244294 37838 244350
rect 37906 244294 37962 244350
rect 37782 244170 37838 244226
rect 37906 244170 37962 244226
rect 37782 244046 37838 244102
rect 37906 244046 37962 244102
rect 37782 243922 37838 243978
rect 37906 243922 37962 243978
rect 68502 244294 68558 244350
rect 68626 244294 68682 244350
rect 68502 244170 68558 244226
rect 68626 244170 68682 244226
rect 68502 244046 68558 244102
rect 68626 244046 68682 244102
rect 68502 243922 68558 243978
rect 68626 243922 68682 243978
rect 99222 244294 99278 244350
rect 99346 244294 99402 244350
rect 99222 244170 99278 244226
rect 99346 244170 99402 244226
rect 99222 244046 99278 244102
rect 99346 244046 99402 244102
rect 99222 243922 99278 243978
rect 99346 243922 99402 243978
rect 129942 244294 129998 244350
rect 130066 244294 130122 244350
rect 129942 244170 129998 244226
rect 130066 244170 130122 244226
rect 129942 244046 129998 244102
rect 130066 244046 130122 244102
rect 129942 243922 129998 243978
rect 130066 243922 130122 243978
rect 22422 238294 22478 238350
rect 22546 238294 22602 238350
rect 22422 238170 22478 238226
rect 22546 238170 22602 238226
rect 22422 238046 22478 238102
rect 22546 238046 22602 238102
rect 22422 237922 22478 237978
rect 22546 237922 22602 237978
rect 53142 238294 53198 238350
rect 53266 238294 53322 238350
rect 53142 238170 53198 238226
rect 53266 238170 53322 238226
rect 53142 238046 53198 238102
rect 53266 238046 53322 238102
rect 53142 237922 53198 237978
rect 53266 237922 53322 237978
rect 83862 238294 83918 238350
rect 83986 238294 84042 238350
rect 83862 238170 83918 238226
rect 83986 238170 84042 238226
rect 83862 238046 83918 238102
rect 83986 238046 84042 238102
rect 83862 237922 83918 237978
rect 83986 237922 84042 237978
rect 114582 238294 114638 238350
rect 114706 238294 114762 238350
rect 114582 238170 114638 238226
rect 114706 238170 114762 238226
rect 114582 238046 114638 238102
rect 114706 238046 114762 238102
rect 114582 237922 114638 237978
rect 114706 237922 114762 237978
rect 145302 238294 145358 238350
rect 145426 238294 145482 238350
rect 145302 238170 145358 238226
rect 145426 238170 145482 238226
rect 145302 238046 145358 238102
rect 145426 238046 145482 238102
rect 145302 237922 145358 237978
rect 145426 237922 145482 237978
rect 37782 226294 37838 226350
rect 37906 226294 37962 226350
rect 37782 226170 37838 226226
rect 37906 226170 37962 226226
rect 37782 226046 37838 226102
rect 37906 226046 37962 226102
rect 37782 225922 37838 225978
rect 37906 225922 37962 225978
rect 68502 226294 68558 226350
rect 68626 226294 68682 226350
rect 68502 226170 68558 226226
rect 68626 226170 68682 226226
rect 68502 226046 68558 226102
rect 68626 226046 68682 226102
rect 68502 225922 68558 225978
rect 68626 225922 68682 225978
rect 99222 226294 99278 226350
rect 99346 226294 99402 226350
rect 99222 226170 99278 226226
rect 99346 226170 99402 226226
rect 99222 226046 99278 226102
rect 99346 226046 99402 226102
rect 99222 225922 99278 225978
rect 99346 225922 99402 225978
rect 129942 226294 129998 226350
rect 130066 226294 130122 226350
rect 129942 226170 129998 226226
rect 130066 226170 130122 226226
rect 129942 226046 129998 226102
rect 130066 226046 130122 226102
rect 129942 225922 129998 225978
rect 130066 225922 130122 225978
rect 22422 220294 22478 220350
rect 22546 220294 22602 220350
rect 22422 220170 22478 220226
rect 22546 220170 22602 220226
rect 22422 220046 22478 220102
rect 22546 220046 22602 220102
rect 22422 219922 22478 219978
rect 22546 219922 22602 219978
rect 53142 220294 53198 220350
rect 53266 220294 53322 220350
rect 53142 220170 53198 220226
rect 53266 220170 53322 220226
rect 53142 220046 53198 220102
rect 53266 220046 53322 220102
rect 53142 219922 53198 219978
rect 53266 219922 53322 219978
rect 83862 220294 83918 220350
rect 83986 220294 84042 220350
rect 83862 220170 83918 220226
rect 83986 220170 84042 220226
rect 83862 220046 83918 220102
rect 83986 220046 84042 220102
rect 83862 219922 83918 219978
rect 83986 219922 84042 219978
rect 114582 220294 114638 220350
rect 114706 220294 114762 220350
rect 114582 220170 114638 220226
rect 114706 220170 114762 220226
rect 114582 220046 114638 220102
rect 114706 220046 114762 220102
rect 114582 219922 114638 219978
rect 114706 219922 114762 219978
rect 145302 220294 145358 220350
rect 145426 220294 145482 220350
rect 145302 220170 145358 220226
rect 145426 220170 145482 220226
rect 145302 220046 145358 220102
rect 145426 220046 145482 220102
rect 145302 219922 145358 219978
rect 145426 219922 145482 219978
rect 37782 208294 37838 208350
rect 37906 208294 37962 208350
rect 37782 208170 37838 208226
rect 37906 208170 37962 208226
rect 37782 208046 37838 208102
rect 37906 208046 37962 208102
rect 37782 207922 37838 207978
rect 37906 207922 37962 207978
rect 68502 208294 68558 208350
rect 68626 208294 68682 208350
rect 68502 208170 68558 208226
rect 68626 208170 68682 208226
rect 68502 208046 68558 208102
rect 68626 208046 68682 208102
rect 68502 207922 68558 207978
rect 68626 207922 68682 207978
rect 99222 208294 99278 208350
rect 99346 208294 99402 208350
rect 99222 208170 99278 208226
rect 99346 208170 99402 208226
rect 99222 208046 99278 208102
rect 99346 208046 99402 208102
rect 99222 207922 99278 207978
rect 99346 207922 99402 207978
rect 129942 208294 129998 208350
rect 130066 208294 130122 208350
rect 129942 208170 129998 208226
rect 130066 208170 130122 208226
rect 129942 208046 129998 208102
rect 130066 208046 130122 208102
rect 129942 207922 129998 207978
rect 130066 207922 130122 207978
rect 22422 202294 22478 202350
rect 22546 202294 22602 202350
rect 22422 202170 22478 202226
rect 22546 202170 22602 202226
rect 22422 202046 22478 202102
rect 22546 202046 22602 202102
rect 22422 201922 22478 201978
rect 22546 201922 22602 201978
rect 53142 202294 53198 202350
rect 53266 202294 53322 202350
rect 53142 202170 53198 202226
rect 53266 202170 53322 202226
rect 53142 202046 53198 202102
rect 53266 202046 53322 202102
rect 53142 201922 53198 201978
rect 53266 201922 53322 201978
rect 83862 202294 83918 202350
rect 83986 202294 84042 202350
rect 83862 202170 83918 202226
rect 83986 202170 84042 202226
rect 83862 202046 83918 202102
rect 83986 202046 84042 202102
rect 83862 201922 83918 201978
rect 83986 201922 84042 201978
rect 114582 202294 114638 202350
rect 114706 202294 114762 202350
rect 114582 202170 114638 202226
rect 114706 202170 114762 202226
rect 114582 202046 114638 202102
rect 114706 202046 114762 202102
rect 114582 201922 114638 201978
rect 114706 201922 114762 201978
rect 145302 202294 145358 202350
rect 145426 202294 145482 202350
rect 145302 202170 145358 202226
rect 145426 202170 145482 202226
rect 145302 202046 145358 202102
rect 145426 202046 145482 202102
rect 145302 201922 145358 201978
rect 145426 201922 145482 201978
rect 37782 190294 37838 190350
rect 37906 190294 37962 190350
rect 37782 190170 37838 190226
rect 37906 190170 37962 190226
rect 37782 190046 37838 190102
rect 37906 190046 37962 190102
rect 37782 189922 37838 189978
rect 37906 189922 37962 189978
rect 68502 190294 68558 190350
rect 68626 190294 68682 190350
rect 68502 190170 68558 190226
rect 68626 190170 68682 190226
rect 68502 190046 68558 190102
rect 68626 190046 68682 190102
rect 68502 189922 68558 189978
rect 68626 189922 68682 189978
rect 99222 190294 99278 190350
rect 99346 190294 99402 190350
rect 99222 190170 99278 190226
rect 99346 190170 99402 190226
rect 99222 190046 99278 190102
rect 99346 190046 99402 190102
rect 99222 189922 99278 189978
rect 99346 189922 99402 189978
rect 129942 190294 129998 190350
rect 130066 190294 130122 190350
rect 129942 190170 129998 190226
rect 130066 190170 130122 190226
rect 129942 190046 129998 190102
rect 130066 190046 130122 190102
rect 129942 189922 129998 189978
rect 130066 189922 130122 189978
rect 22422 184294 22478 184350
rect 22546 184294 22602 184350
rect 22422 184170 22478 184226
rect 22546 184170 22602 184226
rect 22422 184046 22478 184102
rect 22546 184046 22602 184102
rect 22422 183922 22478 183978
rect 22546 183922 22602 183978
rect 53142 184294 53198 184350
rect 53266 184294 53322 184350
rect 53142 184170 53198 184226
rect 53266 184170 53322 184226
rect 53142 184046 53198 184102
rect 53266 184046 53322 184102
rect 53142 183922 53198 183978
rect 53266 183922 53322 183978
rect 83862 184294 83918 184350
rect 83986 184294 84042 184350
rect 83862 184170 83918 184226
rect 83986 184170 84042 184226
rect 83862 184046 83918 184102
rect 83986 184046 84042 184102
rect 83862 183922 83918 183978
rect 83986 183922 84042 183978
rect 114582 184294 114638 184350
rect 114706 184294 114762 184350
rect 114582 184170 114638 184226
rect 114706 184170 114762 184226
rect 114582 184046 114638 184102
rect 114706 184046 114762 184102
rect 114582 183922 114638 183978
rect 114706 183922 114762 183978
rect 145302 184294 145358 184350
rect 145426 184294 145482 184350
rect 145302 184170 145358 184226
rect 145426 184170 145482 184226
rect 145302 184046 145358 184102
rect 145426 184046 145482 184102
rect 145302 183922 145358 183978
rect 145426 183922 145482 183978
rect 37782 172294 37838 172350
rect 37906 172294 37962 172350
rect 37782 172170 37838 172226
rect 37906 172170 37962 172226
rect 37782 172046 37838 172102
rect 37906 172046 37962 172102
rect 37782 171922 37838 171978
rect 37906 171922 37962 171978
rect 68502 172294 68558 172350
rect 68626 172294 68682 172350
rect 68502 172170 68558 172226
rect 68626 172170 68682 172226
rect 68502 172046 68558 172102
rect 68626 172046 68682 172102
rect 68502 171922 68558 171978
rect 68626 171922 68682 171978
rect 99222 172294 99278 172350
rect 99346 172294 99402 172350
rect 99222 172170 99278 172226
rect 99346 172170 99402 172226
rect 99222 172046 99278 172102
rect 99346 172046 99402 172102
rect 99222 171922 99278 171978
rect 99346 171922 99402 171978
rect 129942 172294 129998 172350
rect 130066 172294 130122 172350
rect 129942 172170 129998 172226
rect 130066 172170 130122 172226
rect 129942 172046 129998 172102
rect 130066 172046 130122 172102
rect 129942 171922 129998 171978
rect 130066 171922 130122 171978
rect 22422 166294 22478 166350
rect 22546 166294 22602 166350
rect 22422 166170 22478 166226
rect 22546 166170 22602 166226
rect 22422 166046 22478 166102
rect 22546 166046 22602 166102
rect 22422 165922 22478 165978
rect 22546 165922 22602 165978
rect 53142 166294 53198 166350
rect 53266 166294 53322 166350
rect 53142 166170 53198 166226
rect 53266 166170 53322 166226
rect 53142 166046 53198 166102
rect 53266 166046 53322 166102
rect 53142 165922 53198 165978
rect 53266 165922 53322 165978
rect 83862 166294 83918 166350
rect 83986 166294 84042 166350
rect 83862 166170 83918 166226
rect 83986 166170 84042 166226
rect 83862 166046 83918 166102
rect 83986 166046 84042 166102
rect 83862 165922 83918 165978
rect 83986 165922 84042 165978
rect 114582 166294 114638 166350
rect 114706 166294 114762 166350
rect 114582 166170 114638 166226
rect 114706 166170 114762 166226
rect 114582 166046 114638 166102
rect 114706 166046 114762 166102
rect 114582 165922 114638 165978
rect 114706 165922 114762 165978
rect 145302 166294 145358 166350
rect 145426 166294 145482 166350
rect 145302 166170 145358 166226
rect 145426 166170 145482 166226
rect 145302 166046 145358 166102
rect 145426 166046 145482 166102
rect 145302 165922 145358 165978
rect 145426 165922 145482 165978
rect 37782 154294 37838 154350
rect 37906 154294 37962 154350
rect 37782 154170 37838 154226
rect 37906 154170 37962 154226
rect 37782 154046 37838 154102
rect 37906 154046 37962 154102
rect 37782 153922 37838 153978
rect 37906 153922 37962 153978
rect 68502 154294 68558 154350
rect 68626 154294 68682 154350
rect 68502 154170 68558 154226
rect 68626 154170 68682 154226
rect 68502 154046 68558 154102
rect 68626 154046 68682 154102
rect 68502 153922 68558 153978
rect 68626 153922 68682 153978
rect 99222 154294 99278 154350
rect 99346 154294 99402 154350
rect 99222 154170 99278 154226
rect 99346 154170 99402 154226
rect 99222 154046 99278 154102
rect 99346 154046 99402 154102
rect 99222 153922 99278 153978
rect 99346 153922 99402 153978
rect 129942 154294 129998 154350
rect 130066 154294 130122 154350
rect 129942 154170 129998 154226
rect 130066 154170 130122 154226
rect 129942 154046 129998 154102
rect 130066 154046 130122 154102
rect 129942 153922 129998 153978
rect 130066 153922 130122 153978
rect 22422 148294 22478 148350
rect 22546 148294 22602 148350
rect 22422 148170 22478 148226
rect 22546 148170 22602 148226
rect 22422 148046 22478 148102
rect 22546 148046 22602 148102
rect 22422 147922 22478 147978
rect 22546 147922 22602 147978
rect 53142 148294 53198 148350
rect 53266 148294 53322 148350
rect 53142 148170 53198 148226
rect 53266 148170 53322 148226
rect 53142 148046 53198 148102
rect 53266 148046 53322 148102
rect 53142 147922 53198 147978
rect 53266 147922 53322 147978
rect 83862 148294 83918 148350
rect 83986 148294 84042 148350
rect 83862 148170 83918 148226
rect 83986 148170 84042 148226
rect 83862 148046 83918 148102
rect 83986 148046 84042 148102
rect 83862 147922 83918 147978
rect 83986 147922 84042 147978
rect 114582 148294 114638 148350
rect 114706 148294 114762 148350
rect 114582 148170 114638 148226
rect 114706 148170 114762 148226
rect 114582 148046 114638 148102
rect 114706 148046 114762 148102
rect 114582 147922 114638 147978
rect 114706 147922 114762 147978
rect 145302 148294 145358 148350
rect 145426 148294 145482 148350
rect 145302 148170 145358 148226
rect 145426 148170 145482 148226
rect 145302 148046 145358 148102
rect 145426 148046 145482 148102
rect 145302 147922 145358 147978
rect 145426 147922 145482 147978
rect 37782 136294 37838 136350
rect 37906 136294 37962 136350
rect 37782 136170 37838 136226
rect 37906 136170 37962 136226
rect 37782 136046 37838 136102
rect 37906 136046 37962 136102
rect 37782 135922 37838 135978
rect 37906 135922 37962 135978
rect 68502 136294 68558 136350
rect 68626 136294 68682 136350
rect 68502 136170 68558 136226
rect 68626 136170 68682 136226
rect 68502 136046 68558 136102
rect 68626 136046 68682 136102
rect 68502 135922 68558 135978
rect 68626 135922 68682 135978
rect 99222 136294 99278 136350
rect 99346 136294 99402 136350
rect 99222 136170 99278 136226
rect 99346 136170 99402 136226
rect 99222 136046 99278 136102
rect 99346 136046 99402 136102
rect 99222 135922 99278 135978
rect 99346 135922 99402 135978
rect 129942 136294 129998 136350
rect 130066 136294 130122 136350
rect 129942 136170 129998 136226
rect 130066 136170 130122 136226
rect 129942 136046 129998 136102
rect 130066 136046 130122 136102
rect 129942 135922 129998 135978
rect 130066 135922 130122 135978
rect 22422 130294 22478 130350
rect 22546 130294 22602 130350
rect 22422 130170 22478 130226
rect 22546 130170 22602 130226
rect 22422 130046 22478 130102
rect 22546 130046 22602 130102
rect 22422 129922 22478 129978
rect 22546 129922 22602 129978
rect 53142 130294 53198 130350
rect 53266 130294 53322 130350
rect 53142 130170 53198 130226
rect 53266 130170 53322 130226
rect 53142 130046 53198 130102
rect 53266 130046 53322 130102
rect 53142 129922 53198 129978
rect 53266 129922 53322 129978
rect 83862 130294 83918 130350
rect 83986 130294 84042 130350
rect 83862 130170 83918 130226
rect 83986 130170 84042 130226
rect 83862 130046 83918 130102
rect 83986 130046 84042 130102
rect 83862 129922 83918 129978
rect 83986 129922 84042 129978
rect 114582 130294 114638 130350
rect 114706 130294 114762 130350
rect 114582 130170 114638 130226
rect 114706 130170 114762 130226
rect 114582 130046 114638 130102
rect 114706 130046 114762 130102
rect 114582 129922 114638 129978
rect 114706 129922 114762 129978
rect 145302 130294 145358 130350
rect 145426 130294 145482 130350
rect 145302 130170 145358 130226
rect 145426 130170 145482 130226
rect 145302 130046 145358 130102
rect 145426 130046 145482 130102
rect 145302 129922 145358 129978
rect 145426 129922 145482 129978
rect 37782 118294 37838 118350
rect 37906 118294 37962 118350
rect 37782 118170 37838 118226
rect 37906 118170 37962 118226
rect 37782 118046 37838 118102
rect 37906 118046 37962 118102
rect 37782 117922 37838 117978
rect 37906 117922 37962 117978
rect 68502 118294 68558 118350
rect 68626 118294 68682 118350
rect 68502 118170 68558 118226
rect 68626 118170 68682 118226
rect 68502 118046 68558 118102
rect 68626 118046 68682 118102
rect 68502 117922 68558 117978
rect 68626 117922 68682 117978
rect 99222 118294 99278 118350
rect 99346 118294 99402 118350
rect 99222 118170 99278 118226
rect 99346 118170 99402 118226
rect 99222 118046 99278 118102
rect 99346 118046 99402 118102
rect 99222 117922 99278 117978
rect 99346 117922 99402 117978
rect 129942 118294 129998 118350
rect 130066 118294 130122 118350
rect 129942 118170 129998 118226
rect 130066 118170 130122 118226
rect 129942 118046 129998 118102
rect 130066 118046 130122 118102
rect 129942 117922 129998 117978
rect 130066 117922 130122 117978
rect 22422 112294 22478 112350
rect 22546 112294 22602 112350
rect 22422 112170 22478 112226
rect 22546 112170 22602 112226
rect 22422 112046 22478 112102
rect 22546 112046 22602 112102
rect 22422 111922 22478 111978
rect 22546 111922 22602 111978
rect 53142 112294 53198 112350
rect 53266 112294 53322 112350
rect 53142 112170 53198 112226
rect 53266 112170 53322 112226
rect 53142 112046 53198 112102
rect 53266 112046 53322 112102
rect 53142 111922 53198 111978
rect 53266 111922 53322 111978
rect 83862 112294 83918 112350
rect 83986 112294 84042 112350
rect 83862 112170 83918 112226
rect 83986 112170 84042 112226
rect 83862 112046 83918 112102
rect 83986 112046 84042 112102
rect 83862 111922 83918 111978
rect 83986 111922 84042 111978
rect 114582 112294 114638 112350
rect 114706 112294 114762 112350
rect 114582 112170 114638 112226
rect 114706 112170 114762 112226
rect 114582 112046 114638 112102
rect 114706 112046 114762 112102
rect 114582 111922 114638 111978
rect 114706 111922 114762 111978
rect 145302 112294 145358 112350
rect 145426 112294 145482 112350
rect 145302 112170 145358 112226
rect 145426 112170 145482 112226
rect 145302 112046 145358 112102
rect 145426 112046 145482 112102
rect 145302 111922 145358 111978
rect 145426 111922 145482 111978
rect 37782 100294 37838 100350
rect 37906 100294 37962 100350
rect 37782 100170 37838 100226
rect 37906 100170 37962 100226
rect 37782 100046 37838 100102
rect 37906 100046 37962 100102
rect 37782 99922 37838 99978
rect 37906 99922 37962 99978
rect 68502 100294 68558 100350
rect 68626 100294 68682 100350
rect 68502 100170 68558 100226
rect 68626 100170 68682 100226
rect 68502 100046 68558 100102
rect 68626 100046 68682 100102
rect 68502 99922 68558 99978
rect 68626 99922 68682 99978
rect 99222 100294 99278 100350
rect 99346 100294 99402 100350
rect 99222 100170 99278 100226
rect 99346 100170 99402 100226
rect 99222 100046 99278 100102
rect 99346 100046 99402 100102
rect 99222 99922 99278 99978
rect 99346 99922 99402 99978
rect 129942 100294 129998 100350
rect 130066 100294 130122 100350
rect 129942 100170 129998 100226
rect 130066 100170 130122 100226
rect 129942 100046 129998 100102
rect 130066 100046 130122 100102
rect 129942 99922 129998 99978
rect 130066 99922 130122 99978
rect 22422 94294 22478 94350
rect 22546 94294 22602 94350
rect 22422 94170 22478 94226
rect 22546 94170 22602 94226
rect 22422 94046 22478 94102
rect 22546 94046 22602 94102
rect 22422 93922 22478 93978
rect 22546 93922 22602 93978
rect 53142 94294 53198 94350
rect 53266 94294 53322 94350
rect 53142 94170 53198 94226
rect 53266 94170 53322 94226
rect 53142 94046 53198 94102
rect 53266 94046 53322 94102
rect 53142 93922 53198 93978
rect 53266 93922 53322 93978
rect 83862 94294 83918 94350
rect 83986 94294 84042 94350
rect 83862 94170 83918 94226
rect 83986 94170 84042 94226
rect 83862 94046 83918 94102
rect 83986 94046 84042 94102
rect 83862 93922 83918 93978
rect 83986 93922 84042 93978
rect 114582 94294 114638 94350
rect 114706 94294 114762 94350
rect 114582 94170 114638 94226
rect 114706 94170 114762 94226
rect 114582 94046 114638 94102
rect 114706 94046 114762 94102
rect 114582 93922 114638 93978
rect 114706 93922 114762 93978
rect 145302 94294 145358 94350
rect 145426 94294 145482 94350
rect 145302 94170 145358 94226
rect 145426 94170 145482 94226
rect 145302 94046 145358 94102
rect 145426 94046 145482 94102
rect 145302 93922 145358 93978
rect 145426 93922 145482 93978
rect 37782 82294 37838 82350
rect 37906 82294 37962 82350
rect 37782 82170 37838 82226
rect 37906 82170 37962 82226
rect 37782 82046 37838 82102
rect 37906 82046 37962 82102
rect 37782 81922 37838 81978
rect 37906 81922 37962 81978
rect 68502 82294 68558 82350
rect 68626 82294 68682 82350
rect 68502 82170 68558 82226
rect 68626 82170 68682 82226
rect 68502 82046 68558 82102
rect 68626 82046 68682 82102
rect 68502 81922 68558 81978
rect 68626 81922 68682 81978
rect 99222 82294 99278 82350
rect 99346 82294 99402 82350
rect 99222 82170 99278 82226
rect 99346 82170 99402 82226
rect 99222 82046 99278 82102
rect 99346 82046 99402 82102
rect 99222 81922 99278 81978
rect 99346 81922 99402 81978
rect 129942 82294 129998 82350
rect 130066 82294 130122 82350
rect 129942 82170 129998 82226
rect 130066 82170 130122 82226
rect 129942 82046 129998 82102
rect 130066 82046 130122 82102
rect 129942 81922 129998 81978
rect 130066 81922 130122 81978
rect 22422 76294 22478 76350
rect 22546 76294 22602 76350
rect 22422 76170 22478 76226
rect 22546 76170 22602 76226
rect 22422 76046 22478 76102
rect 22546 76046 22602 76102
rect 22422 75922 22478 75978
rect 22546 75922 22602 75978
rect 53142 76294 53198 76350
rect 53266 76294 53322 76350
rect 53142 76170 53198 76226
rect 53266 76170 53322 76226
rect 53142 76046 53198 76102
rect 53266 76046 53322 76102
rect 53142 75922 53198 75978
rect 53266 75922 53322 75978
rect 83862 76294 83918 76350
rect 83986 76294 84042 76350
rect 83862 76170 83918 76226
rect 83986 76170 84042 76226
rect 83862 76046 83918 76102
rect 83986 76046 84042 76102
rect 83862 75922 83918 75978
rect 83986 75922 84042 75978
rect 114582 76294 114638 76350
rect 114706 76294 114762 76350
rect 114582 76170 114638 76226
rect 114706 76170 114762 76226
rect 114582 76046 114638 76102
rect 114706 76046 114762 76102
rect 114582 75922 114638 75978
rect 114706 75922 114762 75978
rect 145302 76294 145358 76350
rect 145426 76294 145482 76350
rect 145302 76170 145358 76226
rect 145426 76170 145482 76226
rect 145302 76046 145358 76102
rect 145426 76046 145482 76102
rect 145302 75922 145358 75978
rect 145426 75922 145482 75978
rect 37782 64294 37838 64350
rect 37906 64294 37962 64350
rect 37782 64170 37838 64226
rect 37906 64170 37962 64226
rect 37782 64046 37838 64102
rect 37906 64046 37962 64102
rect 37782 63922 37838 63978
rect 37906 63922 37962 63978
rect 68502 64294 68558 64350
rect 68626 64294 68682 64350
rect 68502 64170 68558 64226
rect 68626 64170 68682 64226
rect 68502 64046 68558 64102
rect 68626 64046 68682 64102
rect 68502 63922 68558 63978
rect 68626 63922 68682 63978
rect 99222 64294 99278 64350
rect 99346 64294 99402 64350
rect 99222 64170 99278 64226
rect 99346 64170 99402 64226
rect 99222 64046 99278 64102
rect 99346 64046 99402 64102
rect 99222 63922 99278 63978
rect 99346 63922 99402 63978
rect 129942 64294 129998 64350
rect 130066 64294 130122 64350
rect 129942 64170 129998 64226
rect 130066 64170 130122 64226
rect 129942 64046 129998 64102
rect 130066 64046 130122 64102
rect 129942 63922 129998 63978
rect 130066 63922 130122 63978
rect 22422 58294 22478 58350
rect 22546 58294 22602 58350
rect 22422 58170 22478 58226
rect 22546 58170 22602 58226
rect 22422 58046 22478 58102
rect 22546 58046 22602 58102
rect 22422 57922 22478 57978
rect 22546 57922 22602 57978
rect 53142 58294 53198 58350
rect 53266 58294 53322 58350
rect 53142 58170 53198 58226
rect 53266 58170 53322 58226
rect 53142 58046 53198 58102
rect 53266 58046 53322 58102
rect 53142 57922 53198 57978
rect 53266 57922 53322 57978
rect 83862 58294 83918 58350
rect 83986 58294 84042 58350
rect 83862 58170 83918 58226
rect 83986 58170 84042 58226
rect 83862 58046 83918 58102
rect 83986 58046 84042 58102
rect 83862 57922 83918 57978
rect 83986 57922 84042 57978
rect 114582 58294 114638 58350
rect 114706 58294 114762 58350
rect 114582 58170 114638 58226
rect 114706 58170 114762 58226
rect 114582 58046 114638 58102
rect 114706 58046 114762 58102
rect 114582 57922 114638 57978
rect 114706 57922 114762 57978
rect 145302 58294 145358 58350
rect 145426 58294 145482 58350
rect 145302 58170 145358 58226
rect 145426 58170 145482 58226
rect 145302 58046 145358 58102
rect 145426 58046 145482 58102
rect 145302 57922 145358 57978
rect 145426 57922 145482 57978
rect 37782 46294 37838 46350
rect 37906 46294 37962 46350
rect 37782 46170 37838 46226
rect 37906 46170 37962 46226
rect 37782 46046 37838 46102
rect 37906 46046 37962 46102
rect 37782 45922 37838 45978
rect 37906 45922 37962 45978
rect 68502 46294 68558 46350
rect 68626 46294 68682 46350
rect 68502 46170 68558 46226
rect 68626 46170 68682 46226
rect 68502 46046 68558 46102
rect 68626 46046 68682 46102
rect 68502 45922 68558 45978
rect 68626 45922 68682 45978
rect 99222 46294 99278 46350
rect 99346 46294 99402 46350
rect 99222 46170 99278 46226
rect 99346 46170 99402 46226
rect 99222 46046 99278 46102
rect 99346 46046 99402 46102
rect 99222 45922 99278 45978
rect 99346 45922 99402 45978
rect 129942 46294 129998 46350
rect 130066 46294 130122 46350
rect 129942 46170 129998 46226
rect 130066 46170 130122 46226
rect 129942 46046 129998 46102
rect 130066 46046 130122 46102
rect 129942 45922 129998 45978
rect 130066 45922 130122 45978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 22422 40294 22478 40350
rect 22546 40294 22602 40350
rect 22422 40170 22478 40226
rect 22546 40170 22602 40226
rect 22422 40046 22478 40102
rect 22546 40046 22602 40102
rect 22422 39922 22478 39978
rect 22546 39922 22602 39978
rect 53142 40294 53198 40350
rect 53266 40294 53322 40350
rect 53142 40170 53198 40226
rect 53266 40170 53322 40226
rect 53142 40046 53198 40102
rect 53266 40046 53322 40102
rect 53142 39922 53198 39978
rect 53266 39922 53322 39978
rect 83862 40294 83918 40350
rect 83986 40294 84042 40350
rect 83862 40170 83918 40226
rect 83986 40170 84042 40226
rect 83862 40046 83918 40102
rect 83986 40046 84042 40102
rect 83862 39922 83918 39978
rect 83986 39922 84042 39978
rect 114582 40294 114638 40350
rect 114706 40294 114762 40350
rect 114582 40170 114638 40226
rect 114706 40170 114762 40226
rect 114582 40046 114638 40102
rect 114706 40046 114762 40102
rect 114582 39922 114638 39978
rect 114706 39922 114762 39978
rect 145302 40294 145358 40350
rect 145426 40294 145482 40350
rect 145302 40170 145358 40226
rect 145426 40170 145482 40226
rect 145302 40046 145358 40102
rect 145426 40046 145482 40102
rect 145302 39922 145358 39978
rect 145426 39922 145482 39978
rect 37782 28294 37838 28350
rect 37906 28294 37962 28350
rect 37782 28170 37838 28226
rect 37906 28170 37962 28226
rect 37782 28046 37838 28102
rect 37906 28046 37962 28102
rect 37782 27922 37838 27978
rect 37906 27922 37962 27978
rect 68502 28294 68558 28350
rect 68626 28294 68682 28350
rect 68502 28170 68558 28226
rect 68626 28170 68682 28226
rect 68502 28046 68558 28102
rect 68626 28046 68682 28102
rect 68502 27922 68558 27978
rect 68626 27922 68682 27978
rect 99222 28294 99278 28350
rect 99346 28294 99402 28350
rect 99222 28170 99278 28226
rect 99346 28170 99402 28226
rect 99222 28046 99278 28102
rect 99346 28046 99402 28102
rect 99222 27922 99278 27978
rect 99346 27922 99402 27978
rect 129942 28294 129998 28350
rect 130066 28294 130122 28350
rect 129942 28170 129998 28226
rect 130066 28170 130122 28226
rect 129942 28046 129998 28102
rect 130066 28046 130122 28102
rect 129942 27922 129998 27978
rect 130066 27922 130122 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 23436 13562 23492 13618
rect 17276 9242 17332 9298
rect 11564 5822 11620 5878
rect 26796 6002 26852 6058
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 13356 3302 13412 3358
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 44492 11762 44548 11818
rect 55356 7622 55412 7678
rect 41804 7442 41860 7498
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 159114 346294 159170 346350
rect 159238 346294 159294 346350
rect 159362 346294 159418 346350
rect 159486 346294 159542 346350
rect 159114 346170 159170 346226
rect 159238 346170 159294 346226
rect 159362 346170 159418 346226
rect 159486 346170 159542 346226
rect 159114 346046 159170 346102
rect 159238 346046 159294 346102
rect 159362 346046 159418 346102
rect 159486 346046 159542 346102
rect 159114 345922 159170 345978
rect 159238 345922 159294 345978
rect 159362 345922 159418 345978
rect 159486 345922 159542 345978
rect 159114 328294 159170 328350
rect 159238 328294 159294 328350
rect 159362 328294 159418 328350
rect 159486 328294 159542 328350
rect 159114 328170 159170 328226
rect 159238 328170 159294 328226
rect 159362 328170 159418 328226
rect 159486 328170 159542 328226
rect 159114 328046 159170 328102
rect 159238 328046 159294 328102
rect 159362 328046 159418 328102
rect 159486 328046 159542 328102
rect 159114 327922 159170 327978
rect 159238 327922 159294 327978
rect 159362 327922 159418 327978
rect 159486 327922 159542 327978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 159114 274294 159170 274350
rect 159238 274294 159294 274350
rect 159362 274294 159418 274350
rect 159486 274294 159542 274350
rect 159114 274170 159170 274226
rect 159238 274170 159294 274226
rect 159362 274170 159418 274226
rect 159486 274170 159542 274226
rect 159114 274046 159170 274102
rect 159238 274046 159294 274102
rect 159362 274046 159418 274102
rect 159486 274046 159542 274102
rect 159114 273922 159170 273978
rect 159238 273922 159294 273978
rect 159362 273922 159418 273978
rect 159486 273922 159542 273978
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 159114 202294 159170 202350
rect 159238 202294 159294 202350
rect 159362 202294 159418 202350
rect 159486 202294 159542 202350
rect 159114 202170 159170 202226
rect 159238 202170 159294 202226
rect 159362 202170 159418 202226
rect 159486 202170 159542 202226
rect 159114 202046 159170 202102
rect 159238 202046 159294 202102
rect 159362 202046 159418 202102
rect 159486 202046 159542 202102
rect 159114 201922 159170 201978
rect 159238 201922 159294 201978
rect 159362 201922 159418 201978
rect 159486 201922 159542 201978
rect 159114 184294 159170 184350
rect 159238 184294 159294 184350
rect 159362 184294 159418 184350
rect 159486 184294 159542 184350
rect 159114 184170 159170 184226
rect 159238 184170 159294 184226
rect 159362 184170 159418 184226
rect 159486 184170 159542 184226
rect 159114 184046 159170 184102
rect 159238 184046 159294 184102
rect 159362 184046 159418 184102
rect 159486 184046 159542 184102
rect 159114 183922 159170 183978
rect 159238 183922 159294 183978
rect 159362 183922 159418 183978
rect 159486 183922 159542 183978
rect 159114 166294 159170 166350
rect 159238 166294 159294 166350
rect 159362 166294 159418 166350
rect 159486 166294 159542 166350
rect 159114 166170 159170 166226
rect 159238 166170 159294 166226
rect 159362 166170 159418 166226
rect 159486 166170 159542 166226
rect 159114 166046 159170 166102
rect 159238 166046 159294 166102
rect 159362 166046 159418 166102
rect 159486 166046 159542 166102
rect 159114 165922 159170 165978
rect 159238 165922 159294 165978
rect 159362 165922 159418 165978
rect 159486 165922 159542 165978
rect 159114 148294 159170 148350
rect 159238 148294 159294 148350
rect 159362 148294 159418 148350
rect 159486 148294 159542 148350
rect 159114 148170 159170 148226
rect 159238 148170 159294 148226
rect 159362 148170 159418 148226
rect 159486 148170 159542 148226
rect 159114 148046 159170 148102
rect 159238 148046 159294 148102
rect 159362 148046 159418 148102
rect 159486 148046 159542 148102
rect 159114 147922 159170 147978
rect 159238 147922 159294 147978
rect 159362 147922 159418 147978
rect 159486 147922 159542 147978
rect 159114 130294 159170 130350
rect 159238 130294 159294 130350
rect 159362 130294 159418 130350
rect 159486 130294 159542 130350
rect 159114 130170 159170 130226
rect 159238 130170 159294 130226
rect 159362 130170 159418 130226
rect 159486 130170 159542 130226
rect 159114 130046 159170 130102
rect 159238 130046 159294 130102
rect 159362 130046 159418 130102
rect 159486 130046 159542 130102
rect 159114 129922 159170 129978
rect 159238 129922 159294 129978
rect 159362 129922 159418 129978
rect 159486 129922 159542 129978
rect 159114 112294 159170 112350
rect 159238 112294 159294 112350
rect 159362 112294 159418 112350
rect 159486 112294 159542 112350
rect 159114 112170 159170 112226
rect 159238 112170 159294 112226
rect 159362 112170 159418 112226
rect 159486 112170 159542 112226
rect 159114 112046 159170 112102
rect 159238 112046 159294 112102
rect 159362 112046 159418 112102
rect 159486 112046 159542 112102
rect 159114 111922 159170 111978
rect 159238 111922 159294 111978
rect 159362 111922 159418 111978
rect 159486 111922 159542 111978
rect 159114 94294 159170 94350
rect 159238 94294 159294 94350
rect 159362 94294 159418 94350
rect 159486 94294 159542 94350
rect 159114 94170 159170 94226
rect 159238 94170 159294 94226
rect 159362 94170 159418 94226
rect 159486 94170 159542 94226
rect 159114 94046 159170 94102
rect 159238 94046 159294 94102
rect 159362 94046 159418 94102
rect 159486 94046 159542 94102
rect 159114 93922 159170 93978
rect 159238 93922 159294 93978
rect 159362 93922 159418 93978
rect 159486 93922 159542 93978
rect 159114 76294 159170 76350
rect 159238 76294 159294 76350
rect 159362 76294 159418 76350
rect 159486 76294 159542 76350
rect 159114 76170 159170 76226
rect 159238 76170 159294 76226
rect 159362 76170 159418 76226
rect 159486 76170 159542 76226
rect 159114 76046 159170 76102
rect 159238 76046 159294 76102
rect 159362 76046 159418 76102
rect 159486 76046 159542 76102
rect 159114 75922 159170 75978
rect 159238 75922 159294 75978
rect 159362 75922 159418 75978
rect 159486 75922 159542 75978
rect 159114 58294 159170 58350
rect 159238 58294 159294 58350
rect 159362 58294 159418 58350
rect 159486 58294 159542 58350
rect 159114 58170 159170 58226
rect 159238 58170 159294 58226
rect 159362 58170 159418 58226
rect 159486 58170 159542 58226
rect 159114 58046 159170 58102
rect 159238 58046 159294 58102
rect 159362 58046 159418 58102
rect 159486 58046 159542 58102
rect 159114 57922 159170 57978
rect 159238 57922 159294 57978
rect 159362 57922 159418 57978
rect 159486 57922 159542 57978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 162834 352294 162890 352350
rect 162958 352294 163014 352350
rect 163082 352294 163138 352350
rect 163206 352294 163262 352350
rect 162834 352170 162890 352226
rect 162958 352170 163014 352226
rect 163082 352170 163138 352226
rect 163206 352170 163262 352226
rect 162834 352046 162890 352102
rect 162958 352046 163014 352102
rect 163082 352046 163138 352102
rect 163206 352046 163262 352102
rect 162834 351922 162890 351978
rect 162958 351922 163014 351978
rect 163082 351922 163138 351978
rect 163206 351922 163262 351978
rect 162834 334294 162890 334350
rect 162958 334294 163014 334350
rect 163082 334294 163138 334350
rect 163206 334294 163262 334350
rect 162834 334170 162890 334226
rect 162958 334170 163014 334226
rect 163082 334170 163138 334226
rect 163206 334170 163262 334226
rect 162834 334046 162890 334102
rect 162958 334046 163014 334102
rect 163082 334046 163138 334102
rect 163206 334046 163262 334102
rect 162834 333922 162890 333978
rect 162958 333922 163014 333978
rect 163082 333922 163138 333978
rect 163206 333922 163262 333978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 162834 262294 162890 262350
rect 162958 262294 163014 262350
rect 163082 262294 163138 262350
rect 163206 262294 163262 262350
rect 162834 262170 162890 262226
rect 162958 262170 163014 262226
rect 163082 262170 163138 262226
rect 163206 262170 163262 262226
rect 162834 262046 162890 262102
rect 162958 262046 163014 262102
rect 163082 262046 163138 262102
rect 163206 262046 163262 262102
rect 162834 261922 162890 261978
rect 162958 261922 163014 261978
rect 163082 261922 163138 261978
rect 163206 261922 163262 261978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 162834 208294 162890 208350
rect 162958 208294 163014 208350
rect 163082 208294 163138 208350
rect 163206 208294 163262 208350
rect 162834 208170 162890 208226
rect 162958 208170 163014 208226
rect 163082 208170 163138 208226
rect 163206 208170 163262 208226
rect 162834 208046 162890 208102
rect 162958 208046 163014 208102
rect 163082 208046 163138 208102
rect 163206 208046 163262 208102
rect 162834 207922 162890 207978
rect 162958 207922 163014 207978
rect 163082 207922 163138 207978
rect 163206 207922 163262 207978
rect 162834 190294 162890 190350
rect 162958 190294 163014 190350
rect 163082 190294 163138 190350
rect 163206 190294 163262 190350
rect 162834 190170 162890 190226
rect 162958 190170 163014 190226
rect 163082 190170 163138 190226
rect 163206 190170 163262 190226
rect 162834 190046 162890 190102
rect 162958 190046 163014 190102
rect 163082 190046 163138 190102
rect 163206 190046 163262 190102
rect 162834 189922 162890 189978
rect 162958 189922 163014 189978
rect 163082 189922 163138 189978
rect 163206 189922 163262 189978
rect 162834 172294 162890 172350
rect 162958 172294 163014 172350
rect 163082 172294 163138 172350
rect 163206 172294 163262 172350
rect 162834 172170 162890 172226
rect 162958 172170 163014 172226
rect 163082 172170 163138 172226
rect 163206 172170 163262 172226
rect 162834 172046 162890 172102
rect 162958 172046 163014 172102
rect 163082 172046 163138 172102
rect 163206 172046 163262 172102
rect 162834 171922 162890 171978
rect 162958 171922 163014 171978
rect 163082 171922 163138 171978
rect 163206 171922 163262 171978
rect 162834 154294 162890 154350
rect 162958 154294 163014 154350
rect 163082 154294 163138 154350
rect 163206 154294 163262 154350
rect 162834 154170 162890 154226
rect 162958 154170 163014 154226
rect 163082 154170 163138 154226
rect 163206 154170 163262 154226
rect 162834 154046 162890 154102
rect 162958 154046 163014 154102
rect 163082 154046 163138 154102
rect 163206 154046 163262 154102
rect 162834 153922 162890 153978
rect 162958 153922 163014 153978
rect 163082 153922 163138 153978
rect 163206 153922 163262 153978
rect 162834 136294 162890 136350
rect 162958 136294 163014 136350
rect 163082 136294 163138 136350
rect 163206 136294 163262 136350
rect 162834 136170 162890 136226
rect 162958 136170 163014 136226
rect 163082 136170 163138 136226
rect 163206 136170 163262 136226
rect 162834 136046 162890 136102
rect 162958 136046 163014 136102
rect 163082 136046 163138 136102
rect 163206 136046 163262 136102
rect 162834 135922 162890 135978
rect 162958 135922 163014 135978
rect 163082 135922 163138 135978
rect 163206 135922 163262 135978
rect 162834 118294 162890 118350
rect 162958 118294 163014 118350
rect 163082 118294 163138 118350
rect 163206 118294 163262 118350
rect 162834 118170 162890 118226
rect 162958 118170 163014 118226
rect 163082 118170 163138 118226
rect 163206 118170 163262 118226
rect 162834 118046 162890 118102
rect 162958 118046 163014 118102
rect 163082 118046 163138 118102
rect 163206 118046 163262 118102
rect 162834 117922 162890 117978
rect 162958 117922 163014 117978
rect 163082 117922 163138 117978
rect 163206 117922 163262 117978
rect 162834 100294 162890 100350
rect 162958 100294 163014 100350
rect 163082 100294 163138 100350
rect 163206 100294 163262 100350
rect 162834 100170 162890 100226
rect 162958 100170 163014 100226
rect 163082 100170 163138 100226
rect 163206 100170 163262 100226
rect 162834 100046 162890 100102
rect 162958 100046 163014 100102
rect 163082 100046 163138 100102
rect 163206 100046 163262 100102
rect 162834 99922 162890 99978
rect 162958 99922 163014 99978
rect 163082 99922 163138 99978
rect 163206 99922 163262 99978
rect 162834 82294 162890 82350
rect 162958 82294 163014 82350
rect 163082 82294 163138 82350
rect 163206 82294 163262 82350
rect 162834 82170 162890 82226
rect 162958 82170 163014 82226
rect 163082 82170 163138 82226
rect 163206 82170 163262 82226
rect 162834 82046 162890 82102
rect 162958 82046 163014 82102
rect 163082 82046 163138 82102
rect 163206 82046 163262 82102
rect 162834 81922 162890 81978
rect 162958 81922 163014 81978
rect 163082 81922 163138 81978
rect 163206 81922 163262 81978
rect 162834 64294 162890 64350
rect 162958 64294 163014 64350
rect 163082 64294 163138 64350
rect 163206 64294 163262 64350
rect 162834 64170 162890 64226
rect 162958 64170 163014 64226
rect 163082 64170 163138 64226
rect 163206 64170 163262 64226
rect 162834 64046 162890 64102
rect 162958 64046 163014 64102
rect 163082 64046 163138 64102
rect 163206 64046 163262 64102
rect 162834 63922 162890 63978
rect 162958 63922 163014 63978
rect 163082 63922 163138 63978
rect 163206 63922 163262 63978
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 152012 16622 152068 16678
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 134428 11942 134484 11998
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 193878 370294 193934 370350
rect 194002 370294 194058 370350
rect 193878 370170 193934 370226
rect 194002 370170 194058 370226
rect 193878 370046 193934 370102
rect 194002 370046 194058 370102
rect 193878 369922 193934 369978
rect 194002 369922 194058 369978
rect 224598 370294 224654 370350
rect 224722 370294 224778 370350
rect 224598 370170 224654 370226
rect 224722 370170 224778 370226
rect 224598 370046 224654 370102
rect 224722 370046 224778 370102
rect 224598 369922 224654 369978
rect 224722 369922 224778 369978
rect 255318 370294 255374 370350
rect 255442 370294 255498 370350
rect 255318 370170 255374 370226
rect 255442 370170 255498 370226
rect 255318 370046 255374 370102
rect 255442 370046 255498 370102
rect 255318 369922 255374 369978
rect 255442 369922 255498 369978
rect 286038 370294 286094 370350
rect 286162 370294 286218 370350
rect 286038 370170 286094 370226
rect 286162 370170 286218 370226
rect 286038 370046 286094 370102
rect 286162 370046 286218 370102
rect 286038 369922 286094 369978
rect 286162 369922 286218 369978
rect 316758 370294 316814 370350
rect 316882 370294 316938 370350
rect 316758 370170 316814 370226
rect 316882 370170 316938 370226
rect 316758 370046 316814 370102
rect 316882 370046 316938 370102
rect 316758 369922 316814 369978
rect 316882 369922 316938 369978
rect 347478 370294 347534 370350
rect 347602 370294 347658 370350
rect 347478 370170 347534 370226
rect 347602 370170 347658 370226
rect 347478 370046 347534 370102
rect 347602 370046 347658 370102
rect 347478 369922 347534 369978
rect 347602 369922 347658 369978
rect 378198 370294 378254 370350
rect 378322 370294 378378 370350
rect 378198 370170 378254 370226
rect 378322 370170 378378 370226
rect 378198 370046 378254 370102
rect 378322 370046 378378 370102
rect 378198 369922 378254 369978
rect 378322 369922 378378 369978
rect 408918 370294 408974 370350
rect 409042 370294 409098 370350
rect 408918 370170 408974 370226
rect 409042 370170 409098 370226
rect 408918 370046 408974 370102
rect 409042 370046 409098 370102
rect 408918 369922 408974 369978
rect 409042 369922 409098 369978
rect 178518 364294 178574 364350
rect 178642 364294 178698 364350
rect 178518 364170 178574 364226
rect 178642 364170 178698 364226
rect 178518 364046 178574 364102
rect 178642 364046 178698 364102
rect 178518 363922 178574 363978
rect 178642 363922 178698 363978
rect 209238 364294 209294 364350
rect 209362 364294 209418 364350
rect 209238 364170 209294 364226
rect 209362 364170 209418 364226
rect 209238 364046 209294 364102
rect 209362 364046 209418 364102
rect 209238 363922 209294 363978
rect 209362 363922 209418 363978
rect 239958 364294 240014 364350
rect 240082 364294 240138 364350
rect 239958 364170 240014 364226
rect 240082 364170 240138 364226
rect 239958 364046 240014 364102
rect 240082 364046 240138 364102
rect 239958 363922 240014 363978
rect 240082 363922 240138 363978
rect 270678 364294 270734 364350
rect 270802 364294 270858 364350
rect 270678 364170 270734 364226
rect 270802 364170 270858 364226
rect 270678 364046 270734 364102
rect 270802 364046 270858 364102
rect 270678 363922 270734 363978
rect 270802 363922 270858 363978
rect 301398 364294 301454 364350
rect 301522 364294 301578 364350
rect 301398 364170 301454 364226
rect 301522 364170 301578 364226
rect 301398 364046 301454 364102
rect 301522 364046 301578 364102
rect 301398 363922 301454 363978
rect 301522 363922 301578 363978
rect 332118 364294 332174 364350
rect 332242 364294 332298 364350
rect 332118 364170 332174 364226
rect 332242 364170 332298 364226
rect 332118 364046 332174 364102
rect 332242 364046 332298 364102
rect 332118 363922 332174 363978
rect 332242 363922 332298 363978
rect 362838 364294 362894 364350
rect 362962 364294 363018 364350
rect 362838 364170 362894 364226
rect 362962 364170 363018 364226
rect 362838 364046 362894 364102
rect 362962 364046 363018 364102
rect 362838 363922 362894 363978
rect 362962 363922 363018 363978
rect 393558 364294 393614 364350
rect 393682 364294 393738 364350
rect 393558 364170 393614 364226
rect 393682 364170 393738 364226
rect 393558 364046 393614 364102
rect 393682 364046 393738 364102
rect 393558 363922 393614 363978
rect 393682 363922 393738 363978
rect 193878 352294 193934 352350
rect 194002 352294 194058 352350
rect 193878 352170 193934 352226
rect 194002 352170 194058 352226
rect 193878 352046 193934 352102
rect 194002 352046 194058 352102
rect 193878 351922 193934 351978
rect 194002 351922 194058 351978
rect 224598 352294 224654 352350
rect 224722 352294 224778 352350
rect 224598 352170 224654 352226
rect 224722 352170 224778 352226
rect 224598 352046 224654 352102
rect 224722 352046 224778 352102
rect 224598 351922 224654 351978
rect 224722 351922 224778 351978
rect 255318 352294 255374 352350
rect 255442 352294 255498 352350
rect 255318 352170 255374 352226
rect 255442 352170 255498 352226
rect 255318 352046 255374 352102
rect 255442 352046 255498 352102
rect 255318 351922 255374 351978
rect 255442 351922 255498 351978
rect 286038 352294 286094 352350
rect 286162 352294 286218 352350
rect 286038 352170 286094 352226
rect 286162 352170 286218 352226
rect 286038 352046 286094 352102
rect 286162 352046 286218 352102
rect 286038 351922 286094 351978
rect 286162 351922 286218 351978
rect 316758 352294 316814 352350
rect 316882 352294 316938 352350
rect 316758 352170 316814 352226
rect 316882 352170 316938 352226
rect 316758 352046 316814 352102
rect 316882 352046 316938 352102
rect 316758 351922 316814 351978
rect 316882 351922 316938 351978
rect 347478 352294 347534 352350
rect 347602 352294 347658 352350
rect 347478 352170 347534 352226
rect 347602 352170 347658 352226
rect 347478 352046 347534 352102
rect 347602 352046 347658 352102
rect 347478 351922 347534 351978
rect 347602 351922 347658 351978
rect 378198 352294 378254 352350
rect 378322 352294 378378 352350
rect 378198 352170 378254 352226
rect 378322 352170 378378 352226
rect 378198 352046 378254 352102
rect 378322 352046 378378 352102
rect 378198 351922 378254 351978
rect 378322 351922 378378 351978
rect 408918 352294 408974 352350
rect 409042 352294 409098 352350
rect 408918 352170 408974 352226
rect 409042 352170 409098 352226
rect 408918 352046 408974 352102
rect 409042 352046 409098 352102
rect 408918 351922 408974 351978
rect 409042 351922 409098 351978
rect 178518 346294 178574 346350
rect 178642 346294 178698 346350
rect 178518 346170 178574 346226
rect 178642 346170 178698 346226
rect 178518 346046 178574 346102
rect 178642 346046 178698 346102
rect 178518 345922 178574 345978
rect 178642 345922 178698 345978
rect 209238 346294 209294 346350
rect 209362 346294 209418 346350
rect 209238 346170 209294 346226
rect 209362 346170 209418 346226
rect 209238 346046 209294 346102
rect 209362 346046 209418 346102
rect 209238 345922 209294 345978
rect 209362 345922 209418 345978
rect 239958 346294 240014 346350
rect 240082 346294 240138 346350
rect 239958 346170 240014 346226
rect 240082 346170 240138 346226
rect 239958 346046 240014 346102
rect 240082 346046 240138 346102
rect 239958 345922 240014 345978
rect 240082 345922 240138 345978
rect 270678 346294 270734 346350
rect 270802 346294 270858 346350
rect 270678 346170 270734 346226
rect 270802 346170 270858 346226
rect 270678 346046 270734 346102
rect 270802 346046 270858 346102
rect 270678 345922 270734 345978
rect 270802 345922 270858 345978
rect 301398 346294 301454 346350
rect 301522 346294 301578 346350
rect 301398 346170 301454 346226
rect 301522 346170 301578 346226
rect 301398 346046 301454 346102
rect 301522 346046 301578 346102
rect 301398 345922 301454 345978
rect 301522 345922 301578 345978
rect 332118 346294 332174 346350
rect 332242 346294 332298 346350
rect 332118 346170 332174 346226
rect 332242 346170 332298 346226
rect 332118 346046 332174 346102
rect 332242 346046 332298 346102
rect 332118 345922 332174 345978
rect 332242 345922 332298 345978
rect 362838 346294 362894 346350
rect 362962 346294 363018 346350
rect 362838 346170 362894 346226
rect 362962 346170 363018 346226
rect 362838 346046 362894 346102
rect 362962 346046 363018 346102
rect 362838 345922 362894 345978
rect 362962 345922 363018 345978
rect 393558 346294 393614 346350
rect 393682 346294 393738 346350
rect 393558 346170 393614 346226
rect 393682 346170 393738 346226
rect 393558 346046 393614 346102
rect 393682 346046 393738 346102
rect 393558 345922 393614 345978
rect 393682 345922 393738 345978
rect 173852 304082 173908 304138
rect 193878 334294 193934 334350
rect 194002 334294 194058 334350
rect 193878 334170 193934 334226
rect 194002 334170 194058 334226
rect 193878 334046 193934 334102
rect 194002 334046 194058 334102
rect 193878 333922 193934 333978
rect 194002 333922 194058 333978
rect 224598 334294 224654 334350
rect 224722 334294 224778 334350
rect 224598 334170 224654 334226
rect 224722 334170 224778 334226
rect 224598 334046 224654 334102
rect 224722 334046 224778 334102
rect 224598 333922 224654 333978
rect 224722 333922 224778 333978
rect 255318 334294 255374 334350
rect 255442 334294 255498 334350
rect 255318 334170 255374 334226
rect 255442 334170 255498 334226
rect 255318 334046 255374 334102
rect 255442 334046 255498 334102
rect 255318 333922 255374 333978
rect 255442 333922 255498 333978
rect 286038 334294 286094 334350
rect 286162 334294 286218 334350
rect 286038 334170 286094 334226
rect 286162 334170 286218 334226
rect 286038 334046 286094 334102
rect 286162 334046 286218 334102
rect 286038 333922 286094 333978
rect 286162 333922 286218 333978
rect 316758 334294 316814 334350
rect 316882 334294 316938 334350
rect 316758 334170 316814 334226
rect 316882 334170 316938 334226
rect 316758 334046 316814 334102
rect 316882 334046 316938 334102
rect 316758 333922 316814 333978
rect 316882 333922 316938 333978
rect 347478 334294 347534 334350
rect 347602 334294 347658 334350
rect 347478 334170 347534 334226
rect 347602 334170 347658 334226
rect 347478 334046 347534 334102
rect 347602 334046 347658 334102
rect 347478 333922 347534 333978
rect 347602 333922 347658 333978
rect 378198 334294 378254 334350
rect 378322 334294 378378 334350
rect 378198 334170 378254 334226
rect 378322 334170 378378 334226
rect 378198 334046 378254 334102
rect 378322 334046 378378 334102
rect 378198 333922 378254 333978
rect 378322 333922 378378 333978
rect 408918 334294 408974 334350
rect 409042 334294 409098 334350
rect 408918 334170 408974 334226
rect 409042 334170 409098 334226
rect 408918 334046 408974 334102
rect 409042 334046 409098 334102
rect 408918 333922 408974 333978
rect 409042 333922 409098 333978
rect 178518 328294 178574 328350
rect 178642 328294 178698 328350
rect 178518 328170 178574 328226
rect 178642 328170 178698 328226
rect 178518 328046 178574 328102
rect 178642 328046 178698 328102
rect 178518 327922 178574 327978
rect 178642 327922 178698 327978
rect 209238 328294 209294 328350
rect 209362 328294 209418 328350
rect 209238 328170 209294 328226
rect 209362 328170 209418 328226
rect 209238 328046 209294 328102
rect 209362 328046 209418 328102
rect 209238 327922 209294 327978
rect 209362 327922 209418 327978
rect 239958 328294 240014 328350
rect 240082 328294 240138 328350
rect 239958 328170 240014 328226
rect 240082 328170 240138 328226
rect 239958 328046 240014 328102
rect 240082 328046 240138 328102
rect 239958 327922 240014 327978
rect 240082 327922 240138 327978
rect 270678 328294 270734 328350
rect 270802 328294 270858 328350
rect 270678 328170 270734 328226
rect 270802 328170 270858 328226
rect 270678 328046 270734 328102
rect 270802 328046 270858 328102
rect 270678 327922 270734 327978
rect 270802 327922 270858 327978
rect 301398 328294 301454 328350
rect 301522 328294 301578 328350
rect 301398 328170 301454 328226
rect 301522 328170 301578 328226
rect 301398 328046 301454 328102
rect 301522 328046 301578 328102
rect 301398 327922 301454 327978
rect 301522 327922 301578 327978
rect 332118 328294 332174 328350
rect 332242 328294 332298 328350
rect 332118 328170 332174 328226
rect 332242 328170 332298 328226
rect 332118 328046 332174 328102
rect 332242 328046 332298 328102
rect 332118 327922 332174 327978
rect 332242 327922 332298 327978
rect 362838 328294 362894 328350
rect 362962 328294 363018 328350
rect 362838 328170 362894 328226
rect 362962 328170 363018 328226
rect 362838 328046 362894 328102
rect 362962 328046 363018 328102
rect 362838 327922 362894 327978
rect 362962 327922 363018 327978
rect 393558 328294 393614 328350
rect 393682 328294 393738 328350
rect 393558 328170 393614 328226
rect 393682 328170 393738 328226
rect 393558 328046 393614 328102
rect 393682 328046 393738 328102
rect 393558 327922 393614 327978
rect 393682 327922 393738 327978
rect 193878 316294 193934 316350
rect 194002 316294 194058 316350
rect 193878 316170 193934 316226
rect 194002 316170 194058 316226
rect 193878 316046 193934 316102
rect 194002 316046 194058 316102
rect 193878 315922 193934 315978
rect 194002 315922 194058 315978
rect 224598 316294 224654 316350
rect 224722 316294 224778 316350
rect 224598 316170 224654 316226
rect 224722 316170 224778 316226
rect 224598 316046 224654 316102
rect 224722 316046 224778 316102
rect 224598 315922 224654 315978
rect 224722 315922 224778 315978
rect 255318 316294 255374 316350
rect 255442 316294 255498 316350
rect 255318 316170 255374 316226
rect 255442 316170 255498 316226
rect 255318 316046 255374 316102
rect 255442 316046 255498 316102
rect 255318 315922 255374 315978
rect 255442 315922 255498 315978
rect 286038 316294 286094 316350
rect 286162 316294 286218 316350
rect 286038 316170 286094 316226
rect 286162 316170 286218 316226
rect 286038 316046 286094 316102
rect 286162 316046 286218 316102
rect 286038 315922 286094 315978
rect 286162 315922 286218 315978
rect 316758 316294 316814 316350
rect 316882 316294 316938 316350
rect 316758 316170 316814 316226
rect 316882 316170 316938 316226
rect 316758 316046 316814 316102
rect 316882 316046 316938 316102
rect 316758 315922 316814 315978
rect 316882 315922 316938 315978
rect 347478 316294 347534 316350
rect 347602 316294 347658 316350
rect 347478 316170 347534 316226
rect 347602 316170 347658 316226
rect 347478 316046 347534 316102
rect 347602 316046 347658 316102
rect 347478 315922 347534 315978
rect 347602 315922 347658 315978
rect 378198 316294 378254 316350
rect 378322 316294 378378 316350
rect 378198 316170 378254 316226
rect 378322 316170 378378 316226
rect 378198 316046 378254 316102
rect 378322 316046 378378 316102
rect 378198 315922 378254 315978
rect 378322 315922 378378 315978
rect 408918 316294 408974 316350
rect 409042 316294 409098 316350
rect 408918 316170 408974 316226
rect 409042 316170 409098 316226
rect 408918 316046 408974 316102
rect 409042 316046 409098 316102
rect 408918 315922 408974 315978
rect 409042 315922 409098 315978
rect 272188 304082 272244 304138
rect 228732 301562 228788 301618
rect 218428 301202 218484 301258
rect 229180 301382 229236 301438
rect 260540 301022 260596 301078
rect 242172 300842 242228 300898
rect 237692 300122 237748 300178
rect 217980 299942 218036 299998
rect 223356 299762 223412 299818
rect 178518 292294 178574 292350
rect 178642 292294 178698 292350
rect 178518 292170 178574 292226
rect 178642 292170 178698 292226
rect 178518 292046 178574 292102
rect 178642 292046 178698 292102
rect 178518 291922 178574 291978
rect 178642 291922 178698 291978
rect 209238 292294 209294 292350
rect 209362 292294 209418 292350
rect 209238 292170 209294 292226
rect 209362 292170 209418 292226
rect 209238 292046 209294 292102
rect 209362 292046 209418 292102
rect 209238 291922 209294 291978
rect 209362 291922 209418 291978
rect 239958 292294 240014 292350
rect 240082 292294 240138 292350
rect 239958 292170 240014 292226
rect 240082 292170 240138 292226
rect 239958 292046 240014 292102
rect 240082 292046 240138 292102
rect 239958 291922 240014 291978
rect 240082 291922 240138 291978
rect 270678 292294 270734 292350
rect 270802 292294 270858 292350
rect 270678 292170 270734 292226
rect 270802 292170 270858 292226
rect 270678 292046 270734 292102
rect 270802 292046 270858 292102
rect 270678 291922 270734 291978
rect 270802 291922 270858 291978
rect 281994 292294 282050 292350
rect 282118 292294 282174 292350
rect 282242 292294 282298 292350
rect 282366 292294 282422 292350
rect 281994 292170 282050 292226
rect 282118 292170 282174 292226
rect 282242 292170 282298 292226
rect 282366 292170 282422 292226
rect 281994 292046 282050 292102
rect 282118 292046 282174 292102
rect 282242 292046 282298 292102
rect 282366 292046 282422 292102
rect 281994 291922 282050 291978
rect 282118 291922 282174 291978
rect 282242 291922 282298 291978
rect 282366 291922 282422 291978
rect 193878 280294 193934 280350
rect 194002 280294 194058 280350
rect 193878 280170 193934 280226
rect 194002 280170 194058 280226
rect 193878 280046 193934 280102
rect 194002 280046 194058 280102
rect 193878 279922 193934 279978
rect 194002 279922 194058 279978
rect 224598 280294 224654 280350
rect 224722 280294 224778 280350
rect 224598 280170 224654 280226
rect 224722 280170 224778 280226
rect 224598 280046 224654 280102
rect 224722 280046 224778 280102
rect 224598 279922 224654 279978
rect 224722 279922 224778 279978
rect 255318 280294 255374 280350
rect 255442 280294 255498 280350
rect 255318 280170 255374 280226
rect 255442 280170 255498 280226
rect 255318 280046 255374 280102
rect 255442 280046 255498 280102
rect 255318 279922 255374 279978
rect 255442 279922 255498 279978
rect 178518 274294 178574 274350
rect 178642 274294 178698 274350
rect 178518 274170 178574 274226
rect 178642 274170 178698 274226
rect 178518 274046 178574 274102
rect 178642 274046 178698 274102
rect 178518 273922 178574 273978
rect 178642 273922 178698 273978
rect 209238 274294 209294 274350
rect 209362 274294 209418 274350
rect 209238 274170 209294 274226
rect 209362 274170 209418 274226
rect 209238 274046 209294 274102
rect 209362 274046 209418 274102
rect 209238 273922 209294 273978
rect 209362 273922 209418 273978
rect 239958 274294 240014 274350
rect 240082 274294 240138 274350
rect 239958 274170 240014 274226
rect 240082 274170 240138 274226
rect 239958 274046 240014 274102
rect 240082 274046 240138 274102
rect 239958 273922 240014 273978
rect 240082 273922 240138 273978
rect 270678 274294 270734 274350
rect 270802 274294 270858 274350
rect 270678 274170 270734 274226
rect 270802 274170 270858 274226
rect 270678 274046 270734 274102
rect 270802 274046 270858 274102
rect 270678 273922 270734 273978
rect 270802 273922 270858 273978
rect 193878 262294 193934 262350
rect 194002 262294 194058 262350
rect 193878 262170 193934 262226
rect 194002 262170 194058 262226
rect 193878 262046 193934 262102
rect 194002 262046 194058 262102
rect 193878 261922 193934 261978
rect 194002 261922 194058 261978
rect 224598 262294 224654 262350
rect 224722 262294 224778 262350
rect 224598 262170 224654 262226
rect 224722 262170 224778 262226
rect 224598 262046 224654 262102
rect 224722 262046 224778 262102
rect 224598 261922 224654 261978
rect 224722 261922 224778 261978
rect 255318 262294 255374 262350
rect 255442 262294 255498 262350
rect 255318 262170 255374 262226
rect 255442 262170 255498 262226
rect 255318 262046 255374 262102
rect 255442 262046 255498 262102
rect 255318 261922 255374 261978
rect 255442 261922 255498 261978
rect 178518 256294 178574 256350
rect 178642 256294 178698 256350
rect 178518 256170 178574 256226
rect 178642 256170 178698 256226
rect 178518 256046 178574 256102
rect 178642 256046 178698 256102
rect 178518 255922 178574 255978
rect 178642 255922 178698 255978
rect 209238 256294 209294 256350
rect 209362 256294 209418 256350
rect 209238 256170 209294 256226
rect 209362 256170 209418 256226
rect 209238 256046 209294 256102
rect 209362 256046 209418 256102
rect 209238 255922 209294 255978
rect 209362 255922 209418 255978
rect 239958 256294 240014 256350
rect 240082 256294 240138 256350
rect 239958 256170 240014 256226
rect 240082 256170 240138 256226
rect 239958 256046 240014 256102
rect 240082 256046 240138 256102
rect 239958 255922 240014 255978
rect 240082 255922 240138 255978
rect 270678 256294 270734 256350
rect 270802 256294 270858 256350
rect 270678 256170 270734 256226
rect 270802 256170 270858 256226
rect 270678 256046 270734 256102
rect 270802 256046 270858 256102
rect 270678 255922 270734 255978
rect 270802 255922 270858 255978
rect 193878 244294 193934 244350
rect 194002 244294 194058 244350
rect 193878 244170 193934 244226
rect 194002 244170 194058 244226
rect 193878 244046 193934 244102
rect 194002 244046 194058 244102
rect 193878 243922 193934 243978
rect 194002 243922 194058 243978
rect 224598 244294 224654 244350
rect 224722 244294 224778 244350
rect 224598 244170 224654 244226
rect 224722 244170 224778 244226
rect 224598 244046 224654 244102
rect 224722 244046 224778 244102
rect 224598 243922 224654 243978
rect 224722 243922 224778 243978
rect 255318 244294 255374 244350
rect 255442 244294 255498 244350
rect 255318 244170 255374 244226
rect 255442 244170 255498 244226
rect 255318 244046 255374 244102
rect 255442 244046 255498 244102
rect 255318 243922 255374 243978
rect 255442 243922 255498 243978
rect 178518 238294 178574 238350
rect 178642 238294 178698 238350
rect 178518 238170 178574 238226
rect 178642 238170 178698 238226
rect 178518 238046 178574 238102
rect 178642 238046 178698 238102
rect 178518 237922 178574 237978
rect 178642 237922 178698 237978
rect 209238 238294 209294 238350
rect 209362 238294 209418 238350
rect 209238 238170 209294 238226
rect 209362 238170 209418 238226
rect 209238 238046 209294 238102
rect 209362 238046 209418 238102
rect 209238 237922 209294 237978
rect 209362 237922 209418 237978
rect 239958 238294 240014 238350
rect 240082 238294 240138 238350
rect 239958 238170 240014 238226
rect 240082 238170 240138 238226
rect 239958 238046 240014 238102
rect 240082 238046 240138 238102
rect 239958 237922 240014 237978
rect 240082 237922 240138 237978
rect 270678 238294 270734 238350
rect 270802 238294 270858 238350
rect 270678 238170 270734 238226
rect 270802 238170 270858 238226
rect 270678 238046 270734 238102
rect 270802 238046 270858 238102
rect 270678 237922 270734 237978
rect 270802 237922 270858 237978
rect 193878 226294 193934 226350
rect 194002 226294 194058 226350
rect 193878 226170 193934 226226
rect 194002 226170 194058 226226
rect 193878 226046 193934 226102
rect 194002 226046 194058 226102
rect 193878 225922 193934 225978
rect 194002 225922 194058 225978
rect 224598 226294 224654 226350
rect 224722 226294 224778 226350
rect 224598 226170 224654 226226
rect 224722 226170 224778 226226
rect 224598 226046 224654 226102
rect 224722 226046 224778 226102
rect 224598 225922 224654 225978
rect 224722 225922 224778 225978
rect 255318 226294 255374 226350
rect 255442 226294 255498 226350
rect 255318 226170 255374 226226
rect 255442 226170 255498 226226
rect 255318 226046 255374 226102
rect 255442 226046 255498 226102
rect 255318 225922 255374 225978
rect 255442 225922 255498 225978
rect 178518 220294 178574 220350
rect 178642 220294 178698 220350
rect 178518 220170 178574 220226
rect 178642 220170 178698 220226
rect 178518 220046 178574 220102
rect 178642 220046 178698 220102
rect 178518 219922 178574 219978
rect 178642 219922 178698 219978
rect 209238 220294 209294 220350
rect 209362 220294 209418 220350
rect 209238 220170 209294 220226
rect 209362 220170 209418 220226
rect 209238 220046 209294 220102
rect 209362 220046 209418 220102
rect 209238 219922 209294 219978
rect 209362 219922 209418 219978
rect 239958 220294 240014 220350
rect 240082 220294 240138 220350
rect 239958 220170 240014 220226
rect 240082 220170 240138 220226
rect 239958 220046 240014 220102
rect 240082 220046 240138 220102
rect 239958 219922 240014 219978
rect 240082 219922 240138 219978
rect 270678 220294 270734 220350
rect 270802 220294 270858 220350
rect 270678 220170 270734 220226
rect 270802 220170 270858 220226
rect 270678 220046 270734 220102
rect 270802 220046 270858 220102
rect 270678 219922 270734 219978
rect 270802 219922 270858 219978
rect 193878 208294 193934 208350
rect 194002 208294 194058 208350
rect 193878 208170 193934 208226
rect 194002 208170 194058 208226
rect 193878 208046 193934 208102
rect 194002 208046 194058 208102
rect 193878 207922 193934 207978
rect 194002 207922 194058 207978
rect 224598 208294 224654 208350
rect 224722 208294 224778 208350
rect 224598 208170 224654 208226
rect 224722 208170 224778 208226
rect 224598 208046 224654 208102
rect 224722 208046 224778 208102
rect 224598 207922 224654 207978
rect 224722 207922 224778 207978
rect 255318 208294 255374 208350
rect 255442 208294 255498 208350
rect 255318 208170 255374 208226
rect 255442 208170 255498 208226
rect 255318 208046 255374 208102
rect 255442 208046 255498 208102
rect 255318 207922 255374 207978
rect 255442 207922 255498 207978
rect 178518 202294 178574 202350
rect 178642 202294 178698 202350
rect 178518 202170 178574 202226
rect 178642 202170 178698 202226
rect 178518 202046 178574 202102
rect 178642 202046 178698 202102
rect 178518 201922 178574 201978
rect 178642 201922 178698 201978
rect 209238 202294 209294 202350
rect 209362 202294 209418 202350
rect 209238 202170 209294 202226
rect 209362 202170 209418 202226
rect 209238 202046 209294 202102
rect 209362 202046 209418 202102
rect 209238 201922 209294 201978
rect 209362 201922 209418 201978
rect 239958 202294 240014 202350
rect 240082 202294 240138 202350
rect 239958 202170 240014 202226
rect 240082 202170 240138 202226
rect 239958 202046 240014 202102
rect 240082 202046 240138 202102
rect 239958 201922 240014 201978
rect 240082 201922 240138 201978
rect 270678 202294 270734 202350
rect 270802 202294 270858 202350
rect 270678 202170 270734 202226
rect 270802 202170 270858 202226
rect 270678 202046 270734 202102
rect 270802 202046 270858 202102
rect 270678 201922 270734 201978
rect 270802 201922 270858 201978
rect 193878 190294 193934 190350
rect 194002 190294 194058 190350
rect 193878 190170 193934 190226
rect 194002 190170 194058 190226
rect 193878 190046 193934 190102
rect 194002 190046 194058 190102
rect 193878 189922 193934 189978
rect 194002 189922 194058 189978
rect 224598 190294 224654 190350
rect 224722 190294 224778 190350
rect 224598 190170 224654 190226
rect 224722 190170 224778 190226
rect 224598 190046 224654 190102
rect 224722 190046 224778 190102
rect 224598 189922 224654 189978
rect 224722 189922 224778 189978
rect 255318 190294 255374 190350
rect 255442 190294 255498 190350
rect 255318 190170 255374 190226
rect 255442 190170 255498 190226
rect 255318 190046 255374 190102
rect 255442 190046 255498 190102
rect 255318 189922 255374 189978
rect 255442 189922 255498 189978
rect 178518 184294 178574 184350
rect 178642 184294 178698 184350
rect 178518 184170 178574 184226
rect 178642 184170 178698 184226
rect 178518 184046 178574 184102
rect 178642 184046 178698 184102
rect 178518 183922 178574 183978
rect 178642 183922 178698 183978
rect 209238 184294 209294 184350
rect 209362 184294 209418 184350
rect 209238 184170 209294 184226
rect 209362 184170 209418 184226
rect 209238 184046 209294 184102
rect 209362 184046 209418 184102
rect 209238 183922 209294 183978
rect 209362 183922 209418 183978
rect 239958 184294 240014 184350
rect 240082 184294 240138 184350
rect 239958 184170 240014 184226
rect 240082 184170 240138 184226
rect 239958 184046 240014 184102
rect 240082 184046 240138 184102
rect 239958 183922 240014 183978
rect 240082 183922 240138 183978
rect 270678 184294 270734 184350
rect 270802 184294 270858 184350
rect 270678 184170 270734 184226
rect 270802 184170 270858 184226
rect 270678 184046 270734 184102
rect 270802 184046 270858 184102
rect 270678 183922 270734 183978
rect 270802 183922 270858 183978
rect 193878 172294 193934 172350
rect 194002 172294 194058 172350
rect 193878 172170 193934 172226
rect 194002 172170 194058 172226
rect 193878 172046 193934 172102
rect 194002 172046 194058 172102
rect 193878 171922 193934 171978
rect 194002 171922 194058 171978
rect 224598 172294 224654 172350
rect 224722 172294 224778 172350
rect 224598 172170 224654 172226
rect 224722 172170 224778 172226
rect 224598 172046 224654 172102
rect 224722 172046 224778 172102
rect 224598 171922 224654 171978
rect 224722 171922 224778 171978
rect 255318 172294 255374 172350
rect 255442 172294 255498 172350
rect 255318 172170 255374 172226
rect 255442 172170 255498 172226
rect 255318 172046 255374 172102
rect 255442 172046 255498 172102
rect 255318 171922 255374 171978
rect 255442 171922 255498 171978
rect 178518 166294 178574 166350
rect 178642 166294 178698 166350
rect 178518 166170 178574 166226
rect 178642 166170 178698 166226
rect 178518 166046 178574 166102
rect 178642 166046 178698 166102
rect 178518 165922 178574 165978
rect 178642 165922 178698 165978
rect 209238 166294 209294 166350
rect 209362 166294 209418 166350
rect 209238 166170 209294 166226
rect 209362 166170 209418 166226
rect 209238 166046 209294 166102
rect 209362 166046 209418 166102
rect 209238 165922 209294 165978
rect 209362 165922 209418 165978
rect 239958 166294 240014 166350
rect 240082 166294 240138 166350
rect 239958 166170 240014 166226
rect 240082 166170 240138 166226
rect 239958 166046 240014 166102
rect 240082 166046 240138 166102
rect 239958 165922 240014 165978
rect 240082 165922 240138 165978
rect 270678 166294 270734 166350
rect 270802 166294 270858 166350
rect 270678 166170 270734 166226
rect 270802 166170 270858 166226
rect 270678 166046 270734 166102
rect 270802 166046 270858 166102
rect 270678 165922 270734 165978
rect 270802 165922 270858 165978
rect 193878 154294 193934 154350
rect 194002 154294 194058 154350
rect 193878 154170 193934 154226
rect 194002 154170 194058 154226
rect 193878 154046 193934 154102
rect 194002 154046 194058 154102
rect 193878 153922 193934 153978
rect 194002 153922 194058 153978
rect 224598 154294 224654 154350
rect 224722 154294 224778 154350
rect 224598 154170 224654 154226
rect 224722 154170 224778 154226
rect 224598 154046 224654 154102
rect 224722 154046 224778 154102
rect 224598 153922 224654 153978
rect 224722 153922 224778 153978
rect 255318 154294 255374 154350
rect 255442 154294 255498 154350
rect 255318 154170 255374 154226
rect 255442 154170 255498 154226
rect 255318 154046 255374 154102
rect 255442 154046 255498 154102
rect 255318 153922 255374 153978
rect 255442 153922 255498 153978
rect 178518 148294 178574 148350
rect 178642 148294 178698 148350
rect 178518 148170 178574 148226
rect 178642 148170 178698 148226
rect 178518 148046 178574 148102
rect 178642 148046 178698 148102
rect 178518 147922 178574 147978
rect 178642 147922 178698 147978
rect 209238 148294 209294 148350
rect 209362 148294 209418 148350
rect 209238 148170 209294 148226
rect 209362 148170 209418 148226
rect 209238 148046 209294 148102
rect 209362 148046 209418 148102
rect 209238 147922 209294 147978
rect 209362 147922 209418 147978
rect 239958 148294 240014 148350
rect 240082 148294 240138 148350
rect 239958 148170 240014 148226
rect 240082 148170 240138 148226
rect 239958 148046 240014 148102
rect 240082 148046 240138 148102
rect 239958 147922 240014 147978
rect 240082 147922 240138 147978
rect 270678 148294 270734 148350
rect 270802 148294 270858 148350
rect 270678 148170 270734 148226
rect 270802 148170 270858 148226
rect 270678 148046 270734 148102
rect 270802 148046 270858 148102
rect 270678 147922 270734 147978
rect 270802 147922 270858 147978
rect 193878 136294 193934 136350
rect 194002 136294 194058 136350
rect 193878 136170 193934 136226
rect 194002 136170 194058 136226
rect 193878 136046 193934 136102
rect 194002 136046 194058 136102
rect 193878 135922 193934 135978
rect 194002 135922 194058 135978
rect 224598 136294 224654 136350
rect 224722 136294 224778 136350
rect 224598 136170 224654 136226
rect 224722 136170 224778 136226
rect 224598 136046 224654 136102
rect 224722 136046 224778 136102
rect 224598 135922 224654 135978
rect 224722 135922 224778 135978
rect 255318 136294 255374 136350
rect 255442 136294 255498 136350
rect 255318 136170 255374 136226
rect 255442 136170 255498 136226
rect 255318 136046 255374 136102
rect 255442 136046 255498 136102
rect 255318 135922 255374 135978
rect 255442 135922 255498 135978
rect 178518 130294 178574 130350
rect 178642 130294 178698 130350
rect 178518 130170 178574 130226
rect 178642 130170 178698 130226
rect 178518 130046 178574 130102
rect 178642 130046 178698 130102
rect 178518 129922 178574 129978
rect 178642 129922 178698 129978
rect 209238 130294 209294 130350
rect 209362 130294 209418 130350
rect 209238 130170 209294 130226
rect 209362 130170 209418 130226
rect 209238 130046 209294 130102
rect 209362 130046 209418 130102
rect 209238 129922 209294 129978
rect 209362 129922 209418 129978
rect 239958 130294 240014 130350
rect 240082 130294 240138 130350
rect 239958 130170 240014 130226
rect 240082 130170 240138 130226
rect 239958 130046 240014 130102
rect 240082 130046 240138 130102
rect 239958 129922 240014 129978
rect 240082 129922 240138 129978
rect 270678 130294 270734 130350
rect 270802 130294 270858 130350
rect 270678 130170 270734 130226
rect 270802 130170 270858 130226
rect 270678 130046 270734 130102
rect 270802 130046 270858 130102
rect 270678 129922 270734 129978
rect 270802 129922 270858 129978
rect 193878 118294 193934 118350
rect 194002 118294 194058 118350
rect 193878 118170 193934 118226
rect 194002 118170 194058 118226
rect 193878 118046 193934 118102
rect 194002 118046 194058 118102
rect 193878 117922 193934 117978
rect 194002 117922 194058 117978
rect 224598 118294 224654 118350
rect 224722 118294 224778 118350
rect 224598 118170 224654 118226
rect 224722 118170 224778 118226
rect 224598 118046 224654 118102
rect 224722 118046 224778 118102
rect 224598 117922 224654 117978
rect 224722 117922 224778 117978
rect 255318 118294 255374 118350
rect 255442 118294 255498 118350
rect 255318 118170 255374 118226
rect 255442 118170 255498 118226
rect 255318 118046 255374 118102
rect 255442 118046 255498 118102
rect 255318 117922 255374 117978
rect 255442 117922 255498 117978
rect 178518 112294 178574 112350
rect 178642 112294 178698 112350
rect 178518 112170 178574 112226
rect 178642 112170 178698 112226
rect 178518 112046 178574 112102
rect 178642 112046 178698 112102
rect 178518 111922 178574 111978
rect 178642 111922 178698 111978
rect 209238 112294 209294 112350
rect 209362 112294 209418 112350
rect 209238 112170 209294 112226
rect 209362 112170 209418 112226
rect 209238 112046 209294 112102
rect 209362 112046 209418 112102
rect 209238 111922 209294 111978
rect 209362 111922 209418 111978
rect 239958 112294 240014 112350
rect 240082 112294 240138 112350
rect 239958 112170 240014 112226
rect 240082 112170 240138 112226
rect 239958 112046 240014 112102
rect 240082 112046 240138 112102
rect 239958 111922 240014 111978
rect 240082 111922 240138 111978
rect 270678 112294 270734 112350
rect 270802 112294 270858 112350
rect 270678 112170 270734 112226
rect 270802 112170 270858 112226
rect 270678 112046 270734 112102
rect 270802 112046 270858 112102
rect 270678 111922 270734 111978
rect 270802 111922 270858 111978
rect 271516 108242 271572 108298
rect 189834 94294 189890 94350
rect 189958 94294 190014 94350
rect 190082 94294 190138 94350
rect 190206 94294 190262 94350
rect 189834 94170 189890 94226
rect 189958 94170 190014 94226
rect 190082 94170 190138 94226
rect 190206 94170 190262 94226
rect 189834 94046 189890 94102
rect 189958 94046 190014 94102
rect 190082 94046 190138 94102
rect 190206 94046 190262 94102
rect 189834 93922 189890 93978
rect 189958 93922 190014 93978
rect 190082 93922 190138 93978
rect 190206 93922 190262 93978
rect 189532 86462 189588 86518
rect 181468 81422 181524 81478
rect 189834 76294 189890 76350
rect 189958 76294 190014 76350
rect 190082 76294 190138 76350
rect 190206 76294 190262 76350
rect 189834 76170 189890 76226
rect 189958 76170 190014 76226
rect 190082 76170 190138 76226
rect 190206 76170 190262 76226
rect 189834 76046 189890 76102
rect 189958 76046 190014 76102
rect 190082 76046 190138 76102
rect 190206 76046 190262 76102
rect 189834 75922 189890 75978
rect 189958 75922 190014 75978
rect 190082 75922 190138 75978
rect 190206 75922 190262 75978
rect 193554 99867 193610 99923
rect 193678 99867 193734 99923
rect 193802 99867 193858 99923
rect 193926 99867 193982 99923
rect 243516 101942 243572 101998
rect 226604 101762 226660 101818
rect 220554 94294 220610 94350
rect 220678 94294 220734 94350
rect 220802 94294 220858 94350
rect 220926 94294 220982 94350
rect 220554 94170 220610 94226
rect 220678 94170 220734 94226
rect 220802 94170 220858 94226
rect 220926 94170 220982 94226
rect 220554 94046 220610 94102
rect 220678 94046 220734 94102
rect 220802 94046 220858 94102
rect 220926 94046 220982 94102
rect 220554 93922 220610 93978
rect 220678 93922 220734 93978
rect 220802 93922 220858 93978
rect 220926 93922 220982 93978
rect 206556 88442 206612 88498
rect 193554 82294 193610 82350
rect 193678 82294 193734 82350
rect 193802 82294 193858 82350
rect 193926 82294 193982 82350
rect 193554 82170 193610 82226
rect 193678 82170 193734 82226
rect 193802 82170 193858 82226
rect 193926 82170 193982 82226
rect 193554 82046 193610 82102
rect 193678 82046 193734 82102
rect 193802 82046 193858 82102
rect 193926 82046 193982 82102
rect 193554 81922 193610 81978
rect 193678 81922 193734 81978
rect 193802 81922 193858 81978
rect 193926 81922 193982 81978
rect 202524 88262 202580 88318
rect 204876 88082 204932 88138
rect 213948 85022 214004 85078
rect 214844 84842 214900 84898
rect 220554 76294 220610 76350
rect 220678 76294 220734 76350
rect 220802 76294 220858 76350
rect 220926 76294 220982 76350
rect 220554 76170 220610 76226
rect 220678 76170 220734 76226
rect 220802 76170 220858 76226
rect 220926 76170 220982 76226
rect 220554 76046 220610 76102
rect 220678 76046 220734 76102
rect 220802 76046 220858 76102
rect 220926 76046 220982 76102
rect 220554 75922 220610 75978
rect 220678 75922 220734 75978
rect 220802 75922 220858 75978
rect 220926 75922 220982 75978
rect 224274 99867 224330 99923
rect 224398 99867 224454 99923
rect 224522 99867 224578 99923
rect 224646 99867 224702 99923
rect 224274 82294 224330 82350
rect 224398 82294 224454 82350
rect 224522 82294 224578 82350
rect 224646 82294 224702 82350
rect 224274 82170 224330 82226
rect 224398 82170 224454 82226
rect 224522 82170 224578 82226
rect 224646 82170 224702 82226
rect 224274 82046 224330 82102
rect 224398 82046 224454 82102
rect 224522 82046 224578 82102
rect 224646 82046 224702 82102
rect 224274 81922 224330 81978
rect 224398 81922 224454 81978
rect 224522 81922 224578 81978
rect 224646 81922 224702 81978
rect 226716 101582 226772 101638
rect 235116 98522 235172 98578
rect 233436 98342 233492 98398
rect 230076 98162 230132 98218
rect 228396 96542 228452 96598
rect 229964 92402 230020 92458
rect 232092 89882 232148 89938
rect 241836 96722 241892 96778
rect 234780 80522 234836 80578
rect 236796 94922 236852 94978
rect 238476 93122 238532 93178
rect 267932 104102 267988 104158
rect 251274 94294 251330 94350
rect 251398 94294 251454 94350
rect 251522 94294 251578 94350
rect 251646 94294 251702 94350
rect 251274 94170 251330 94226
rect 251398 94170 251454 94226
rect 251522 94170 251578 94226
rect 251646 94170 251702 94226
rect 251274 94046 251330 94102
rect 251398 94046 251454 94102
rect 251522 94046 251578 94102
rect 251646 94046 251702 94102
rect 251274 93922 251330 93978
rect 251398 93922 251454 93978
rect 251522 93922 251578 93978
rect 251646 93922 251702 93978
rect 245196 91502 245252 91558
rect 249564 89162 249620 89218
rect 246876 87362 246932 87418
rect 229964 80342 230020 80398
rect 231420 80162 231476 80218
rect 230748 79802 230804 79858
rect 232764 79982 232820 80038
rect 227276 78902 227332 78958
rect 250908 78002 250964 78058
rect 254994 99867 255050 99923
rect 255118 99867 255174 99923
rect 255242 99867 255298 99923
rect 255366 99867 255422 99923
rect 254716 91142 254772 91198
rect 253484 90962 253540 91018
rect 251916 90782 251972 90838
rect 252924 80882 252980 80938
rect 254492 82682 254548 82738
rect 254994 82294 255050 82350
rect 255118 82294 255174 82350
rect 255242 82294 255298 82350
rect 255366 82294 255422 82350
rect 254994 82170 255050 82226
rect 255118 82170 255174 82226
rect 255242 82170 255298 82226
rect 255366 82170 255422 82226
rect 254994 82046 255050 82102
rect 255118 82046 255174 82102
rect 255242 82046 255298 82102
rect 255366 82046 255422 82102
rect 254994 81922 255050 81978
rect 255118 81922 255174 81978
rect 255242 81922 255298 81978
rect 255366 81922 255422 81978
rect 251274 76294 251330 76350
rect 251398 76294 251454 76350
rect 251522 76294 251578 76350
rect 251646 76294 251702 76350
rect 251274 76170 251330 76226
rect 251398 76170 251454 76226
rect 251522 76170 251578 76226
rect 251646 76170 251702 76226
rect 251274 76046 251330 76102
rect 251398 76046 251454 76102
rect 251522 76046 251578 76102
rect 251646 76046 251702 76102
rect 251274 75922 251330 75978
rect 251398 75922 251454 75978
rect 251522 75922 251578 75978
rect 251646 75922 251702 75978
rect 259644 89342 259700 89398
rect 256956 80702 257012 80758
rect 185878 64294 185934 64350
rect 186002 64294 186058 64350
rect 185878 64170 185934 64226
rect 186002 64170 186058 64226
rect 185878 64046 185934 64102
rect 186002 64046 186058 64102
rect 185878 63922 185934 63978
rect 186002 63922 186058 63978
rect 216598 64294 216654 64350
rect 216722 64294 216778 64350
rect 216598 64170 216654 64226
rect 216722 64170 216778 64226
rect 216598 64046 216654 64102
rect 216722 64046 216778 64102
rect 216598 63922 216654 63978
rect 216722 63922 216778 63978
rect 247318 64294 247374 64350
rect 247442 64294 247498 64350
rect 247318 64170 247374 64226
rect 247442 64170 247498 64226
rect 247318 64046 247374 64102
rect 247442 64046 247498 64102
rect 247318 63922 247374 63978
rect 247442 63922 247498 63978
rect 170518 58294 170574 58350
rect 170642 58294 170698 58350
rect 170518 58170 170574 58226
rect 170642 58170 170698 58226
rect 170518 58046 170574 58102
rect 170642 58046 170698 58102
rect 170518 57922 170574 57978
rect 170642 57922 170698 57978
rect 201238 58294 201294 58350
rect 201362 58294 201418 58350
rect 201238 58170 201294 58226
rect 201362 58170 201418 58226
rect 201238 58046 201294 58102
rect 201362 58046 201418 58102
rect 201238 57922 201294 57978
rect 201362 57922 201418 57978
rect 231958 58294 232014 58350
rect 232082 58294 232138 58350
rect 231958 58170 232014 58226
rect 232082 58170 232138 58226
rect 231958 58046 232014 58102
rect 232082 58046 232138 58102
rect 231958 57922 232014 57978
rect 232082 57922 232138 57978
rect 262678 58294 262734 58350
rect 262802 58294 262858 58350
rect 262678 58170 262734 58226
rect 262802 58170 262858 58226
rect 262678 58046 262734 58102
rect 262802 58046 262858 58102
rect 262678 57922 262734 57978
rect 262802 57922 262858 57978
rect 264572 54602 264628 54658
rect 185878 46294 185934 46350
rect 186002 46294 186058 46350
rect 185878 46170 185934 46226
rect 186002 46170 186058 46226
rect 185878 46046 185934 46102
rect 186002 46046 186058 46102
rect 185878 45922 185934 45978
rect 186002 45922 186058 45978
rect 216598 46294 216654 46350
rect 216722 46294 216778 46350
rect 216598 46170 216654 46226
rect 216722 46170 216778 46226
rect 216598 46046 216654 46102
rect 216722 46046 216778 46102
rect 216598 45922 216654 45978
rect 216722 45922 216778 45978
rect 247318 46294 247374 46350
rect 247442 46294 247498 46350
rect 247318 46170 247374 46226
rect 247442 46170 247498 46226
rect 247318 46046 247374 46102
rect 247442 46046 247498 46102
rect 247318 45922 247374 45978
rect 247442 45922 247498 45978
rect 170518 40294 170574 40350
rect 170642 40294 170698 40350
rect 170518 40170 170574 40226
rect 170642 40170 170698 40226
rect 170518 40046 170574 40102
rect 170642 40046 170698 40102
rect 170518 39922 170574 39978
rect 170642 39922 170698 39978
rect 201238 40294 201294 40350
rect 201362 40294 201418 40350
rect 201238 40170 201294 40226
rect 201362 40170 201418 40226
rect 201238 40046 201294 40102
rect 201362 40046 201418 40102
rect 201238 39922 201294 39978
rect 201362 39922 201418 39978
rect 231958 40294 232014 40350
rect 232082 40294 232138 40350
rect 231958 40170 232014 40226
rect 232082 40170 232138 40226
rect 231958 40046 232014 40102
rect 232082 40046 232138 40102
rect 231958 39922 232014 39978
rect 232082 39922 232138 39978
rect 262678 40294 262734 40350
rect 262802 40294 262858 40350
rect 262678 40170 262734 40226
rect 262802 40170 262858 40226
rect 262678 40046 262734 40102
rect 262802 40046 262858 40102
rect 262678 39922 262734 39978
rect 262802 39922 262858 39978
rect 185878 28294 185934 28350
rect 186002 28294 186058 28350
rect 185878 28170 185934 28226
rect 186002 28170 186058 28226
rect 185878 28046 185934 28102
rect 186002 28046 186058 28102
rect 185878 27922 185934 27978
rect 186002 27922 186058 27978
rect 216598 28294 216654 28350
rect 216722 28294 216778 28350
rect 216598 28170 216654 28226
rect 216722 28170 216778 28226
rect 216598 28046 216654 28102
rect 216722 28046 216778 28102
rect 216598 27922 216654 27978
rect 216722 27922 216778 27978
rect 247318 28294 247374 28350
rect 247442 28294 247498 28350
rect 247318 28170 247374 28226
rect 247442 28170 247498 28226
rect 247318 28046 247374 28102
rect 247442 28046 247498 28102
rect 247318 27922 247374 27978
rect 247442 27922 247498 27978
rect 170518 22294 170574 22350
rect 170642 22294 170698 22350
rect 170518 22170 170574 22226
rect 170642 22170 170698 22226
rect 170518 22046 170574 22102
rect 170642 22046 170698 22102
rect 170518 21922 170574 21978
rect 170642 21922 170698 21978
rect 201238 22294 201294 22350
rect 201362 22294 201418 22350
rect 201238 22170 201294 22226
rect 201362 22170 201418 22226
rect 201238 22046 201294 22102
rect 201362 22046 201418 22102
rect 201238 21922 201294 21978
rect 201362 21922 201418 21978
rect 231958 22294 232014 22350
rect 232082 22294 232138 22350
rect 231958 22170 232014 22226
rect 232082 22170 232138 22226
rect 231958 22046 232014 22102
rect 232082 22046 232138 22102
rect 231958 21922 232014 21978
rect 232082 21922 232138 21978
rect 262678 22294 262734 22350
rect 262802 22294 262858 22350
rect 262678 22170 262734 22226
rect 262802 22170 262858 22226
rect 262678 22046 262734 22102
rect 262802 22046 262858 22102
rect 262678 21922 262734 21978
rect 262802 21922 262858 21978
rect 241948 21302 242004 21358
rect 240604 21122 240660 21178
rect 240380 20942 240436 20998
rect 231196 19862 231252 19918
rect 169596 13382 169652 13438
rect 187068 13562 187124 13618
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 184940 5822 184996 5878
rect 186172 9242 186228 9298
rect 186844 11762 186900 11818
rect 188188 7442 188244 7498
rect 186508 6002 186564 6058
rect 185052 3302 185108 3358
rect 190540 11942 190596 11998
rect 190428 7622 190484 7678
rect 217308 16100 217364 16138
rect 217308 16082 217364 16100
rect 218652 13562 218708 13618
rect 209692 13412 209748 13438
rect 209692 13382 209748 13412
rect 210140 13412 210196 13438
rect 210140 13382 210196 13412
rect 209916 13202 209972 13258
rect 209468 13022 209524 13078
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 221340 13922 221396 13978
rect 222236 13742 222292 13798
rect 222012 9602 222068 9658
rect 223356 6362 223412 6418
rect 226268 16802 226324 16858
rect 230748 17162 230804 17218
rect 239260 19502 239316 19558
rect 236572 19322 236628 19378
rect 236796 16982 236852 17038
rect 226044 15902 226100 15958
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 226604 8342 226660 8398
rect 225036 6182 225092 6238
rect 224924 6002 224980 6058
rect 228396 7622 228452 7678
rect 231420 9242 231476 9298
rect 236124 11582 236180 11638
rect 241948 19862 242004 19918
rect 243740 19862 243796 19918
rect 241948 19682 242004 19738
rect 245084 17522 245140 17578
rect 245308 16268 245364 16318
rect 245308 16262 245364 16268
rect 238588 15182 238644 15238
rect 230076 7442 230132 7498
rect 238252 7982 238308 8038
rect 231756 6542 231812 6598
rect 226716 5822 226772 5878
rect 238364 2762 238420 2818
rect 243068 14282 243124 14338
rect 240044 2402 240100 2458
rect 238476 782 238532 838
rect 241500 11402 241556 11458
rect 241052 7802 241108 7858
rect 242396 9422 242452 9478
rect 241724 3122 241780 3178
rect 240156 602 240212 658
rect 243292 242 243348 298
rect 245980 12842 246036 12898
rect 243516 11762 243572 11818
rect 245084 4742 245140 4798
rect 246876 4922 246932 4978
rect 245196 3302 245252 3358
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 243404 62 243460 118
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 256956 17162 257012 17218
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 264684 20042 264740 20098
rect 265468 12482 265524 12538
rect 266364 85742 266420 85798
rect 266364 17522 266420 17578
rect 268156 87542 268212 87598
rect 268044 85202 268100 85258
rect 266588 21302 266644 21358
rect 267932 77282 267988 77338
rect 266924 72962 266980 73018
rect 266700 19862 266756 19918
rect 266812 69722 266868 69778
rect 267820 15902 267876 15958
rect 267932 13382 267988 13438
rect 265468 2762 265524 2818
rect 268828 85922 268884 85978
rect 268156 16262 268212 16318
rect 268268 84122 268324 84178
rect 268940 82862 268996 82918
rect 268716 77642 268772 77698
rect 268604 74042 268660 74098
rect 268380 14282 268436 14338
rect 268492 73142 268548 73198
rect 268268 13202 268324 13258
rect 268604 13922 268660 13978
rect 269052 16262 269108 16318
rect 268940 13022 268996 13078
rect 269948 86642 270004 86698
rect 269612 11402 269668 11458
rect 267148 2582 267204 2638
rect 269948 12842 270004 12898
rect 270732 83042 270788 83098
rect 270284 21122 270340 21178
rect 270508 20942 270564 20998
rect 272972 104102 273028 104158
rect 271702 76294 271758 76350
rect 271826 76294 271882 76350
rect 271702 76170 271758 76226
rect 271826 76170 271882 76226
rect 271702 76046 271758 76102
rect 271826 76046 271882 76102
rect 271702 75922 271758 75978
rect 271826 75922 271882 75978
rect 271702 58294 271758 58350
rect 271826 58294 271882 58350
rect 271702 58170 271758 58226
rect 271826 58170 271882 58226
rect 271702 58046 271758 58102
rect 271826 58046 271882 58102
rect 271702 57922 271758 57978
rect 271826 57922 271882 57978
rect 271702 40294 271758 40350
rect 271826 40294 271882 40350
rect 271702 40170 271758 40226
rect 271826 40170 271882 40226
rect 271702 40046 271758 40102
rect 271826 40046 271882 40102
rect 271702 39922 271758 39978
rect 271826 39922 271882 39978
rect 271702 22294 271758 22350
rect 271826 22294 271882 22350
rect 271702 22170 271758 22226
rect 271826 22170 271882 22226
rect 271702 22046 271758 22102
rect 271826 22046 271882 22102
rect 271702 21922 271758 21978
rect 271826 21922 271882 21978
rect 271292 19502 271348 19558
rect 273084 54602 273140 54658
rect 273308 73142 273364 73198
rect 281994 274294 282050 274350
rect 282118 274294 282174 274350
rect 282242 274294 282298 274350
rect 282366 274294 282422 274350
rect 281994 274170 282050 274226
rect 282118 274170 282174 274226
rect 282242 274170 282298 274226
rect 282366 274170 282422 274226
rect 281994 274046 282050 274102
rect 282118 274046 282174 274102
rect 282242 274046 282298 274102
rect 282366 274046 282422 274102
rect 281994 273922 282050 273978
rect 282118 273922 282174 273978
rect 282242 273922 282298 273978
rect 282366 273922 282422 273978
rect 281994 256294 282050 256350
rect 282118 256294 282174 256350
rect 282242 256294 282298 256350
rect 282366 256294 282422 256350
rect 281994 256170 282050 256226
rect 282118 256170 282174 256226
rect 282242 256170 282298 256226
rect 282366 256170 282422 256226
rect 281994 256046 282050 256102
rect 282118 256046 282174 256102
rect 282242 256046 282298 256102
rect 282366 256046 282422 256102
rect 281994 255922 282050 255978
rect 282118 255922 282174 255978
rect 282242 255922 282298 255978
rect 282366 255922 282422 255978
rect 281994 238294 282050 238350
rect 282118 238294 282174 238350
rect 282242 238294 282298 238350
rect 282366 238294 282422 238350
rect 281994 238170 282050 238226
rect 282118 238170 282174 238226
rect 282242 238170 282298 238226
rect 282366 238170 282422 238226
rect 281994 238046 282050 238102
rect 282118 238046 282174 238102
rect 282242 238046 282298 238102
rect 282366 238046 282422 238102
rect 281994 237922 282050 237978
rect 282118 237922 282174 237978
rect 282242 237922 282298 237978
rect 282366 237922 282422 237978
rect 281994 220294 282050 220350
rect 282118 220294 282174 220350
rect 282242 220294 282298 220350
rect 282366 220294 282422 220350
rect 281994 220170 282050 220226
rect 282118 220170 282174 220226
rect 282242 220170 282298 220226
rect 282366 220170 282422 220226
rect 281994 220046 282050 220102
rect 282118 220046 282174 220102
rect 282242 220046 282298 220102
rect 282366 220046 282422 220102
rect 281994 219922 282050 219978
rect 282118 219922 282174 219978
rect 282242 219922 282298 219978
rect 282366 219922 282422 219978
rect 281994 202294 282050 202350
rect 282118 202294 282174 202350
rect 282242 202294 282298 202350
rect 282366 202294 282422 202350
rect 281994 202170 282050 202226
rect 282118 202170 282174 202226
rect 282242 202170 282298 202226
rect 282366 202170 282422 202226
rect 281994 202046 282050 202102
rect 282118 202046 282174 202102
rect 282242 202046 282298 202102
rect 282366 202046 282422 202102
rect 281994 201922 282050 201978
rect 282118 201922 282174 201978
rect 282242 201922 282298 201978
rect 282366 201922 282422 201978
rect 281994 184294 282050 184350
rect 282118 184294 282174 184350
rect 282242 184294 282298 184350
rect 282366 184294 282422 184350
rect 281994 184170 282050 184226
rect 282118 184170 282174 184226
rect 282242 184170 282298 184226
rect 282366 184170 282422 184226
rect 281994 184046 282050 184102
rect 282118 184046 282174 184102
rect 282242 184046 282298 184102
rect 282366 184046 282422 184102
rect 281994 183922 282050 183978
rect 282118 183922 282174 183978
rect 282242 183922 282298 183978
rect 282366 183922 282422 183978
rect 281994 166294 282050 166350
rect 282118 166294 282174 166350
rect 282242 166294 282298 166350
rect 282366 166294 282422 166350
rect 281994 166170 282050 166226
rect 282118 166170 282174 166226
rect 282242 166170 282298 166226
rect 282366 166170 282422 166226
rect 281994 166046 282050 166102
rect 282118 166046 282174 166102
rect 282242 166046 282298 166102
rect 282366 166046 282422 166102
rect 281994 165922 282050 165978
rect 282118 165922 282174 165978
rect 282242 165922 282298 165978
rect 282366 165922 282422 165978
rect 281994 148294 282050 148350
rect 282118 148294 282174 148350
rect 282242 148294 282298 148350
rect 282366 148294 282422 148350
rect 281994 148170 282050 148226
rect 282118 148170 282174 148226
rect 282242 148170 282298 148226
rect 282366 148170 282422 148226
rect 281994 148046 282050 148102
rect 282118 148046 282174 148102
rect 282242 148046 282298 148102
rect 282366 148046 282422 148102
rect 281994 147922 282050 147978
rect 282118 147922 282174 147978
rect 282242 147922 282298 147978
rect 282366 147922 282422 147978
rect 281994 130294 282050 130350
rect 282118 130294 282174 130350
rect 282242 130294 282298 130350
rect 282366 130294 282422 130350
rect 281994 130170 282050 130226
rect 282118 130170 282174 130226
rect 282242 130170 282298 130226
rect 282366 130170 282422 130226
rect 281994 130046 282050 130102
rect 282118 130046 282174 130102
rect 282242 130046 282298 130102
rect 282366 130046 282422 130102
rect 281994 129922 282050 129978
rect 282118 129922 282174 129978
rect 282242 129922 282298 129978
rect 282366 129922 282422 129978
rect 281994 112294 282050 112350
rect 282118 112294 282174 112350
rect 282242 112294 282298 112350
rect 282366 112294 282422 112350
rect 281994 112170 282050 112226
rect 282118 112170 282174 112226
rect 282242 112170 282298 112226
rect 282366 112170 282422 112226
rect 281994 112046 282050 112102
rect 282118 112046 282174 112102
rect 282242 112046 282298 112102
rect 282366 112046 282422 112102
rect 281994 111922 282050 111978
rect 282118 111922 282174 111978
rect 282242 111922 282298 111978
rect 282366 111922 282422 111978
rect 281994 94294 282050 94350
rect 282118 94294 282174 94350
rect 282242 94294 282298 94350
rect 282366 94294 282422 94350
rect 281994 94170 282050 94226
rect 282118 94170 282174 94226
rect 282242 94170 282298 94226
rect 282366 94170 282422 94226
rect 273980 92402 274036 92458
rect 281994 94046 282050 94102
rect 282118 94046 282174 94102
rect 282242 94046 282298 94102
rect 282366 94046 282422 94102
rect 281994 93922 282050 93978
rect 282118 93922 282174 93978
rect 282242 93922 282298 93978
rect 282366 93922 282422 93978
rect 273868 81422 273924 81478
rect 273532 72962 273588 73018
rect 282604 86462 282660 86518
rect 285714 298294 285770 298350
rect 285838 298294 285894 298350
rect 285962 298294 286018 298350
rect 286086 298294 286142 298350
rect 285714 298170 285770 298226
rect 285838 298170 285894 298226
rect 285962 298170 286018 298226
rect 286086 298170 286142 298226
rect 285714 298046 285770 298102
rect 285838 298046 285894 298102
rect 285962 298046 286018 298102
rect 286086 298046 286142 298102
rect 285714 297922 285770 297978
rect 285838 297922 285894 297978
rect 285962 297922 286018 297978
rect 286086 297922 286142 297978
rect 285714 280294 285770 280350
rect 285838 280294 285894 280350
rect 285962 280294 286018 280350
rect 286086 280294 286142 280350
rect 285714 280170 285770 280226
rect 285838 280170 285894 280226
rect 285962 280170 286018 280226
rect 286086 280170 286142 280226
rect 285714 280046 285770 280102
rect 285838 280046 285894 280102
rect 285962 280046 286018 280102
rect 286086 280046 286142 280102
rect 285714 279922 285770 279978
rect 285838 279922 285894 279978
rect 285962 279922 286018 279978
rect 286086 279922 286142 279978
rect 285714 262294 285770 262350
rect 285838 262294 285894 262350
rect 285962 262294 286018 262350
rect 286086 262294 286142 262350
rect 285714 262170 285770 262226
rect 285838 262170 285894 262226
rect 285962 262170 286018 262226
rect 286086 262170 286142 262226
rect 285714 262046 285770 262102
rect 285838 262046 285894 262102
rect 285962 262046 286018 262102
rect 286086 262046 286142 262102
rect 285714 261922 285770 261978
rect 285838 261922 285894 261978
rect 285962 261922 286018 261978
rect 286086 261922 286142 261978
rect 285714 244294 285770 244350
rect 285838 244294 285894 244350
rect 285962 244294 286018 244350
rect 286086 244294 286142 244350
rect 285714 244170 285770 244226
rect 285838 244170 285894 244226
rect 285962 244170 286018 244226
rect 286086 244170 286142 244226
rect 285714 244046 285770 244102
rect 285838 244046 285894 244102
rect 285962 244046 286018 244102
rect 286086 244046 286142 244102
rect 285714 243922 285770 243978
rect 285838 243922 285894 243978
rect 285962 243922 286018 243978
rect 286086 243922 286142 243978
rect 285714 226294 285770 226350
rect 285838 226294 285894 226350
rect 285962 226294 286018 226350
rect 286086 226294 286142 226350
rect 285714 226170 285770 226226
rect 285838 226170 285894 226226
rect 285962 226170 286018 226226
rect 286086 226170 286142 226226
rect 285714 226046 285770 226102
rect 285838 226046 285894 226102
rect 285962 226046 286018 226102
rect 286086 226046 286142 226102
rect 285714 225922 285770 225978
rect 285838 225922 285894 225978
rect 285962 225922 286018 225978
rect 286086 225922 286142 225978
rect 285714 208294 285770 208350
rect 285838 208294 285894 208350
rect 285962 208294 286018 208350
rect 286086 208294 286142 208350
rect 285714 208170 285770 208226
rect 285838 208170 285894 208226
rect 285962 208170 286018 208226
rect 286086 208170 286142 208226
rect 285714 208046 285770 208102
rect 285838 208046 285894 208102
rect 285962 208046 286018 208102
rect 286086 208046 286142 208102
rect 285714 207922 285770 207978
rect 285838 207922 285894 207978
rect 285962 207922 286018 207978
rect 286086 207922 286142 207978
rect 285714 190294 285770 190350
rect 285838 190294 285894 190350
rect 285962 190294 286018 190350
rect 286086 190294 286142 190350
rect 285714 190170 285770 190226
rect 285838 190170 285894 190226
rect 285962 190170 286018 190226
rect 286086 190170 286142 190226
rect 285714 190046 285770 190102
rect 285838 190046 285894 190102
rect 285962 190046 286018 190102
rect 286086 190046 286142 190102
rect 285714 189922 285770 189978
rect 285838 189922 285894 189978
rect 285962 189922 286018 189978
rect 286086 189922 286142 189978
rect 285714 172294 285770 172350
rect 285838 172294 285894 172350
rect 285962 172294 286018 172350
rect 286086 172294 286142 172350
rect 285714 172170 285770 172226
rect 285838 172170 285894 172226
rect 285962 172170 286018 172226
rect 286086 172170 286142 172226
rect 285714 172046 285770 172102
rect 285838 172046 285894 172102
rect 285962 172046 286018 172102
rect 286086 172046 286142 172102
rect 285714 171922 285770 171978
rect 285838 171922 285894 171978
rect 285962 171922 286018 171978
rect 286086 171922 286142 171978
rect 285714 154294 285770 154350
rect 285838 154294 285894 154350
rect 285962 154294 286018 154350
rect 286086 154294 286142 154350
rect 285714 154170 285770 154226
rect 285838 154170 285894 154226
rect 285962 154170 286018 154226
rect 286086 154170 286142 154226
rect 285714 154046 285770 154102
rect 285838 154046 285894 154102
rect 285962 154046 286018 154102
rect 286086 154046 286142 154102
rect 285714 153922 285770 153978
rect 285838 153922 285894 153978
rect 285962 153922 286018 153978
rect 286086 153922 286142 153978
rect 285714 136294 285770 136350
rect 285838 136294 285894 136350
rect 285962 136294 286018 136350
rect 286086 136294 286142 136350
rect 285714 136170 285770 136226
rect 285838 136170 285894 136226
rect 285962 136170 286018 136226
rect 286086 136170 286142 136226
rect 285714 136046 285770 136102
rect 285838 136046 285894 136102
rect 285962 136046 286018 136102
rect 286086 136046 286142 136102
rect 285714 135922 285770 135978
rect 285838 135922 285894 135978
rect 285962 135922 286018 135978
rect 286086 135922 286142 135978
rect 285714 118294 285770 118350
rect 285838 118294 285894 118350
rect 285962 118294 286018 118350
rect 286086 118294 286142 118350
rect 285714 118170 285770 118226
rect 285838 118170 285894 118226
rect 285962 118170 286018 118226
rect 286086 118170 286142 118226
rect 285714 118046 285770 118102
rect 285838 118046 285894 118102
rect 285962 118046 286018 118102
rect 286086 118046 286142 118102
rect 285714 117922 285770 117978
rect 285838 117922 285894 117978
rect 285962 117922 286018 117978
rect 286086 117922 286142 117978
rect 286300 108242 286356 108298
rect 285714 100294 285770 100350
rect 285838 100294 285894 100350
rect 285962 100294 286018 100350
rect 286086 100294 286142 100350
rect 285714 100170 285770 100226
rect 285838 100170 285894 100226
rect 285962 100170 286018 100226
rect 286086 100170 286142 100226
rect 285714 100046 285770 100102
rect 285838 100046 285894 100102
rect 285962 100046 286018 100102
rect 286086 100046 286142 100102
rect 285714 99922 285770 99978
rect 285838 99922 285894 99978
rect 285962 99922 286018 99978
rect 286086 99922 286142 99978
rect 283836 85202 283892 85258
rect 290668 88262 290724 88318
rect 294028 88442 294084 88498
rect 292348 88082 292404 88138
rect 296492 85022 296548 85078
rect 310828 304982 310884 305038
rect 309148 303182 309204 303238
rect 310604 301202 310660 301258
rect 310828 301202 310884 301258
rect 315084 301562 315140 301618
rect 312714 292294 312770 292350
rect 312838 292294 312894 292350
rect 312962 292294 313018 292350
rect 313086 292294 313142 292350
rect 312714 292170 312770 292226
rect 312838 292170 312894 292226
rect 312962 292170 313018 292226
rect 313086 292170 313142 292226
rect 312714 292046 312770 292102
rect 312838 292046 312894 292102
rect 312962 292046 313018 292102
rect 313086 292046 313142 292102
rect 312714 291922 312770 291978
rect 312838 291922 312894 291978
rect 312962 291922 313018 291978
rect 313086 291922 313142 291978
rect 312714 274294 312770 274350
rect 312838 274294 312894 274350
rect 312962 274294 313018 274350
rect 313086 274294 313142 274350
rect 312714 274170 312770 274226
rect 312838 274170 312894 274226
rect 312962 274170 313018 274226
rect 313086 274170 313142 274226
rect 312714 274046 312770 274102
rect 312838 274046 312894 274102
rect 312962 274046 313018 274102
rect 313086 274046 313142 274102
rect 312714 273922 312770 273978
rect 312838 273922 312894 273978
rect 312962 273922 313018 273978
rect 313086 273922 313142 273978
rect 312714 256294 312770 256350
rect 312838 256294 312894 256350
rect 312962 256294 313018 256350
rect 313086 256294 313142 256350
rect 312714 256170 312770 256226
rect 312838 256170 312894 256226
rect 312962 256170 313018 256226
rect 313086 256170 313142 256226
rect 312714 256046 312770 256102
rect 312838 256046 312894 256102
rect 312962 256046 313018 256102
rect 313086 256046 313142 256102
rect 312714 255922 312770 255978
rect 312838 255922 312894 255978
rect 312962 255922 313018 255978
rect 313086 255922 313142 255978
rect 312714 238294 312770 238350
rect 312838 238294 312894 238350
rect 312962 238294 313018 238350
rect 313086 238294 313142 238350
rect 312714 238170 312770 238226
rect 312838 238170 312894 238226
rect 312962 238170 313018 238226
rect 313086 238170 313142 238226
rect 312714 238046 312770 238102
rect 312838 238046 312894 238102
rect 312962 238046 313018 238102
rect 313086 238046 313142 238102
rect 312714 237922 312770 237978
rect 312838 237922 312894 237978
rect 312962 237922 313018 237978
rect 313086 237922 313142 237978
rect 312714 220294 312770 220350
rect 312838 220294 312894 220350
rect 312962 220294 313018 220350
rect 313086 220294 313142 220350
rect 312714 220170 312770 220226
rect 312838 220170 312894 220226
rect 312962 220170 313018 220226
rect 313086 220170 313142 220226
rect 312714 220046 312770 220102
rect 312838 220046 312894 220102
rect 312962 220046 313018 220102
rect 313086 220046 313142 220102
rect 312714 219922 312770 219978
rect 312838 219922 312894 219978
rect 312962 219922 313018 219978
rect 313086 219922 313142 219978
rect 312714 202294 312770 202350
rect 312838 202294 312894 202350
rect 312962 202294 313018 202350
rect 313086 202294 313142 202350
rect 312714 202170 312770 202226
rect 312838 202170 312894 202226
rect 312962 202170 313018 202226
rect 313086 202170 313142 202226
rect 312714 202046 312770 202102
rect 312838 202046 312894 202102
rect 312962 202046 313018 202102
rect 313086 202046 313142 202102
rect 312714 201922 312770 201978
rect 312838 201922 312894 201978
rect 312962 201922 313018 201978
rect 313086 201922 313142 201978
rect 312714 184294 312770 184350
rect 312838 184294 312894 184350
rect 312962 184294 313018 184350
rect 313086 184294 313142 184350
rect 312714 184170 312770 184226
rect 312838 184170 312894 184226
rect 312962 184170 313018 184226
rect 313086 184170 313142 184226
rect 312714 184046 312770 184102
rect 312838 184046 312894 184102
rect 312962 184046 313018 184102
rect 313086 184046 313142 184102
rect 312714 183922 312770 183978
rect 312838 183922 312894 183978
rect 312962 183922 313018 183978
rect 313086 183922 313142 183978
rect 312714 166294 312770 166350
rect 312838 166294 312894 166350
rect 312962 166294 313018 166350
rect 313086 166294 313142 166350
rect 312714 166170 312770 166226
rect 312838 166170 312894 166226
rect 312962 166170 313018 166226
rect 313086 166170 313142 166226
rect 312714 166046 312770 166102
rect 312838 166046 312894 166102
rect 312962 166046 313018 166102
rect 313086 166046 313142 166102
rect 312714 165922 312770 165978
rect 312838 165922 312894 165978
rect 312962 165922 313018 165978
rect 313086 165922 313142 165978
rect 312714 148294 312770 148350
rect 312838 148294 312894 148350
rect 312962 148294 313018 148350
rect 313086 148294 313142 148350
rect 312714 148170 312770 148226
rect 312838 148170 312894 148226
rect 312962 148170 313018 148226
rect 313086 148170 313142 148226
rect 312714 148046 312770 148102
rect 312838 148046 312894 148102
rect 312962 148046 313018 148102
rect 313086 148046 313142 148102
rect 312714 147922 312770 147978
rect 312838 147922 312894 147978
rect 312962 147922 313018 147978
rect 313086 147922 313142 147978
rect 312714 130294 312770 130350
rect 312838 130294 312894 130350
rect 312962 130294 313018 130350
rect 313086 130294 313142 130350
rect 312714 130170 312770 130226
rect 312838 130170 312894 130226
rect 312962 130170 313018 130226
rect 313086 130170 313142 130226
rect 312714 130046 312770 130102
rect 312838 130046 312894 130102
rect 312962 130046 313018 130102
rect 313086 130046 313142 130102
rect 312714 129922 312770 129978
rect 312838 129922 312894 129978
rect 312962 129922 313018 129978
rect 313086 129922 313142 129978
rect 312714 112294 312770 112350
rect 312838 112294 312894 112350
rect 312962 112294 313018 112350
rect 313086 112294 313142 112350
rect 312714 112170 312770 112226
rect 312838 112170 312894 112226
rect 312962 112170 313018 112226
rect 313086 112170 313142 112226
rect 312714 112046 312770 112102
rect 312838 112046 312894 112102
rect 312962 112046 313018 112102
rect 313086 112046 313142 112102
rect 312714 111922 312770 111978
rect 312838 111922 312894 111978
rect 312962 111922 313018 111978
rect 313086 111922 313142 111978
rect 312714 94294 312770 94350
rect 312838 94294 312894 94350
rect 312962 94294 313018 94350
rect 313086 94294 313142 94350
rect 312714 94170 312770 94226
rect 312838 94170 312894 94226
rect 312962 94170 313018 94226
rect 313086 94170 313142 94226
rect 312714 94046 312770 94102
rect 312838 94046 312894 94102
rect 312962 94046 313018 94102
rect 313086 94046 313142 94102
rect 312714 93922 312770 93978
rect 312838 93922 312894 93978
rect 312962 93922 313018 93978
rect 313086 93922 313142 93978
rect 299068 84842 299124 84898
rect 285714 82294 285770 82350
rect 285838 82294 285894 82350
rect 285962 82294 286018 82350
rect 286086 82294 286142 82350
rect 285714 82170 285770 82226
rect 285838 82170 285894 82226
rect 285962 82170 286018 82226
rect 286086 82170 286142 82226
rect 285714 82046 285770 82102
rect 285838 82046 285894 82102
rect 285962 82046 286018 82102
rect 286086 82046 286142 82102
rect 285714 81922 285770 81978
rect 285838 81922 285894 81978
rect 285962 81922 286018 81978
rect 286086 81922 286142 81978
rect 319004 302462 319060 302518
rect 324156 304802 324212 304858
rect 324604 303362 324660 303418
rect 324492 303182 324548 303238
rect 327740 304982 327796 305038
rect 327292 303182 327348 303238
rect 330428 304082 330484 304138
rect 330876 303722 330932 303778
rect 320796 302282 320852 302338
rect 329868 302282 329924 302338
rect 320684 302102 320740 302158
rect 329420 302102 329476 302158
rect 316434 298294 316490 298350
rect 316558 298294 316614 298350
rect 316682 298294 316738 298350
rect 316806 298294 316862 298350
rect 316434 298170 316490 298226
rect 316558 298170 316614 298226
rect 316682 298170 316738 298226
rect 316806 298170 316862 298226
rect 316434 298046 316490 298102
rect 316558 298046 316614 298102
rect 316682 298046 316738 298102
rect 316806 298046 316862 298102
rect 316434 297922 316490 297978
rect 316558 297922 316614 297978
rect 316682 297922 316738 297978
rect 316806 297922 316862 297978
rect 316434 280294 316490 280350
rect 316558 280294 316614 280350
rect 316682 280294 316738 280350
rect 316806 280294 316862 280350
rect 316434 280170 316490 280226
rect 316558 280170 316614 280226
rect 316682 280170 316738 280226
rect 316806 280170 316862 280226
rect 316434 280046 316490 280102
rect 316558 280046 316614 280102
rect 316682 280046 316738 280102
rect 316806 280046 316862 280102
rect 316434 279922 316490 279978
rect 316558 279922 316614 279978
rect 316682 279922 316738 279978
rect 316806 279922 316862 279978
rect 316434 262294 316490 262350
rect 316558 262294 316614 262350
rect 316682 262294 316738 262350
rect 316806 262294 316862 262350
rect 316434 262170 316490 262226
rect 316558 262170 316614 262226
rect 316682 262170 316738 262226
rect 316806 262170 316862 262226
rect 316434 262046 316490 262102
rect 316558 262046 316614 262102
rect 316682 262046 316738 262102
rect 316806 262046 316862 262102
rect 316434 261922 316490 261978
rect 316558 261922 316614 261978
rect 316682 261922 316738 261978
rect 316806 261922 316862 261978
rect 316434 244294 316490 244350
rect 316558 244294 316614 244350
rect 316682 244294 316738 244350
rect 316806 244294 316862 244350
rect 316434 244170 316490 244226
rect 316558 244170 316614 244226
rect 316682 244170 316738 244226
rect 316806 244170 316862 244226
rect 316434 244046 316490 244102
rect 316558 244046 316614 244102
rect 316682 244046 316738 244102
rect 316806 244046 316862 244102
rect 316434 243922 316490 243978
rect 316558 243922 316614 243978
rect 316682 243922 316738 243978
rect 316806 243922 316862 243978
rect 316434 226294 316490 226350
rect 316558 226294 316614 226350
rect 316682 226294 316738 226350
rect 316806 226294 316862 226350
rect 316434 226170 316490 226226
rect 316558 226170 316614 226226
rect 316682 226170 316738 226226
rect 316806 226170 316862 226226
rect 316434 226046 316490 226102
rect 316558 226046 316614 226102
rect 316682 226046 316738 226102
rect 316806 226046 316862 226102
rect 316434 225922 316490 225978
rect 316558 225922 316614 225978
rect 316682 225922 316738 225978
rect 316806 225922 316862 225978
rect 316434 208294 316490 208350
rect 316558 208294 316614 208350
rect 316682 208294 316738 208350
rect 316806 208294 316862 208350
rect 316434 208170 316490 208226
rect 316558 208170 316614 208226
rect 316682 208170 316738 208226
rect 316806 208170 316862 208226
rect 316434 208046 316490 208102
rect 316558 208046 316614 208102
rect 316682 208046 316738 208102
rect 316806 208046 316862 208102
rect 316434 207922 316490 207978
rect 316558 207922 316614 207978
rect 316682 207922 316738 207978
rect 316806 207922 316862 207978
rect 316434 190294 316490 190350
rect 316558 190294 316614 190350
rect 316682 190294 316738 190350
rect 316806 190294 316862 190350
rect 316434 190170 316490 190226
rect 316558 190170 316614 190226
rect 316682 190170 316738 190226
rect 316806 190170 316862 190226
rect 316434 190046 316490 190102
rect 316558 190046 316614 190102
rect 316682 190046 316738 190102
rect 316806 190046 316862 190102
rect 316434 189922 316490 189978
rect 316558 189922 316614 189978
rect 316682 189922 316738 189978
rect 316806 189922 316862 189978
rect 316434 172294 316490 172350
rect 316558 172294 316614 172350
rect 316682 172294 316738 172350
rect 316806 172294 316862 172350
rect 316434 172170 316490 172226
rect 316558 172170 316614 172226
rect 316682 172170 316738 172226
rect 316806 172170 316862 172226
rect 316434 172046 316490 172102
rect 316558 172046 316614 172102
rect 316682 172046 316738 172102
rect 316806 172046 316862 172102
rect 316434 171922 316490 171978
rect 316558 171922 316614 171978
rect 316682 171922 316738 171978
rect 316806 171922 316862 171978
rect 316434 154294 316490 154350
rect 316558 154294 316614 154350
rect 316682 154294 316738 154350
rect 316806 154294 316862 154350
rect 316434 154170 316490 154226
rect 316558 154170 316614 154226
rect 316682 154170 316738 154226
rect 316806 154170 316862 154226
rect 316434 154046 316490 154102
rect 316558 154046 316614 154102
rect 316682 154046 316738 154102
rect 316806 154046 316862 154102
rect 316434 153922 316490 153978
rect 316558 153922 316614 153978
rect 316682 153922 316738 153978
rect 316806 153922 316862 153978
rect 316434 136294 316490 136350
rect 316558 136294 316614 136350
rect 316682 136294 316738 136350
rect 316806 136294 316862 136350
rect 316434 136170 316490 136226
rect 316558 136170 316614 136226
rect 316682 136170 316738 136226
rect 316806 136170 316862 136226
rect 316434 136046 316490 136102
rect 316558 136046 316614 136102
rect 316682 136046 316738 136102
rect 316806 136046 316862 136102
rect 316434 135922 316490 135978
rect 316558 135922 316614 135978
rect 316682 135922 316738 135978
rect 316806 135922 316862 135978
rect 316434 118294 316490 118350
rect 316558 118294 316614 118350
rect 316682 118294 316738 118350
rect 316806 118294 316862 118350
rect 316434 118170 316490 118226
rect 316558 118170 316614 118226
rect 316682 118170 316738 118226
rect 316806 118170 316862 118226
rect 316434 118046 316490 118102
rect 316558 118046 316614 118102
rect 316682 118046 316738 118102
rect 316806 118046 316862 118102
rect 316434 117922 316490 117978
rect 316558 117922 316614 117978
rect 316682 117922 316738 117978
rect 316806 117922 316862 117978
rect 316434 100294 316490 100350
rect 316558 100294 316614 100350
rect 316682 100294 316738 100350
rect 316806 100294 316862 100350
rect 316434 100170 316490 100226
rect 316558 100170 316614 100226
rect 316682 100170 316738 100226
rect 316806 100170 316862 100226
rect 316434 100046 316490 100102
rect 316558 100046 316614 100102
rect 316682 100046 316738 100102
rect 316806 100046 316862 100102
rect 316434 99922 316490 99978
rect 316558 99922 316614 99978
rect 316682 99922 316738 99978
rect 316806 99922 316862 99978
rect 318332 301382 318388 301438
rect 317436 86642 317492 86698
rect 317436 84302 317492 84358
rect 332556 302462 332612 302518
rect 336476 304982 336532 305038
rect 336028 303542 336084 303598
rect 342524 304262 342580 304318
rect 344652 304802 344708 304858
rect 342972 303902 343028 303958
rect 342636 303362 342692 303418
rect 344428 303182 344484 303238
rect 344316 301562 344372 301618
rect 347788 303722 347844 303778
rect 351372 304082 351428 304138
rect 351036 303542 351092 303598
rect 355852 304982 355908 305038
rect 352380 304082 352436 304138
rect 357756 304802 357812 304858
rect 357756 304262 357812 304318
rect 360892 303542 360948 303598
rect 362684 303182 362740 303238
rect 363468 303902 363524 303958
rect 369404 303902 369460 303958
rect 364588 302282 364644 302338
rect 364812 301562 364868 301618
rect 367612 301562 367668 301618
rect 376460 304802 376516 304858
rect 372428 304082 372484 304138
rect 374556 302282 374612 302338
rect 374332 301742 374388 301798
rect 381052 304802 381108 304858
rect 379596 303722 379652 303778
rect 381388 303542 381444 303598
rect 379708 303182 379764 303238
rect 389900 303902 389956 303958
rect 401548 304802 401604 304858
rect 394492 303182 394548 303238
rect 398412 303722 398468 303778
rect 393148 302102 393204 302158
rect 399756 302102 399812 302158
rect 394828 301742 394884 301798
rect 388108 301562 388164 301618
rect 347154 298294 347210 298350
rect 347278 298294 347334 298350
rect 347402 298294 347458 298350
rect 347526 298294 347582 298350
rect 347154 298170 347210 298226
rect 347278 298170 347334 298226
rect 347402 298170 347458 298226
rect 347526 298170 347582 298226
rect 347154 298046 347210 298102
rect 347278 298046 347334 298102
rect 347402 298046 347458 298102
rect 347526 298046 347582 298102
rect 347154 297922 347210 297978
rect 347278 297922 347334 297978
rect 347402 297922 347458 297978
rect 347526 297922 347582 297978
rect 377874 298294 377930 298350
rect 377998 298294 378054 298350
rect 378122 298294 378178 298350
rect 378246 298294 378302 298350
rect 377874 298170 377930 298226
rect 377998 298170 378054 298226
rect 378122 298170 378178 298226
rect 378246 298170 378302 298226
rect 377874 298046 377930 298102
rect 377998 298046 378054 298102
rect 378122 298046 378178 298102
rect 378246 298046 378302 298102
rect 377874 297922 377930 297978
rect 377998 297922 378054 297978
rect 378122 297922 378178 297978
rect 378246 297922 378302 297978
rect 408594 298294 408650 298350
rect 408718 298294 408774 298350
rect 408842 298294 408898 298350
rect 408966 298294 409022 298350
rect 408594 298170 408650 298226
rect 408718 298170 408774 298226
rect 408842 298170 408898 298226
rect 408966 298170 409022 298226
rect 408594 298046 408650 298102
rect 408718 298046 408774 298102
rect 408842 298046 408898 298102
rect 408966 298046 409022 298102
rect 408594 297922 408650 297978
rect 408718 297922 408774 297978
rect 408842 297922 408898 297978
rect 408966 297922 409022 297978
rect 414988 303182 415044 303238
rect 324518 292294 324574 292350
rect 324642 292294 324698 292350
rect 324518 292170 324574 292226
rect 324642 292170 324698 292226
rect 324518 292046 324574 292102
rect 324642 292046 324698 292102
rect 324518 291922 324574 291978
rect 324642 291922 324698 291978
rect 355238 292294 355294 292350
rect 355362 292294 355418 292350
rect 355238 292170 355294 292226
rect 355362 292170 355418 292226
rect 355238 292046 355294 292102
rect 355362 292046 355418 292102
rect 355238 291922 355294 291978
rect 355362 291922 355418 291978
rect 385958 292294 386014 292350
rect 386082 292294 386138 292350
rect 385958 292170 386014 292226
rect 386082 292170 386138 292226
rect 385958 292046 386014 292102
rect 386082 292046 386138 292102
rect 385958 291922 386014 291978
rect 386082 291922 386138 291978
rect 416678 292294 416734 292350
rect 416802 292294 416858 292350
rect 416678 292170 416734 292226
rect 416802 292170 416858 292226
rect 416678 292046 416734 292102
rect 416802 292046 416858 292102
rect 416678 291922 416734 291978
rect 416802 291922 416858 291978
rect 339878 280294 339934 280350
rect 340002 280294 340058 280350
rect 339878 280170 339934 280226
rect 340002 280170 340058 280226
rect 339878 280046 339934 280102
rect 340002 280046 340058 280102
rect 339878 279922 339934 279978
rect 340002 279922 340058 279978
rect 370598 280294 370654 280350
rect 370722 280294 370778 280350
rect 370598 280170 370654 280226
rect 370722 280170 370778 280226
rect 370598 280046 370654 280102
rect 370722 280046 370778 280102
rect 370598 279922 370654 279978
rect 370722 279922 370778 279978
rect 401318 280294 401374 280350
rect 401442 280294 401498 280350
rect 401318 280170 401374 280226
rect 401442 280170 401498 280226
rect 401318 280046 401374 280102
rect 401442 280046 401498 280102
rect 401318 279922 401374 279978
rect 401442 279922 401498 279978
rect 324518 274294 324574 274350
rect 324642 274294 324698 274350
rect 324518 274170 324574 274226
rect 324642 274170 324698 274226
rect 324518 274046 324574 274102
rect 324642 274046 324698 274102
rect 324518 273922 324574 273978
rect 324642 273922 324698 273978
rect 355238 274294 355294 274350
rect 355362 274294 355418 274350
rect 355238 274170 355294 274226
rect 355362 274170 355418 274226
rect 355238 274046 355294 274102
rect 355362 274046 355418 274102
rect 355238 273922 355294 273978
rect 355362 273922 355418 273978
rect 385958 274294 386014 274350
rect 386082 274294 386138 274350
rect 385958 274170 386014 274226
rect 386082 274170 386138 274226
rect 385958 274046 386014 274102
rect 386082 274046 386138 274102
rect 385958 273922 386014 273978
rect 386082 273922 386138 273978
rect 416678 274294 416734 274350
rect 416802 274294 416858 274350
rect 416678 274170 416734 274226
rect 416802 274170 416858 274226
rect 416678 274046 416734 274102
rect 416802 274046 416858 274102
rect 416678 273922 416734 273978
rect 416802 273922 416858 273978
rect 339878 262294 339934 262350
rect 340002 262294 340058 262350
rect 339878 262170 339934 262226
rect 340002 262170 340058 262226
rect 339878 262046 339934 262102
rect 340002 262046 340058 262102
rect 339878 261922 339934 261978
rect 340002 261922 340058 261978
rect 370598 262294 370654 262350
rect 370722 262294 370778 262350
rect 370598 262170 370654 262226
rect 370722 262170 370778 262226
rect 370598 262046 370654 262102
rect 370722 262046 370778 262102
rect 370598 261922 370654 261978
rect 370722 261922 370778 261978
rect 401318 262294 401374 262350
rect 401442 262294 401498 262350
rect 401318 262170 401374 262226
rect 401442 262170 401498 262226
rect 401318 262046 401374 262102
rect 401442 262046 401498 262102
rect 401318 261922 401374 261978
rect 401442 261922 401498 261978
rect 324518 256294 324574 256350
rect 324642 256294 324698 256350
rect 324518 256170 324574 256226
rect 324642 256170 324698 256226
rect 324518 256046 324574 256102
rect 324642 256046 324698 256102
rect 324518 255922 324574 255978
rect 324642 255922 324698 255978
rect 355238 256294 355294 256350
rect 355362 256294 355418 256350
rect 355238 256170 355294 256226
rect 355362 256170 355418 256226
rect 355238 256046 355294 256102
rect 355362 256046 355418 256102
rect 355238 255922 355294 255978
rect 355362 255922 355418 255978
rect 385958 256294 386014 256350
rect 386082 256294 386138 256350
rect 385958 256170 386014 256226
rect 386082 256170 386138 256226
rect 385958 256046 386014 256102
rect 386082 256046 386138 256102
rect 385958 255922 386014 255978
rect 386082 255922 386138 255978
rect 416678 256294 416734 256350
rect 416802 256294 416858 256350
rect 416678 256170 416734 256226
rect 416802 256170 416858 256226
rect 416678 256046 416734 256102
rect 416802 256046 416858 256102
rect 416678 255922 416734 255978
rect 416802 255922 416858 255978
rect 339878 244294 339934 244350
rect 340002 244294 340058 244350
rect 339878 244170 339934 244226
rect 340002 244170 340058 244226
rect 339878 244046 339934 244102
rect 340002 244046 340058 244102
rect 339878 243922 339934 243978
rect 340002 243922 340058 243978
rect 370598 244294 370654 244350
rect 370722 244294 370778 244350
rect 370598 244170 370654 244226
rect 370722 244170 370778 244226
rect 370598 244046 370654 244102
rect 370722 244046 370778 244102
rect 370598 243922 370654 243978
rect 370722 243922 370778 243978
rect 401318 244294 401374 244350
rect 401442 244294 401498 244350
rect 401318 244170 401374 244226
rect 401442 244170 401498 244226
rect 401318 244046 401374 244102
rect 401442 244046 401498 244102
rect 401318 243922 401374 243978
rect 401442 243922 401498 243978
rect 324518 238294 324574 238350
rect 324642 238294 324698 238350
rect 324518 238170 324574 238226
rect 324642 238170 324698 238226
rect 324518 238046 324574 238102
rect 324642 238046 324698 238102
rect 324518 237922 324574 237978
rect 324642 237922 324698 237978
rect 355238 238294 355294 238350
rect 355362 238294 355418 238350
rect 355238 238170 355294 238226
rect 355362 238170 355418 238226
rect 355238 238046 355294 238102
rect 355362 238046 355418 238102
rect 355238 237922 355294 237978
rect 355362 237922 355418 237978
rect 385958 238294 386014 238350
rect 386082 238294 386138 238350
rect 385958 238170 386014 238226
rect 386082 238170 386138 238226
rect 385958 238046 386014 238102
rect 386082 238046 386138 238102
rect 385958 237922 386014 237978
rect 386082 237922 386138 237978
rect 416678 238294 416734 238350
rect 416802 238294 416858 238350
rect 416678 238170 416734 238226
rect 416802 238170 416858 238226
rect 416678 238046 416734 238102
rect 416802 238046 416858 238102
rect 416678 237922 416734 237978
rect 416802 237922 416858 237978
rect 339878 226294 339934 226350
rect 340002 226294 340058 226350
rect 339878 226170 339934 226226
rect 340002 226170 340058 226226
rect 339878 226046 339934 226102
rect 340002 226046 340058 226102
rect 339878 225922 339934 225978
rect 340002 225922 340058 225978
rect 370598 226294 370654 226350
rect 370722 226294 370778 226350
rect 370598 226170 370654 226226
rect 370722 226170 370778 226226
rect 370598 226046 370654 226102
rect 370722 226046 370778 226102
rect 370598 225922 370654 225978
rect 370722 225922 370778 225978
rect 401318 226294 401374 226350
rect 401442 226294 401498 226350
rect 401318 226170 401374 226226
rect 401442 226170 401498 226226
rect 401318 226046 401374 226102
rect 401442 226046 401498 226102
rect 401318 225922 401374 225978
rect 401442 225922 401498 225978
rect 324518 220294 324574 220350
rect 324642 220294 324698 220350
rect 324518 220170 324574 220226
rect 324642 220170 324698 220226
rect 324518 220046 324574 220102
rect 324642 220046 324698 220102
rect 324518 219922 324574 219978
rect 324642 219922 324698 219978
rect 355238 220294 355294 220350
rect 355362 220294 355418 220350
rect 355238 220170 355294 220226
rect 355362 220170 355418 220226
rect 355238 220046 355294 220102
rect 355362 220046 355418 220102
rect 355238 219922 355294 219978
rect 355362 219922 355418 219978
rect 385958 220294 386014 220350
rect 386082 220294 386138 220350
rect 385958 220170 386014 220226
rect 386082 220170 386138 220226
rect 385958 220046 386014 220102
rect 386082 220046 386138 220102
rect 385958 219922 386014 219978
rect 386082 219922 386138 219978
rect 416678 220294 416734 220350
rect 416802 220294 416858 220350
rect 416678 220170 416734 220226
rect 416802 220170 416858 220226
rect 416678 220046 416734 220102
rect 416802 220046 416858 220102
rect 416678 219922 416734 219978
rect 416802 219922 416858 219978
rect 339878 208294 339934 208350
rect 340002 208294 340058 208350
rect 339878 208170 339934 208226
rect 340002 208170 340058 208226
rect 339878 208046 339934 208102
rect 340002 208046 340058 208102
rect 339878 207922 339934 207978
rect 340002 207922 340058 207978
rect 370598 208294 370654 208350
rect 370722 208294 370778 208350
rect 370598 208170 370654 208226
rect 370722 208170 370778 208226
rect 370598 208046 370654 208102
rect 370722 208046 370778 208102
rect 370598 207922 370654 207978
rect 370722 207922 370778 207978
rect 401318 208294 401374 208350
rect 401442 208294 401498 208350
rect 401318 208170 401374 208226
rect 401442 208170 401498 208226
rect 401318 208046 401374 208102
rect 401442 208046 401498 208102
rect 401318 207922 401374 207978
rect 401442 207922 401498 207978
rect 324518 202294 324574 202350
rect 324642 202294 324698 202350
rect 324518 202170 324574 202226
rect 324642 202170 324698 202226
rect 324518 202046 324574 202102
rect 324642 202046 324698 202102
rect 324518 201922 324574 201978
rect 324642 201922 324698 201978
rect 355238 202294 355294 202350
rect 355362 202294 355418 202350
rect 355238 202170 355294 202226
rect 355362 202170 355418 202226
rect 355238 202046 355294 202102
rect 355362 202046 355418 202102
rect 355238 201922 355294 201978
rect 355362 201922 355418 201978
rect 385958 202294 386014 202350
rect 386082 202294 386138 202350
rect 385958 202170 386014 202226
rect 386082 202170 386138 202226
rect 385958 202046 386014 202102
rect 386082 202046 386138 202102
rect 385958 201922 386014 201978
rect 386082 201922 386138 201978
rect 416678 202294 416734 202350
rect 416802 202294 416858 202350
rect 416678 202170 416734 202226
rect 416802 202170 416858 202226
rect 416678 202046 416734 202102
rect 416802 202046 416858 202102
rect 416678 201922 416734 201978
rect 416802 201922 416858 201978
rect 339878 190294 339934 190350
rect 340002 190294 340058 190350
rect 339878 190170 339934 190226
rect 340002 190170 340058 190226
rect 339878 190046 339934 190102
rect 340002 190046 340058 190102
rect 339878 189922 339934 189978
rect 340002 189922 340058 189978
rect 370598 190294 370654 190350
rect 370722 190294 370778 190350
rect 370598 190170 370654 190226
rect 370722 190170 370778 190226
rect 370598 190046 370654 190102
rect 370722 190046 370778 190102
rect 370598 189922 370654 189978
rect 370722 189922 370778 189978
rect 401318 190294 401374 190350
rect 401442 190294 401498 190350
rect 401318 190170 401374 190226
rect 401442 190170 401498 190226
rect 401318 190046 401374 190102
rect 401442 190046 401498 190102
rect 401318 189922 401374 189978
rect 401442 189922 401498 189978
rect 324518 184294 324574 184350
rect 324642 184294 324698 184350
rect 324518 184170 324574 184226
rect 324642 184170 324698 184226
rect 324518 184046 324574 184102
rect 324642 184046 324698 184102
rect 324518 183922 324574 183978
rect 324642 183922 324698 183978
rect 355238 184294 355294 184350
rect 355362 184294 355418 184350
rect 355238 184170 355294 184226
rect 355362 184170 355418 184226
rect 355238 184046 355294 184102
rect 355362 184046 355418 184102
rect 355238 183922 355294 183978
rect 355362 183922 355418 183978
rect 385958 184294 386014 184350
rect 386082 184294 386138 184350
rect 385958 184170 386014 184226
rect 386082 184170 386138 184226
rect 385958 184046 386014 184102
rect 386082 184046 386138 184102
rect 385958 183922 386014 183978
rect 386082 183922 386138 183978
rect 416678 184294 416734 184350
rect 416802 184294 416858 184350
rect 416678 184170 416734 184226
rect 416802 184170 416858 184226
rect 416678 184046 416734 184102
rect 416802 184046 416858 184102
rect 416678 183922 416734 183978
rect 416802 183922 416858 183978
rect 339878 172294 339934 172350
rect 340002 172294 340058 172350
rect 339878 172170 339934 172226
rect 340002 172170 340058 172226
rect 339878 172046 339934 172102
rect 340002 172046 340058 172102
rect 339878 171922 339934 171978
rect 340002 171922 340058 171978
rect 370598 172294 370654 172350
rect 370722 172294 370778 172350
rect 370598 172170 370654 172226
rect 370722 172170 370778 172226
rect 370598 172046 370654 172102
rect 370722 172046 370778 172102
rect 370598 171922 370654 171978
rect 370722 171922 370778 171978
rect 401318 172294 401374 172350
rect 401442 172294 401498 172350
rect 401318 172170 401374 172226
rect 401442 172170 401498 172226
rect 401318 172046 401374 172102
rect 401442 172046 401498 172102
rect 401318 171922 401374 171978
rect 401442 171922 401498 171978
rect 324518 166294 324574 166350
rect 324642 166294 324698 166350
rect 324518 166170 324574 166226
rect 324642 166170 324698 166226
rect 324518 166046 324574 166102
rect 324642 166046 324698 166102
rect 324518 165922 324574 165978
rect 324642 165922 324698 165978
rect 355238 166294 355294 166350
rect 355362 166294 355418 166350
rect 355238 166170 355294 166226
rect 355362 166170 355418 166226
rect 355238 166046 355294 166102
rect 355362 166046 355418 166102
rect 355238 165922 355294 165978
rect 355362 165922 355418 165978
rect 385958 166294 386014 166350
rect 386082 166294 386138 166350
rect 385958 166170 386014 166226
rect 386082 166170 386138 166226
rect 385958 166046 386014 166102
rect 386082 166046 386138 166102
rect 385958 165922 386014 165978
rect 386082 165922 386138 165978
rect 416678 166294 416734 166350
rect 416802 166294 416858 166350
rect 416678 166170 416734 166226
rect 416802 166170 416858 166226
rect 416678 166046 416734 166102
rect 416802 166046 416858 166102
rect 416678 165922 416734 165978
rect 416802 165922 416858 165978
rect 339878 154294 339934 154350
rect 340002 154294 340058 154350
rect 339878 154170 339934 154226
rect 340002 154170 340058 154226
rect 339878 154046 339934 154102
rect 340002 154046 340058 154102
rect 339878 153922 339934 153978
rect 340002 153922 340058 153978
rect 370598 154294 370654 154350
rect 370722 154294 370778 154350
rect 370598 154170 370654 154226
rect 370722 154170 370778 154226
rect 370598 154046 370654 154102
rect 370722 154046 370778 154102
rect 370598 153922 370654 153978
rect 370722 153922 370778 153978
rect 401318 154294 401374 154350
rect 401442 154294 401498 154350
rect 401318 154170 401374 154226
rect 401442 154170 401498 154226
rect 401318 154046 401374 154102
rect 401442 154046 401498 154102
rect 401318 153922 401374 153978
rect 401442 153922 401498 153978
rect 324518 148294 324574 148350
rect 324642 148294 324698 148350
rect 324518 148170 324574 148226
rect 324642 148170 324698 148226
rect 324518 148046 324574 148102
rect 324642 148046 324698 148102
rect 324518 147922 324574 147978
rect 324642 147922 324698 147978
rect 355238 148294 355294 148350
rect 355362 148294 355418 148350
rect 355238 148170 355294 148226
rect 355362 148170 355418 148226
rect 355238 148046 355294 148102
rect 355362 148046 355418 148102
rect 355238 147922 355294 147978
rect 355362 147922 355418 147978
rect 385958 148294 386014 148350
rect 386082 148294 386138 148350
rect 385958 148170 386014 148226
rect 386082 148170 386138 148226
rect 385958 148046 386014 148102
rect 386082 148046 386138 148102
rect 385958 147922 386014 147978
rect 386082 147922 386138 147978
rect 416678 148294 416734 148350
rect 416802 148294 416858 148350
rect 416678 148170 416734 148226
rect 416802 148170 416858 148226
rect 416678 148046 416734 148102
rect 416802 148046 416858 148102
rect 416678 147922 416734 147978
rect 416802 147922 416858 147978
rect 339878 136294 339934 136350
rect 340002 136294 340058 136350
rect 339878 136170 339934 136226
rect 340002 136170 340058 136226
rect 339878 136046 339934 136102
rect 340002 136046 340058 136102
rect 339878 135922 339934 135978
rect 340002 135922 340058 135978
rect 370598 136294 370654 136350
rect 370722 136294 370778 136350
rect 370598 136170 370654 136226
rect 370722 136170 370778 136226
rect 370598 136046 370654 136102
rect 370722 136046 370778 136102
rect 370598 135922 370654 135978
rect 370722 135922 370778 135978
rect 401318 136294 401374 136350
rect 401442 136294 401498 136350
rect 401318 136170 401374 136226
rect 401442 136170 401498 136226
rect 401318 136046 401374 136102
rect 401442 136046 401498 136102
rect 401318 135922 401374 135978
rect 401442 135922 401498 135978
rect 324518 130294 324574 130350
rect 324642 130294 324698 130350
rect 324518 130170 324574 130226
rect 324642 130170 324698 130226
rect 324518 130046 324574 130102
rect 324642 130046 324698 130102
rect 324518 129922 324574 129978
rect 324642 129922 324698 129978
rect 355238 130294 355294 130350
rect 355362 130294 355418 130350
rect 355238 130170 355294 130226
rect 355362 130170 355418 130226
rect 355238 130046 355294 130102
rect 355362 130046 355418 130102
rect 355238 129922 355294 129978
rect 355362 129922 355418 129978
rect 385958 130294 386014 130350
rect 386082 130294 386138 130350
rect 385958 130170 386014 130226
rect 386082 130170 386138 130226
rect 385958 130046 386014 130102
rect 386082 130046 386138 130102
rect 385958 129922 386014 129978
rect 386082 129922 386138 129978
rect 416678 130294 416734 130350
rect 416802 130294 416858 130350
rect 416678 130170 416734 130226
rect 416802 130170 416858 130226
rect 416678 130046 416734 130102
rect 416802 130046 416858 130102
rect 416678 129922 416734 129978
rect 416802 129922 416858 129978
rect 339878 118294 339934 118350
rect 340002 118294 340058 118350
rect 339878 118170 339934 118226
rect 340002 118170 340058 118226
rect 339878 118046 339934 118102
rect 340002 118046 340058 118102
rect 339878 117922 339934 117978
rect 340002 117922 340058 117978
rect 370598 118294 370654 118350
rect 370722 118294 370778 118350
rect 370598 118170 370654 118226
rect 370722 118170 370778 118226
rect 370598 118046 370654 118102
rect 370722 118046 370778 118102
rect 370598 117922 370654 117978
rect 370722 117922 370778 117978
rect 401318 118294 401374 118350
rect 401442 118294 401498 118350
rect 401318 118170 401374 118226
rect 401442 118170 401498 118226
rect 401318 118046 401374 118102
rect 401442 118046 401498 118102
rect 401318 117922 401374 117978
rect 401442 117922 401498 117978
rect 324518 112294 324574 112350
rect 324642 112294 324698 112350
rect 324518 112170 324574 112226
rect 324642 112170 324698 112226
rect 324518 112046 324574 112102
rect 324642 112046 324698 112102
rect 324518 111922 324574 111978
rect 324642 111922 324698 111978
rect 355238 112294 355294 112350
rect 355362 112294 355418 112350
rect 355238 112170 355294 112226
rect 355362 112170 355418 112226
rect 355238 112046 355294 112102
rect 355362 112046 355418 112102
rect 355238 111922 355294 111978
rect 355362 111922 355418 111978
rect 385958 112294 386014 112350
rect 386082 112294 386138 112350
rect 385958 112170 386014 112226
rect 386082 112170 386138 112226
rect 385958 112046 386014 112102
rect 386082 112046 386138 112102
rect 385958 111922 386014 111978
rect 386082 111922 386138 111978
rect 416678 112294 416734 112350
rect 416802 112294 416858 112350
rect 416678 112170 416734 112226
rect 416802 112170 416858 112226
rect 416678 112046 416734 112102
rect 416802 112046 416858 112102
rect 416678 111922 416734 111978
rect 416802 111922 416858 111978
rect 347154 100294 347210 100350
rect 347278 100294 347334 100350
rect 347402 100294 347458 100350
rect 347526 100294 347582 100350
rect 347154 100170 347210 100226
rect 347278 100170 347334 100226
rect 347402 100170 347458 100226
rect 347526 100170 347582 100226
rect 347154 100046 347210 100102
rect 347278 100046 347334 100102
rect 347402 100046 347458 100102
rect 347526 100046 347582 100102
rect 347154 99922 347210 99978
rect 347278 99922 347334 99978
rect 347402 99922 347458 99978
rect 347526 99922 347582 99978
rect 317436 83042 317492 83098
rect 316434 82294 316490 82350
rect 316558 82294 316614 82350
rect 316682 82294 316738 82350
rect 316806 82294 316862 82350
rect 316434 82170 316490 82226
rect 316558 82170 316614 82226
rect 316682 82170 316738 82226
rect 316806 82170 316862 82226
rect 316434 82046 316490 82102
rect 316558 82046 316614 82102
rect 316682 82046 316738 82102
rect 316806 82046 316862 82102
rect 316434 81922 316490 81978
rect 316558 81922 316614 81978
rect 316682 81922 316738 81978
rect 316806 81922 316862 81978
rect 347154 82294 347210 82350
rect 347278 82294 347334 82350
rect 347402 82294 347458 82350
rect 347526 82294 347582 82350
rect 347154 82170 347210 82226
rect 347278 82170 347334 82226
rect 347402 82170 347458 82226
rect 347526 82170 347582 82226
rect 347154 82046 347210 82102
rect 347278 82046 347334 82102
rect 347402 82046 347458 82102
rect 347526 82046 347582 82102
rect 347154 81922 347210 81978
rect 347278 81922 347334 81978
rect 347402 81922 347458 81978
rect 347526 81922 347582 81978
rect 377874 100294 377930 100350
rect 377998 100294 378054 100350
rect 378122 100294 378178 100350
rect 378246 100294 378302 100350
rect 377874 100170 377930 100226
rect 377998 100170 378054 100226
rect 378122 100170 378178 100226
rect 378246 100170 378302 100226
rect 377874 100046 377930 100102
rect 377998 100046 378054 100102
rect 378122 100046 378178 100102
rect 378246 100046 378302 100102
rect 377874 99922 377930 99978
rect 377998 99922 378054 99978
rect 378122 99922 378178 99978
rect 378246 99922 378302 99978
rect 377874 82294 377930 82350
rect 377998 82294 378054 82350
rect 378122 82294 378178 82350
rect 378246 82294 378302 82350
rect 377874 82170 377930 82226
rect 377998 82170 378054 82226
rect 378122 82170 378178 82226
rect 378246 82170 378302 82226
rect 377874 82046 377930 82102
rect 377998 82046 378054 82102
rect 378122 82046 378178 82102
rect 378246 82046 378302 82102
rect 377874 81922 377930 81978
rect 377998 81922 378054 81978
rect 378122 81922 378178 81978
rect 378246 81922 378302 81978
rect 408594 100294 408650 100350
rect 408718 100294 408774 100350
rect 408842 100294 408898 100350
rect 408966 100294 409022 100350
rect 408594 100170 408650 100226
rect 408718 100170 408774 100226
rect 408842 100170 408898 100226
rect 408966 100170 409022 100226
rect 408594 100046 408650 100102
rect 408718 100046 408774 100102
rect 408842 100046 408898 100102
rect 408966 100046 409022 100102
rect 408594 99922 408650 99978
rect 408718 99922 408774 99978
rect 408842 99922 408898 99978
rect 408966 99922 409022 99978
rect 408594 82294 408650 82350
rect 408718 82294 408774 82350
rect 408842 82294 408898 82350
rect 408966 82294 409022 82350
rect 408594 82170 408650 82226
rect 408718 82170 408774 82226
rect 408842 82170 408898 82226
rect 408966 82170 409022 82226
rect 408594 82046 408650 82102
rect 408718 82046 408774 82102
rect 408842 82046 408898 82102
rect 408966 82046 409022 82102
rect 408594 81922 408650 81978
rect 408718 81922 408774 81978
rect 408842 81922 408898 81978
rect 408966 81922 409022 81978
rect 314972 78902 315028 78958
rect 302422 76294 302478 76350
rect 302546 76294 302602 76350
rect 302422 76170 302478 76226
rect 302546 76170 302602 76226
rect 302422 76046 302478 76102
rect 302546 76046 302602 76102
rect 302422 75922 302478 75978
rect 302546 75922 302602 75978
rect 333142 76294 333198 76350
rect 333266 76294 333322 76350
rect 333142 76170 333198 76226
rect 333266 76170 333322 76226
rect 333142 76046 333198 76102
rect 333266 76046 333322 76102
rect 333142 75922 333198 75978
rect 333266 75922 333322 75978
rect 363862 76294 363918 76350
rect 363986 76294 364042 76350
rect 363862 76170 363918 76226
rect 363986 76170 364042 76226
rect 363862 76046 363918 76102
rect 363986 76046 364042 76102
rect 363862 75922 363918 75978
rect 363986 75922 364042 75978
rect 394582 76294 394638 76350
rect 394706 76294 394762 76350
rect 394582 76170 394638 76226
rect 394706 76170 394762 76226
rect 394582 76046 394638 76102
rect 394706 76046 394762 76102
rect 394582 75922 394638 75978
rect 394706 75922 394762 75978
rect 274092 74042 274148 74098
rect 273644 69722 273700 69778
rect 287062 64294 287118 64350
rect 287186 64294 287242 64350
rect 287062 64170 287118 64226
rect 287186 64170 287242 64226
rect 287062 64046 287118 64102
rect 287186 64046 287242 64102
rect 287062 63922 287118 63978
rect 287186 63922 287242 63978
rect 317782 64294 317838 64350
rect 317906 64294 317962 64350
rect 317782 64170 317838 64226
rect 317906 64170 317962 64226
rect 317782 64046 317838 64102
rect 317906 64046 317962 64102
rect 317782 63922 317838 63978
rect 317906 63922 317962 63978
rect 348502 64294 348558 64350
rect 348626 64294 348682 64350
rect 348502 64170 348558 64226
rect 348626 64170 348682 64226
rect 348502 64046 348558 64102
rect 348626 64046 348682 64102
rect 348502 63922 348558 63978
rect 348626 63922 348682 63978
rect 379222 64294 379278 64350
rect 379346 64294 379402 64350
rect 379222 64170 379278 64226
rect 379346 64170 379402 64226
rect 379222 64046 379278 64102
rect 379346 64046 379402 64102
rect 379222 63922 379278 63978
rect 379346 63922 379402 63978
rect 409942 64294 409998 64350
rect 410066 64294 410122 64350
rect 409942 64170 409998 64226
rect 410066 64170 410122 64226
rect 409942 64046 409998 64102
rect 410066 64046 410122 64102
rect 409942 63922 409998 63978
rect 410066 63922 410122 63978
rect 302422 58294 302478 58350
rect 302546 58294 302602 58350
rect 302422 58170 302478 58226
rect 302546 58170 302602 58226
rect 302422 58046 302478 58102
rect 302546 58046 302602 58102
rect 302422 57922 302478 57978
rect 302546 57922 302602 57978
rect 333142 58294 333198 58350
rect 333266 58294 333322 58350
rect 333142 58170 333198 58226
rect 333266 58170 333322 58226
rect 333142 58046 333198 58102
rect 333266 58046 333322 58102
rect 333142 57922 333198 57978
rect 333266 57922 333322 57978
rect 363862 58294 363918 58350
rect 363986 58294 364042 58350
rect 363862 58170 363918 58226
rect 363986 58170 364042 58226
rect 363862 58046 363918 58102
rect 363986 58046 364042 58102
rect 363862 57922 363918 57978
rect 363986 57922 364042 57978
rect 394582 58294 394638 58350
rect 394706 58294 394762 58350
rect 394582 58170 394638 58226
rect 394706 58170 394762 58226
rect 394582 58046 394638 58102
rect 394706 58046 394762 58102
rect 394582 57922 394638 57978
rect 394706 57922 394762 57978
rect 287062 46294 287118 46350
rect 287186 46294 287242 46350
rect 287062 46170 287118 46226
rect 287186 46170 287242 46226
rect 287062 46046 287118 46102
rect 287186 46046 287242 46102
rect 287062 45922 287118 45978
rect 287186 45922 287242 45978
rect 317782 46294 317838 46350
rect 317906 46294 317962 46350
rect 317782 46170 317838 46226
rect 317906 46170 317962 46226
rect 317782 46046 317838 46102
rect 317906 46046 317962 46102
rect 317782 45922 317838 45978
rect 317906 45922 317962 45978
rect 348502 46294 348558 46350
rect 348626 46294 348682 46350
rect 348502 46170 348558 46226
rect 348626 46170 348682 46226
rect 348502 46046 348558 46102
rect 348626 46046 348682 46102
rect 348502 45922 348558 45978
rect 348626 45922 348682 45978
rect 379222 46294 379278 46350
rect 379346 46294 379402 46350
rect 379222 46170 379278 46226
rect 379346 46170 379402 46226
rect 379222 46046 379278 46102
rect 379346 46046 379402 46102
rect 379222 45922 379278 45978
rect 379346 45922 379402 45978
rect 409942 46294 409998 46350
rect 410066 46294 410122 46350
rect 409942 46170 409998 46226
rect 410066 46170 410122 46226
rect 409942 46046 409998 46102
rect 410066 46046 410122 46102
rect 409942 45922 409998 45978
rect 410066 45922 410122 45978
rect 302422 40294 302478 40350
rect 302546 40294 302602 40350
rect 302422 40170 302478 40226
rect 302546 40170 302602 40226
rect 302422 40046 302478 40102
rect 302546 40046 302602 40102
rect 302422 39922 302478 39978
rect 302546 39922 302602 39978
rect 333142 40294 333198 40350
rect 333266 40294 333322 40350
rect 333142 40170 333198 40226
rect 333266 40170 333322 40226
rect 333142 40046 333198 40102
rect 333266 40046 333322 40102
rect 333142 39922 333198 39978
rect 333266 39922 333322 39978
rect 363862 40294 363918 40350
rect 363986 40294 364042 40350
rect 363862 40170 363918 40226
rect 363986 40170 364042 40226
rect 363862 40046 363918 40102
rect 363986 40046 364042 40102
rect 363862 39922 363918 39978
rect 363986 39922 364042 39978
rect 394582 40294 394638 40350
rect 394706 40294 394762 40350
rect 394582 40170 394638 40226
rect 394706 40170 394762 40226
rect 394582 40046 394638 40102
rect 394706 40046 394762 40102
rect 394582 39922 394638 39978
rect 394706 39922 394762 39978
rect 287062 28294 287118 28350
rect 287186 28294 287242 28350
rect 287062 28170 287118 28226
rect 287186 28170 287242 28226
rect 287062 28046 287118 28102
rect 287186 28046 287242 28102
rect 287062 27922 287118 27978
rect 287186 27922 287242 27978
rect 317782 28294 317838 28350
rect 317906 28294 317962 28350
rect 317782 28170 317838 28226
rect 317906 28170 317962 28226
rect 317782 28046 317838 28102
rect 317906 28046 317962 28102
rect 317782 27922 317838 27978
rect 317906 27922 317962 27978
rect 348502 28294 348558 28350
rect 348626 28294 348682 28350
rect 348502 28170 348558 28226
rect 348626 28170 348682 28226
rect 348502 28046 348558 28102
rect 348626 28046 348682 28102
rect 348502 27922 348558 27978
rect 348626 27922 348682 27978
rect 379222 28294 379278 28350
rect 379346 28294 379402 28350
rect 379222 28170 379278 28226
rect 379346 28170 379402 28226
rect 379222 28046 379278 28102
rect 379346 28046 379402 28102
rect 379222 27922 379278 27978
rect 379346 27922 379402 27978
rect 409942 28294 409998 28350
rect 410066 28294 410122 28350
rect 409942 28170 409998 28226
rect 410066 28170 410122 28226
rect 409942 28046 409998 28102
rect 410066 28046 410122 28102
rect 409942 27922 409998 27978
rect 410066 27922 410122 27978
rect 302422 22294 302478 22350
rect 302546 22294 302602 22350
rect 302422 22170 302478 22226
rect 302546 22170 302602 22226
rect 302422 22046 302478 22102
rect 302546 22046 302602 22102
rect 302422 21922 302478 21978
rect 302546 21922 302602 21978
rect 333142 22294 333198 22350
rect 333266 22294 333322 22350
rect 333142 22170 333198 22226
rect 333266 22170 333322 22226
rect 333142 22046 333198 22102
rect 333266 22046 333322 22102
rect 333142 21922 333198 21978
rect 333266 21922 333322 21978
rect 363862 22294 363918 22350
rect 363986 22294 364042 22350
rect 363862 22170 363918 22226
rect 363986 22170 364042 22226
rect 363862 22046 363918 22102
rect 363986 22046 364042 22102
rect 363862 21922 363918 21978
rect 363986 21922 364042 21978
rect 394582 22294 394638 22350
rect 394706 22294 394762 22350
rect 394582 22170 394638 22226
rect 394706 22170 394762 22226
rect 394582 22046 394638 22102
rect 394706 22046 394762 22102
rect 394582 21922 394638 21978
rect 394706 21922 394762 21978
rect 273420 20042 273476 20098
rect 273196 19682 273252 19738
rect 272972 19322 273028 19378
rect 273308 16982 273364 17038
rect 272860 16802 272916 16858
rect 272188 16082 272244 16138
rect 272076 15182 272132 15238
rect 270396 2762 270452 2818
rect 273196 16262 273252 16318
rect 272972 13742 273028 13798
rect 273084 12482 273140 12538
rect 274092 13562 274148 13618
rect 273420 11762 273476 11818
rect 273868 11582 273924 11638
rect 288988 9602 289044 9658
rect 273420 2942 273476 2998
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 277228 2402 277284 2458
rect 271292 422 271348 478
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 304108 2582 304164 2638
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 394044 6542 394100 6598
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 420812 67922 420868 67978
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 423500 301022 423556 301078
rect 424172 101942 424228 101998
rect 424172 13382 424228 13438
rect 425302 76294 425358 76350
rect 425426 76294 425482 76350
rect 425302 76170 425358 76226
rect 425426 76170 425482 76226
rect 425302 76046 425358 76102
rect 425426 76046 425482 76102
rect 425302 75922 425358 75978
rect 425426 75922 425482 75978
rect 425302 58294 425358 58350
rect 425426 58294 425482 58350
rect 425302 58170 425358 58226
rect 425426 58170 425482 58226
rect 425302 58046 425358 58102
rect 425426 58046 425482 58102
rect 425302 57922 425358 57978
rect 425426 57922 425482 57978
rect 425302 40294 425358 40350
rect 425426 40294 425482 40350
rect 425302 40170 425358 40226
rect 425426 40170 425482 40226
rect 425302 40046 425358 40102
rect 425426 40046 425482 40102
rect 425302 39922 425358 39978
rect 425426 39922 425482 39978
rect 425302 22294 425358 22350
rect 425426 22294 425482 22350
rect 425302 22170 425358 22226
rect 425426 22170 425482 22226
rect 425302 22046 425358 22102
rect 425426 22046 425482 22102
rect 425302 21922 425358 21978
rect 425426 21922 425482 21978
rect 425852 79802 425908 79858
rect 427532 79982 427588 80038
rect 428092 75482 428148 75538
rect 428204 13382 428260 13438
rect 428652 75482 428708 75538
rect 431788 299942 431844 299998
rect 431228 89342 431284 89398
rect 432460 90962 432516 91018
rect 432684 98522 432740 98578
rect 432572 89882 432628 89938
rect 433132 91142 433188 91198
rect 433020 89162 433076 89218
rect 432908 85922 432964 85978
rect 432684 20042 432740 20098
rect 433356 90782 433412 90838
rect 435594 382294 435650 382350
rect 435718 382294 435774 382350
rect 435842 382294 435898 382350
rect 435966 382294 436022 382350
rect 435594 382170 435650 382226
rect 435718 382170 435774 382226
rect 435842 382170 435898 382226
rect 435966 382170 436022 382226
rect 435594 382046 435650 382102
rect 435718 382046 435774 382102
rect 435842 382046 435898 382102
rect 435966 382046 436022 382102
rect 435594 381922 435650 381978
rect 435718 381922 435774 381978
rect 435842 381922 435898 381978
rect 435966 381922 436022 381978
rect 434252 80162 434308 80218
rect 434364 301202 434420 301258
rect 435594 364294 435650 364350
rect 435718 364294 435774 364350
rect 435842 364294 435898 364350
rect 435966 364294 436022 364350
rect 435594 364170 435650 364226
rect 435718 364170 435774 364226
rect 435842 364170 435898 364226
rect 435966 364170 436022 364226
rect 435594 364046 435650 364102
rect 435718 364046 435774 364102
rect 435842 364046 435898 364102
rect 435966 364046 436022 364102
rect 435594 363922 435650 363978
rect 435718 363922 435774 363978
rect 435842 363922 435898 363978
rect 435966 363922 436022 363978
rect 435594 346294 435650 346350
rect 435718 346294 435774 346350
rect 435842 346294 435898 346350
rect 435966 346294 436022 346350
rect 435594 346170 435650 346226
rect 435718 346170 435774 346226
rect 435842 346170 435898 346226
rect 435966 346170 436022 346226
rect 435594 346046 435650 346102
rect 435718 346046 435774 346102
rect 435842 346046 435898 346102
rect 435966 346046 436022 346102
rect 435594 345922 435650 345978
rect 435718 345922 435774 345978
rect 435842 345922 435898 345978
rect 435966 345922 436022 345978
rect 435594 328294 435650 328350
rect 435718 328294 435774 328350
rect 435842 328294 435898 328350
rect 435966 328294 436022 328350
rect 435594 328170 435650 328226
rect 435718 328170 435774 328226
rect 435842 328170 435898 328226
rect 435966 328170 436022 328226
rect 435594 328046 435650 328102
rect 435718 328046 435774 328102
rect 435842 328046 435898 328102
rect 435966 328046 436022 328102
rect 435594 327922 435650 327978
rect 435718 327922 435774 327978
rect 435842 327922 435898 327978
rect 435966 327922 436022 327978
rect 435594 310294 435650 310350
rect 435718 310294 435774 310350
rect 435842 310294 435898 310350
rect 435966 310294 436022 310350
rect 435594 310170 435650 310226
rect 435718 310170 435774 310226
rect 435842 310170 435898 310226
rect 435966 310170 436022 310226
rect 435594 310046 435650 310102
rect 435718 310046 435774 310102
rect 435842 310046 435898 310102
rect 435966 310046 436022 310102
rect 435594 309922 435650 309978
rect 435718 309922 435774 309978
rect 435842 309922 435898 309978
rect 435966 309922 436022 309978
rect 435594 292294 435650 292350
rect 435718 292294 435774 292350
rect 435842 292294 435898 292350
rect 435966 292294 436022 292350
rect 435594 292170 435650 292226
rect 435718 292170 435774 292226
rect 435842 292170 435898 292226
rect 435966 292170 436022 292226
rect 435594 292046 435650 292102
rect 435718 292046 435774 292102
rect 435842 292046 435898 292102
rect 435966 292046 436022 292102
rect 435594 291922 435650 291978
rect 435718 291922 435774 291978
rect 435842 291922 435898 291978
rect 435966 291922 436022 291978
rect 435594 274294 435650 274350
rect 435718 274294 435774 274350
rect 435842 274294 435898 274350
rect 435966 274294 436022 274350
rect 435594 274170 435650 274226
rect 435718 274170 435774 274226
rect 435842 274170 435898 274226
rect 435966 274170 436022 274226
rect 435594 274046 435650 274102
rect 435718 274046 435774 274102
rect 435842 274046 435898 274102
rect 435966 274046 436022 274102
rect 435594 273922 435650 273978
rect 435718 273922 435774 273978
rect 435842 273922 435898 273978
rect 435966 273922 436022 273978
rect 435594 256294 435650 256350
rect 435718 256294 435774 256350
rect 435842 256294 435898 256350
rect 435966 256294 436022 256350
rect 435594 256170 435650 256226
rect 435718 256170 435774 256226
rect 435842 256170 435898 256226
rect 435966 256170 436022 256226
rect 435594 256046 435650 256102
rect 435718 256046 435774 256102
rect 435842 256046 435898 256102
rect 435966 256046 436022 256102
rect 435594 255922 435650 255978
rect 435718 255922 435774 255978
rect 435842 255922 435898 255978
rect 435966 255922 436022 255978
rect 435594 238294 435650 238350
rect 435718 238294 435774 238350
rect 435842 238294 435898 238350
rect 435966 238294 436022 238350
rect 435594 238170 435650 238226
rect 435718 238170 435774 238226
rect 435842 238170 435898 238226
rect 435966 238170 436022 238226
rect 435594 238046 435650 238102
rect 435718 238046 435774 238102
rect 435842 238046 435898 238102
rect 435966 238046 436022 238102
rect 435594 237922 435650 237978
rect 435718 237922 435774 237978
rect 435842 237922 435898 237978
rect 435966 237922 436022 237978
rect 435594 220294 435650 220350
rect 435718 220294 435774 220350
rect 435842 220294 435898 220350
rect 435966 220294 436022 220350
rect 435594 220170 435650 220226
rect 435718 220170 435774 220226
rect 435842 220170 435898 220226
rect 435966 220170 436022 220226
rect 435594 220046 435650 220102
rect 435718 220046 435774 220102
rect 435842 220046 435898 220102
rect 435966 220046 436022 220102
rect 435594 219922 435650 219978
rect 435718 219922 435774 219978
rect 435842 219922 435898 219978
rect 435966 219922 436022 219978
rect 435594 202294 435650 202350
rect 435718 202294 435774 202350
rect 435842 202294 435898 202350
rect 435966 202294 436022 202350
rect 435594 202170 435650 202226
rect 435718 202170 435774 202226
rect 435842 202170 435898 202226
rect 435966 202170 436022 202226
rect 435594 202046 435650 202102
rect 435718 202046 435774 202102
rect 435842 202046 435898 202102
rect 435966 202046 436022 202102
rect 435594 201922 435650 201978
rect 435718 201922 435774 201978
rect 435842 201922 435898 201978
rect 435966 201922 436022 201978
rect 435594 184294 435650 184350
rect 435718 184294 435774 184350
rect 435842 184294 435898 184350
rect 435966 184294 436022 184350
rect 435594 184170 435650 184226
rect 435718 184170 435774 184226
rect 435842 184170 435898 184226
rect 435966 184170 436022 184226
rect 435594 184046 435650 184102
rect 435718 184046 435774 184102
rect 435842 184046 435898 184102
rect 435966 184046 436022 184102
rect 435594 183922 435650 183978
rect 435718 183922 435774 183978
rect 435842 183922 435898 183978
rect 435966 183922 436022 183978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 434476 80342 434532 80398
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 436268 93122 436324 93178
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 436268 82862 436324 82918
rect 436828 299762 436884 299818
rect 436492 87542 436548 87598
rect 436604 84302 436660 84358
rect 436604 15902 436660 15958
rect 436716 77642 436772 77698
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 439314 388294 439370 388350
rect 439438 388294 439494 388350
rect 439562 388294 439618 388350
rect 439686 388294 439742 388350
rect 439314 388170 439370 388226
rect 439438 388170 439494 388226
rect 439562 388170 439618 388226
rect 439686 388170 439742 388226
rect 439314 388046 439370 388102
rect 439438 388046 439494 388102
rect 439562 388046 439618 388102
rect 439686 388046 439742 388102
rect 439314 387922 439370 387978
rect 439438 387922 439494 387978
rect 439562 387922 439618 387978
rect 439686 387922 439742 387978
rect 437724 96722 437780 96778
rect 437836 300842 437892 300898
rect 437612 94922 437668 94978
rect 439314 370294 439370 370350
rect 439438 370294 439494 370350
rect 439562 370294 439618 370350
rect 439686 370294 439742 370350
rect 439314 370170 439370 370226
rect 439438 370170 439494 370226
rect 439562 370170 439618 370226
rect 439686 370170 439742 370226
rect 439314 370046 439370 370102
rect 439438 370046 439494 370102
rect 439562 370046 439618 370102
rect 439686 370046 439742 370102
rect 439314 369922 439370 369978
rect 439438 369922 439494 369978
rect 439562 369922 439618 369978
rect 439686 369922 439742 369978
rect 437948 91502 438004 91558
rect 439314 352294 439370 352350
rect 439438 352294 439494 352350
rect 439562 352294 439618 352350
rect 439686 352294 439742 352350
rect 439314 352170 439370 352226
rect 439438 352170 439494 352226
rect 439562 352170 439618 352226
rect 439686 352170 439742 352226
rect 439314 352046 439370 352102
rect 439438 352046 439494 352102
rect 439562 352046 439618 352102
rect 439686 352046 439742 352102
rect 439314 351922 439370 351978
rect 439438 351922 439494 351978
rect 439562 351922 439618 351978
rect 439686 351922 439742 351978
rect 439314 334294 439370 334350
rect 439438 334294 439494 334350
rect 439562 334294 439618 334350
rect 439686 334294 439742 334350
rect 439314 334170 439370 334226
rect 439438 334170 439494 334226
rect 439562 334170 439618 334226
rect 439686 334170 439742 334226
rect 439314 334046 439370 334102
rect 439438 334046 439494 334102
rect 439562 334046 439618 334102
rect 439686 334046 439742 334102
rect 439314 333922 439370 333978
rect 439438 333922 439494 333978
rect 439562 333922 439618 333978
rect 439686 333922 439742 333978
rect 439314 316294 439370 316350
rect 439438 316294 439494 316350
rect 439562 316294 439618 316350
rect 439686 316294 439742 316350
rect 439314 316170 439370 316226
rect 439438 316170 439494 316226
rect 439562 316170 439618 316226
rect 439686 316170 439742 316226
rect 439314 316046 439370 316102
rect 439438 316046 439494 316102
rect 439562 316046 439618 316102
rect 439686 316046 439742 316102
rect 439314 315922 439370 315978
rect 439438 315922 439494 315978
rect 439562 315922 439618 315978
rect 439686 315922 439742 315978
rect 439314 298294 439370 298350
rect 439438 298294 439494 298350
rect 439562 298294 439618 298350
rect 439686 298294 439742 298350
rect 439314 298170 439370 298226
rect 439438 298170 439494 298226
rect 439562 298170 439618 298226
rect 439686 298170 439742 298226
rect 439314 298046 439370 298102
rect 439438 298046 439494 298102
rect 439562 298046 439618 298102
rect 439686 298046 439742 298102
rect 439314 297922 439370 297978
rect 439438 297922 439494 297978
rect 439562 297922 439618 297978
rect 439686 297922 439742 297978
rect 439314 280294 439370 280350
rect 439438 280294 439494 280350
rect 439562 280294 439618 280350
rect 439686 280294 439742 280350
rect 439314 280170 439370 280226
rect 439438 280170 439494 280226
rect 439562 280170 439618 280226
rect 439686 280170 439742 280226
rect 439314 280046 439370 280102
rect 439438 280046 439494 280102
rect 439562 280046 439618 280102
rect 439686 280046 439742 280102
rect 439314 279922 439370 279978
rect 439438 279922 439494 279978
rect 439562 279922 439618 279978
rect 439686 279922 439742 279978
rect 439314 262294 439370 262350
rect 439438 262294 439494 262350
rect 439562 262294 439618 262350
rect 439686 262294 439742 262350
rect 439314 262170 439370 262226
rect 439438 262170 439494 262226
rect 439562 262170 439618 262226
rect 439686 262170 439742 262226
rect 439314 262046 439370 262102
rect 439438 262046 439494 262102
rect 439562 262046 439618 262102
rect 439686 262046 439742 262102
rect 439314 261922 439370 261978
rect 439438 261922 439494 261978
rect 439562 261922 439618 261978
rect 439686 261922 439742 261978
rect 439314 244294 439370 244350
rect 439438 244294 439494 244350
rect 439562 244294 439618 244350
rect 439686 244294 439742 244350
rect 439314 244170 439370 244226
rect 439438 244170 439494 244226
rect 439562 244170 439618 244226
rect 439686 244170 439742 244226
rect 439314 244046 439370 244102
rect 439438 244046 439494 244102
rect 439562 244046 439618 244102
rect 439686 244046 439742 244102
rect 439314 243922 439370 243978
rect 439438 243922 439494 243978
rect 439562 243922 439618 243978
rect 439686 243922 439742 243978
rect 439314 226294 439370 226350
rect 439438 226294 439494 226350
rect 439562 226294 439618 226350
rect 439686 226294 439742 226350
rect 439314 226170 439370 226226
rect 439438 226170 439494 226226
rect 439562 226170 439618 226226
rect 439686 226170 439742 226226
rect 439314 226046 439370 226102
rect 439438 226046 439494 226102
rect 439562 226046 439618 226102
rect 439686 226046 439742 226102
rect 439314 225922 439370 225978
rect 439438 225922 439494 225978
rect 439562 225922 439618 225978
rect 439686 225922 439742 225978
rect 439314 208294 439370 208350
rect 439438 208294 439494 208350
rect 439562 208294 439618 208350
rect 439686 208294 439742 208350
rect 439314 208170 439370 208226
rect 439438 208170 439494 208226
rect 439562 208170 439618 208226
rect 439686 208170 439742 208226
rect 439314 208046 439370 208102
rect 439438 208046 439494 208102
rect 439562 208046 439618 208102
rect 439686 208046 439742 208102
rect 439314 207922 439370 207978
rect 439438 207922 439494 207978
rect 439562 207922 439618 207978
rect 439686 207922 439742 207978
rect 439314 190294 439370 190350
rect 439438 190294 439494 190350
rect 439562 190294 439618 190350
rect 439686 190294 439742 190350
rect 439314 190170 439370 190226
rect 439438 190170 439494 190226
rect 439562 190170 439618 190226
rect 439686 190170 439742 190226
rect 439314 190046 439370 190102
rect 439438 190046 439494 190102
rect 439562 190046 439618 190102
rect 439686 190046 439742 190102
rect 439314 189922 439370 189978
rect 439438 189922 439494 189978
rect 439562 189922 439618 189978
rect 439686 189922 439742 189978
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439068 82682 439124 82738
rect 438844 80882 438900 80938
rect 438620 78002 438676 78058
rect 439964 392282 440020 392338
rect 440076 98342 440132 98398
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 440076 87362 440132 87418
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439964 77282 440020 77338
rect 442652 80522 442708 80578
rect 442764 300122 442820 300178
rect 442652 67922 442708 67978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 443100 392462 443156 392518
rect 442876 96542 442932 96598
rect 442876 84122 442932 84178
rect 443212 101762 443268 101818
rect 548044 392462 548100 392518
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 558474 472294 558530 472350
rect 558598 472294 558654 472350
rect 558722 472294 558778 472350
rect 558846 472294 558902 472350
rect 558474 472170 558530 472226
rect 558598 472170 558654 472226
rect 558722 472170 558778 472226
rect 558846 472170 558902 472226
rect 558474 472046 558530 472102
rect 558598 472046 558654 472102
rect 558722 472046 558778 472102
rect 558846 472046 558902 472102
rect 558474 471922 558530 471978
rect 558598 471922 558654 471978
rect 558722 471922 558778 471978
rect 558846 471922 558902 471978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 558474 382294 558530 382350
rect 558598 382294 558654 382350
rect 558722 382294 558778 382350
rect 558846 382294 558902 382350
rect 558474 382170 558530 382226
rect 558598 382170 558654 382226
rect 558722 382170 558778 382226
rect 558846 382170 558902 382226
rect 558474 382046 558530 382102
rect 558598 382046 558654 382102
rect 558722 382046 558778 382102
rect 558846 382046 558902 382102
rect 558474 381922 558530 381978
rect 558598 381922 558654 381978
rect 558722 381922 558778 381978
rect 558846 381922 558902 381978
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 590828 392282 590884 392338
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 463878 370294 463934 370350
rect 464002 370294 464058 370350
rect 463878 370170 463934 370226
rect 464002 370170 464058 370226
rect 463878 370046 463934 370102
rect 464002 370046 464058 370102
rect 463878 369922 463934 369978
rect 464002 369922 464058 369978
rect 494598 370294 494654 370350
rect 494722 370294 494778 370350
rect 494598 370170 494654 370226
rect 494722 370170 494778 370226
rect 494598 370046 494654 370102
rect 494722 370046 494778 370102
rect 494598 369922 494654 369978
rect 494722 369922 494778 369978
rect 525318 370294 525374 370350
rect 525442 370294 525498 370350
rect 525318 370170 525374 370226
rect 525442 370170 525498 370226
rect 525318 370046 525374 370102
rect 525442 370046 525498 370102
rect 525318 369922 525374 369978
rect 525442 369922 525498 369978
rect 556038 370294 556094 370350
rect 556162 370294 556218 370350
rect 556038 370170 556094 370226
rect 556162 370170 556218 370226
rect 556038 370046 556094 370102
rect 556162 370046 556218 370102
rect 556038 369922 556094 369978
rect 556162 369922 556218 369978
rect 448518 364294 448574 364350
rect 448642 364294 448698 364350
rect 448518 364170 448574 364226
rect 448642 364170 448698 364226
rect 448518 364046 448574 364102
rect 448642 364046 448698 364102
rect 448518 363922 448574 363978
rect 448642 363922 448698 363978
rect 479238 364294 479294 364350
rect 479362 364294 479418 364350
rect 479238 364170 479294 364226
rect 479362 364170 479418 364226
rect 479238 364046 479294 364102
rect 479362 364046 479418 364102
rect 479238 363922 479294 363978
rect 479362 363922 479418 363978
rect 509958 364294 510014 364350
rect 510082 364294 510138 364350
rect 509958 364170 510014 364226
rect 510082 364170 510138 364226
rect 509958 364046 510014 364102
rect 510082 364046 510138 364102
rect 509958 363922 510014 363978
rect 510082 363922 510138 363978
rect 540678 364294 540734 364350
rect 540802 364294 540858 364350
rect 540678 364170 540734 364226
rect 540802 364170 540858 364226
rect 540678 364046 540734 364102
rect 540802 364046 540858 364102
rect 540678 363922 540734 363978
rect 540802 363922 540858 363978
rect 571398 364294 571454 364350
rect 571522 364294 571578 364350
rect 571398 364170 571454 364226
rect 571522 364170 571578 364226
rect 571398 364046 571454 364102
rect 571522 364046 571578 364102
rect 571398 363922 571454 363978
rect 571522 363922 571578 363978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 463878 352294 463934 352350
rect 464002 352294 464058 352350
rect 463878 352170 463934 352226
rect 464002 352170 464058 352226
rect 463878 352046 463934 352102
rect 464002 352046 464058 352102
rect 463878 351922 463934 351978
rect 464002 351922 464058 351978
rect 494598 352294 494654 352350
rect 494722 352294 494778 352350
rect 494598 352170 494654 352226
rect 494722 352170 494778 352226
rect 494598 352046 494654 352102
rect 494722 352046 494778 352102
rect 494598 351922 494654 351978
rect 494722 351922 494778 351978
rect 525318 352294 525374 352350
rect 525442 352294 525498 352350
rect 525318 352170 525374 352226
rect 525442 352170 525498 352226
rect 525318 352046 525374 352102
rect 525442 352046 525498 352102
rect 525318 351922 525374 351978
rect 525442 351922 525498 351978
rect 556038 352294 556094 352350
rect 556162 352294 556218 352350
rect 556038 352170 556094 352226
rect 556162 352170 556218 352226
rect 556038 352046 556094 352102
rect 556162 352046 556218 352102
rect 556038 351922 556094 351978
rect 556162 351922 556218 351978
rect 448518 346294 448574 346350
rect 448642 346294 448698 346350
rect 448518 346170 448574 346226
rect 448642 346170 448698 346226
rect 448518 346046 448574 346102
rect 448642 346046 448698 346102
rect 448518 345922 448574 345978
rect 448642 345922 448698 345978
rect 479238 346294 479294 346350
rect 479362 346294 479418 346350
rect 479238 346170 479294 346226
rect 479362 346170 479418 346226
rect 479238 346046 479294 346102
rect 479362 346046 479418 346102
rect 479238 345922 479294 345978
rect 479362 345922 479418 345978
rect 509958 346294 510014 346350
rect 510082 346294 510138 346350
rect 509958 346170 510014 346226
rect 510082 346170 510138 346226
rect 509958 346046 510014 346102
rect 510082 346046 510138 346102
rect 509958 345922 510014 345978
rect 510082 345922 510138 345978
rect 540678 346294 540734 346350
rect 540802 346294 540858 346350
rect 540678 346170 540734 346226
rect 540802 346170 540858 346226
rect 540678 346046 540734 346102
rect 540802 346046 540858 346102
rect 540678 345922 540734 345978
rect 540802 345922 540858 345978
rect 571398 346294 571454 346350
rect 571522 346294 571578 346350
rect 571398 346170 571454 346226
rect 571522 346170 571578 346226
rect 571398 346046 571454 346102
rect 571522 346046 571578 346102
rect 571398 345922 571454 345978
rect 571522 345922 571578 345978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 463878 334294 463934 334350
rect 464002 334294 464058 334350
rect 463878 334170 463934 334226
rect 464002 334170 464058 334226
rect 463878 334046 463934 334102
rect 464002 334046 464058 334102
rect 463878 333922 463934 333978
rect 464002 333922 464058 333978
rect 494598 334294 494654 334350
rect 494722 334294 494778 334350
rect 494598 334170 494654 334226
rect 494722 334170 494778 334226
rect 494598 334046 494654 334102
rect 494722 334046 494778 334102
rect 494598 333922 494654 333978
rect 494722 333922 494778 333978
rect 525318 334294 525374 334350
rect 525442 334294 525498 334350
rect 525318 334170 525374 334226
rect 525442 334170 525498 334226
rect 525318 334046 525374 334102
rect 525442 334046 525498 334102
rect 525318 333922 525374 333978
rect 525442 333922 525498 333978
rect 556038 334294 556094 334350
rect 556162 334294 556218 334350
rect 556038 334170 556094 334226
rect 556162 334170 556218 334226
rect 556038 334046 556094 334102
rect 556162 334046 556218 334102
rect 556038 333922 556094 333978
rect 556162 333922 556218 333978
rect 448518 328294 448574 328350
rect 448642 328294 448698 328350
rect 448518 328170 448574 328226
rect 448642 328170 448698 328226
rect 448518 328046 448574 328102
rect 448642 328046 448698 328102
rect 448518 327922 448574 327978
rect 448642 327922 448698 327978
rect 479238 328294 479294 328350
rect 479362 328294 479418 328350
rect 479238 328170 479294 328226
rect 479362 328170 479418 328226
rect 479238 328046 479294 328102
rect 479362 328046 479418 328102
rect 479238 327922 479294 327978
rect 479362 327922 479418 327978
rect 509958 328294 510014 328350
rect 510082 328294 510138 328350
rect 509958 328170 510014 328226
rect 510082 328170 510138 328226
rect 509958 328046 510014 328102
rect 510082 328046 510138 328102
rect 509958 327922 510014 327978
rect 510082 327922 510138 327978
rect 540678 328294 540734 328350
rect 540802 328294 540858 328350
rect 540678 328170 540734 328226
rect 540802 328170 540858 328226
rect 540678 328046 540734 328102
rect 540802 328046 540858 328102
rect 540678 327922 540734 327978
rect 540802 327922 540858 327978
rect 571398 328294 571454 328350
rect 571522 328294 571578 328350
rect 571398 328170 571454 328226
rect 571522 328170 571578 328226
rect 571398 328046 571454 328102
rect 571522 328046 571578 328102
rect 571398 327922 571454 327978
rect 571522 327922 571578 327978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 463878 316294 463934 316350
rect 464002 316294 464058 316350
rect 463878 316170 463934 316226
rect 464002 316170 464058 316226
rect 463878 316046 463934 316102
rect 464002 316046 464058 316102
rect 463878 315922 463934 315978
rect 464002 315922 464058 315978
rect 494598 316294 494654 316350
rect 494722 316294 494778 316350
rect 494598 316170 494654 316226
rect 494722 316170 494778 316226
rect 494598 316046 494654 316102
rect 494722 316046 494778 316102
rect 494598 315922 494654 315978
rect 494722 315922 494778 315978
rect 525318 316294 525374 316350
rect 525442 316294 525498 316350
rect 525318 316170 525374 316226
rect 525442 316170 525498 316226
rect 525318 316046 525374 316102
rect 525442 316046 525498 316102
rect 525318 315922 525374 315978
rect 525442 315922 525498 315978
rect 556038 316294 556094 316350
rect 556162 316294 556218 316350
rect 556038 316170 556094 316226
rect 556162 316170 556218 316226
rect 556038 316046 556094 316102
rect 556162 316046 556218 316102
rect 556038 315922 556094 315978
rect 556162 315922 556218 315978
rect 448518 310294 448574 310350
rect 448642 310294 448698 310350
rect 448518 310170 448574 310226
rect 448642 310170 448698 310226
rect 448518 310046 448574 310102
rect 448642 310046 448698 310102
rect 448518 309922 448574 309978
rect 448642 309922 448698 309978
rect 479238 310294 479294 310350
rect 479362 310294 479418 310350
rect 479238 310170 479294 310226
rect 479362 310170 479418 310226
rect 479238 310046 479294 310102
rect 479362 310046 479418 310102
rect 479238 309922 479294 309978
rect 479362 309922 479418 309978
rect 509958 310294 510014 310350
rect 510082 310294 510138 310350
rect 509958 310170 510014 310226
rect 510082 310170 510138 310226
rect 509958 310046 510014 310102
rect 510082 310046 510138 310102
rect 509958 309922 510014 309978
rect 510082 309922 510138 309978
rect 540678 310294 540734 310350
rect 540802 310294 540858 310350
rect 540678 310170 540734 310226
rect 540802 310170 540858 310226
rect 540678 310046 540734 310102
rect 540802 310046 540858 310102
rect 540678 309922 540734 309978
rect 540802 309922 540858 309978
rect 571398 310294 571454 310350
rect 571522 310294 571578 310350
rect 571398 310170 571454 310226
rect 571522 310170 571578 310226
rect 571398 310046 571454 310102
rect 571522 310046 571578 310102
rect 571398 309922 571454 309978
rect 571522 309922 571578 309978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 463878 298294 463934 298350
rect 464002 298294 464058 298350
rect 463878 298170 463934 298226
rect 464002 298170 464058 298226
rect 463878 298046 463934 298102
rect 464002 298046 464058 298102
rect 463878 297922 463934 297978
rect 464002 297922 464058 297978
rect 494598 298294 494654 298350
rect 494722 298294 494778 298350
rect 494598 298170 494654 298226
rect 494722 298170 494778 298226
rect 494598 298046 494654 298102
rect 494722 298046 494778 298102
rect 494598 297922 494654 297978
rect 494722 297922 494778 297978
rect 525318 298294 525374 298350
rect 525442 298294 525498 298350
rect 525318 298170 525374 298226
rect 525442 298170 525498 298226
rect 525318 298046 525374 298102
rect 525442 298046 525498 298102
rect 525318 297922 525374 297978
rect 525442 297922 525498 297978
rect 556038 298294 556094 298350
rect 556162 298294 556218 298350
rect 556038 298170 556094 298226
rect 556162 298170 556218 298226
rect 556038 298046 556094 298102
rect 556162 298046 556218 298102
rect 556038 297922 556094 297978
rect 556162 297922 556218 297978
rect 448518 292294 448574 292350
rect 448642 292294 448698 292350
rect 448518 292170 448574 292226
rect 448642 292170 448698 292226
rect 448518 292046 448574 292102
rect 448642 292046 448698 292102
rect 448518 291922 448574 291978
rect 448642 291922 448698 291978
rect 479238 292294 479294 292350
rect 479362 292294 479418 292350
rect 479238 292170 479294 292226
rect 479362 292170 479418 292226
rect 479238 292046 479294 292102
rect 479362 292046 479418 292102
rect 479238 291922 479294 291978
rect 479362 291922 479418 291978
rect 509958 292294 510014 292350
rect 510082 292294 510138 292350
rect 509958 292170 510014 292226
rect 510082 292170 510138 292226
rect 509958 292046 510014 292102
rect 510082 292046 510138 292102
rect 509958 291922 510014 291978
rect 510082 291922 510138 291978
rect 540678 292294 540734 292350
rect 540802 292294 540858 292350
rect 540678 292170 540734 292226
rect 540802 292170 540858 292226
rect 540678 292046 540734 292102
rect 540802 292046 540858 292102
rect 540678 291922 540734 291978
rect 540802 291922 540858 291978
rect 571398 292294 571454 292350
rect 571522 292294 571578 292350
rect 571398 292170 571454 292226
rect 571522 292170 571578 292226
rect 571398 292046 571454 292102
rect 571522 292046 571578 292102
rect 571398 291922 571454 291978
rect 571522 291922 571578 291978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 463878 280294 463934 280350
rect 464002 280294 464058 280350
rect 463878 280170 463934 280226
rect 464002 280170 464058 280226
rect 463878 280046 463934 280102
rect 464002 280046 464058 280102
rect 463878 279922 463934 279978
rect 464002 279922 464058 279978
rect 494598 280294 494654 280350
rect 494722 280294 494778 280350
rect 494598 280170 494654 280226
rect 494722 280170 494778 280226
rect 494598 280046 494654 280102
rect 494722 280046 494778 280102
rect 494598 279922 494654 279978
rect 494722 279922 494778 279978
rect 525318 280294 525374 280350
rect 525442 280294 525498 280350
rect 525318 280170 525374 280226
rect 525442 280170 525498 280226
rect 525318 280046 525374 280102
rect 525442 280046 525498 280102
rect 525318 279922 525374 279978
rect 525442 279922 525498 279978
rect 556038 280294 556094 280350
rect 556162 280294 556218 280350
rect 556038 280170 556094 280226
rect 556162 280170 556218 280226
rect 556038 280046 556094 280102
rect 556162 280046 556218 280102
rect 556038 279922 556094 279978
rect 556162 279922 556218 279978
rect 448518 274294 448574 274350
rect 448642 274294 448698 274350
rect 448518 274170 448574 274226
rect 448642 274170 448698 274226
rect 448518 274046 448574 274102
rect 448642 274046 448698 274102
rect 448518 273922 448574 273978
rect 448642 273922 448698 273978
rect 479238 274294 479294 274350
rect 479362 274294 479418 274350
rect 479238 274170 479294 274226
rect 479362 274170 479418 274226
rect 479238 274046 479294 274102
rect 479362 274046 479418 274102
rect 479238 273922 479294 273978
rect 479362 273922 479418 273978
rect 509958 274294 510014 274350
rect 510082 274294 510138 274350
rect 509958 274170 510014 274226
rect 510082 274170 510138 274226
rect 509958 274046 510014 274102
rect 510082 274046 510138 274102
rect 509958 273922 510014 273978
rect 510082 273922 510138 273978
rect 540678 274294 540734 274350
rect 540802 274294 540858 274350
rect 540678 274170 540734 274226
rect 540802 274170 540858 274226
rect 540678 274046 540734 274102
rect 540802 274046 540858 274102
rect 540678 273922 540734 273978
rect 540802 273922 540858 273978
rect 571398 274294 571454 274350
rect 571522 274294 571578 274350
rect 571398 274170 571454 274226
rect 571522 274170 571578 274226
rect 571398 274046 571454 274102
rect 571522 274046 571578 274102
rect 571398 273922 571454 273978
rect 571522 273922 571578 273978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 463878 262294 463934 262350
rect 464002 262294 464058 262350
rect 463878 262170 463934 262226
rect 464002 262170 464058 262226
rect 463878 262046 463934 262102
rect 464002 262046 464058 262102
rect 463878 261922 463934 261978
rect 464002 261922 464058 261978
rect 494598 262294 494654 262350
rect 494722 262294 494778 262350
rect 494598 262170 494654 262226
rect 494722 262170 494778 262226
rect 494598 262046 494654 262102
rect 494722 262046 494778 262102
rect 494598 261922 494654 261978
rect 494722 261922 494778 261978
rect 525318 262294 525374 262350
rect 525442 262294 525498 262350
rect 525318 262170 525374 262226
rect 525442 262170 525498 262226
rect 525318 262046 525374 262102
rect 525442 262046 525498 262102
rect 525318 261922 525374 261978
rect 525442 261922 525498 261978
rect 556038 262294 556094 262350
rect 556162 262294 556218 262350
rect 556038 262170 556094 262226
rect 556162 262170 556218 262226
rect 556038 262046 556094 262102
rect 556162 262046 556218 262102
rect 556038 261922 556094 261978
rect 556162 261922 556218 261978
rect 448518 256294 448574 256350
rect 448642 256294 448698 256350
rect 448518 256170 448574 256226
rect 448642 256170 448698 256226
rect 448518 256046 448574 256102
rect 448642 256046 448698 256102
rect 448518 255922 448574 255978
rect 448642 255922 448698 255978
rect 479238 256294 479294 256350
rect 479362 256294 479418 256350
rect 479238 256170 479294 256226
rect 479362 256170 479418 256226
rect 479238 256046 479294 256102
rect 479362 256046 479418 256102
rect 479238 255922 479294 255978
rect 479362 255922 479418 255978
rect 509958 256294 510014 256350
rect 510082 256294 510138 256350
rect 509958 256170 510014 256226
rect 510082 256170 510138 256226
rect 509958 256046 510014 256102
rect 510082 256046 510138 256102
rect 509958 255922 510014 255978
rect 510082 255922 510138 255978
rect 540678 256294 540734 256350
rect 540802 256294 540858 256350
rect 540678 256170 540734 256226
rect 540802 256170 540858 256226
rect 540678 256046 540734 256102
rect 540802 256046 540858 256102
rect 540678 255922 540734 255978
rect 540802 255922 540858 255978
rect 571398 256294 571454 256350
rect 571522 256294 571578 256350
rect 571398 256170 571454 256226
rect 571522 256170 571578 256226
rect 571398 256046 571454 256102
rect 571522 256046 571578 256102
rect 571398 255922 571454 255978
rect 571522 255922 571578 255978
rect 463878 244294 463934 244350
rect 464002 244294 464058 244350
rect 463878 244170 463934 244226
rect 464002 244170 464058 244226
rect 463878 244046 463934 244102
rect 464002 244046 464058 244102
rect 463878 243922 463934 243978
rect 464002 243922 464058 243978
rect 494598 244294 494654 244350
rect 494722 244294 494778 244350
rect 494598 244170 494654 244226
rect 494722 244170 494778 244226
rect 494598 244046 494654 244102
rect 494722 244046 494778 244102
rect 494598 243922 494654 243978
rect 494722 243922 494778 243978
rect 525318 244294 525374 244350
rect 525442 244294 525498 244350
rect 525318 244170 525374 244226
rect 525442 244170 525498 244226
rect 525318 244046 525374 244102
rect 525442 244046 525498 244102
rect 525318 243922 525374 243978
rect 525442 243922 525498 243978
rect 556038 244294 556094 244350
rect 556162 244294 556218 244350
rect 556038 244170 556094 244226
rect 556162 244170 556218 244226
rect 556038 244046 556094 244102
rect 556162 244046 556218 244102
rect 556038 243922 556094 243978
rect 556162 243922 556218 243978
rect 448518 238294 448574 238350
rect 448642 238294 448698 238350
rect 448518 238170 448574 238226
rect 448642 238170 448698 238226
rect 448518 238046 448574 238102
rect 448642 238046 448698 238102
rect 448518 237922 448574 237978
rect 448642 237922 448698 237978
rect 479238 238294 479294 238350
rect 479362 238294 479418 238350
rect 479238 238170 479294 238226
rect 479362 238170 479418 238226
rect 479238 238046 479294 238102
rect 479362 238046 479418 238102
rect 479238 237922 479294 237978
rect 479362 237922 479418 237978
rect 509958 238294 510014 238350
rect 510082 238294 510138 238350
rect 509958 238170 510014 238226
rect 510082 238170 510138 238226
rect 509958 238046 510014 238102
rect 510082 238046 510138 238102
rect 509958 237922 510014 237978
rect 510082 237922 510138 237978
rect 540678 238294 540734 238350
rect 540802 238294 540858 238350
rect 540678 238170 540734 238226
rect 540802 238170 540858 238226
rect 540678 238046 540734 238102
rect 540802 238046 540858 238102
rect 540678 237922 540734 237978
rect 540802 237922 540858 237978
rect 571398 238294 571454 238350
rect 571522 238294 571578 238350
rect 571398 238170 571454 238226
rect 571522 238170 571578 238226
rect 571398 238046 571454 238102
rect 571522 238046 571578 238102
rect 571398 237922 571454 237978
rect 571522 237922 571578 237978
rect 463878 226294 463934 226350
rect 464002 226294 464058 226350
rect 463878 226170 463934 226226
rect 464002 226170 464058 226226
rect 463878 226046 463934 226102
rect 464002 226046 464058 226102
rect 463878 225922 463934 225978
rect 464002 225922 464058 225978
rect 494598 226294 494654 226350
rect 494722 226294 494778 226350
rect 494598 226170 494654 226226
rect 494722 226170 494778 226226
rect 494598 226046 494654 226102
rect 494722 226046 494778 226102
rect 494598 225922 494654 225978
rect 494722 225922 494778 225978
rect 525318 226294 525374 226350
rect 525442 226294 525498 226350
rect 525318 226170 525374 226226
rect 525442 226170 525498 226226
rect 525318 226046 525374 226102
rect 525442 226046 525498 226102
rect 525318 225922 525374 225978
rect 525442 225922 525498 225978
rect 556038 226294 556094 226350
rect 556162 226294 556218 226350
rect 556038 226170 556094 226226
rect 556162 226170 556218 226226
rect 556038 226046 556094 226102
rect 556162 226046 556218 226102
rect 556038 225922 556094 225978
rect 556162 225922 556218 225978
rect 448518 220294 448574 220350
rect 448642 220294 448698 220350
rect 448518 220170 448574 220226
rect 448642 220170 448698 220226
rect 448518 220046 448574 220102
rect 448642 220046 448698 220102
rect 448518 219922 448574 219978
rect 448642 219922 448698 219978
rect 479238 220294 479294 220350
rect 479362 220294 479418 220350
rect 479238 220170 479294 220226
rect 479362 220170 479418 220226
rect 479238 220046 479294 220102
rect 479362 220046 479418 220102
rect 479238 219922 479294 219978
rect 479362 219922 479418 219978
rect 509958 220294 510014 220350
rect 510082 220294 510138 220350
rect 509958 220170 510014 220226
rect 510082 220170 510138 220226
rect 509958 220046 510014 220102
rect 510082 220046 510138 220102
rect 509958 219922 510014 219978
rect 510082 219922 510138 219978
rect 540678 220294 540734 220350
rect 540802 220294 540858 220350
rect 540678 220170 540734 220226
rect 540802 220170 540858 220226
rect 540678 220046 540734 220102
rect 540802 220046 540858 220102
rect 540678 219922 540734 219978
rect 540802 219922 540858 219978
rect 571398 220294 571454 220350
rect 571522 220294 571578 220350
rect 571398 220170 571454 220226
rect 571522 220170 571578 220226
rect 571398 220046 571454 220102
rect 571522 220046 571578 220102
rect 571398 219922 571454 219978
rect 571522 219922 571578 219978
rect 463878 208294 463934 208350
rect 464002 208294 464058 208350
rect 463878 208170 463934 208226
rect 464002 208170 464058 208226
rect 463878 208046 463934 208102
rect 464002 208046 464058 208102
rect 463878 207922 463934 207978
rect 464002 207922 464058 207978
rect 494598 208294 494654 208350
rect 494722 208294 494778 208350
rect 494598 208170 494654 208226
rect 494722 208170 494778 208226
rect 494598 208046 494654 208102
rect 494722 208046 494778 208102
rect 494598 207922 494654 207978
rect 494722 207922 494778 207978
rect 525318 208294 525374 208350
rect 525442 208294 525498 208350
rect 525318 208170 525374 208226
rect 525442 208170 525498 208226
rect 525318 208046 525374 208102
rect 525442 208046 525498 208102
rect 525318 207922 525374 207978
rect 525442 207922 525498 207978
rect 556038 208294 556094 208350
rect 556162 208294 556218 208350
rect 556038 208170 556094 208226
rect 556162 208170 556218 208226
rect 556038 208046 556094 208102
rect 556162 208046 556218 208102
rect 556038 207922 556094 207978
rect 556162 207922 556218 207978
rect 448518 202294 448574 202350
rect 448642 202294 448698 202350
rect 448518 202170 448574 202226
rect 448642 202170 448698 202226
rect 448518 202046 448574 202102
rect 448642 202046 448698 202102
rect 448518 201922 448574 201978
rect 448642 201922 448698 201978
rect 479238 202294 479294 202350
rect 479362 202294 479418 202350
rect 479238 202170 479294 202226
rect 479362 202170 479418 202226
rect 479238 202046 479294 202102
rect 479362 202046 479418 202102
rect 479238 201922 479294 201978
rect 479362 201922 479418 201978
rect 509958 202294 510014 202350
rect 510082 202294 510138 202350
rect 509958 202170 510014 202226
rect 510082 202170 510138 202226
rect 509958 202046 510014 202102
rect 510082 202046 510138 202102
rect 509958 201922 510014 201978
rect 510082 201922 510138 201978
rect 540678 202294 540734 202350
rect 540802 202294 540858 202350
rect 540678 202170 540734 202226
rect 540802 202170 540858 202226
rect 540678 202046 540734 202102
rect 540802 202046 540858 202102
rect 540678 201922 540734 201978
rect 540802 201922 540858 201978
rect 571398 202294 571454 202350
rect 571522 202294 571578 202350
rect 571398 202170 571454 202226
rect 571522 202170 571578 202226
rect 571398 202046 571454 202102
rect 571522 202046 571578 202102
rect 571398 201922 571454 201978
rect 571522 201922 571578 201978
rect 463878 190294 463934 190350
rect 464002 190294 464058 190350
rect 463878 190170 463934 190226
rect 464002 190170 464058 190226
rect 463878 190046 463934 190102
rect 464002 190046 464058 190102
rect 463878 189922 463934 189978
rect 464002 189922 464058 189978
rect 494598 190294 494654 190350
rect 494722 190294 494778 190350
rect 494598 190170 494654 190226
rect 494722 190170 494778 190226
rect 494598 190046 494654 190102
rect 494722 190046 494778 190102
rect 494598 189922 494654 189978
rect 494722 189922 494778 189978
rect 525318 190294 525374 190350
rect 525442 190294 525498 190350
rect 525318 190170 525374 190226
rect 525442 190170 525498 190226
rect 525318 190046 525374 190102
rect 525442 190046 525498 190102
rect 525318 189922 525374 189978
rect 525442 189922 525498 189978
rect 556038 190294 556094 190350
rect 556162 190294 556218 190350
rect 556038 190170 556094 190226
rect 556162 190170 556218 190226
rect 556038 190046 556094 190102
rect 556162 190046 556218 190102
rect 556038 189922 556094 189978
rect 556162 189922 556218 189978
rect 448518 184294 448574 184350
rect 448642 184294 448698 184350
rect 448518 184170 448574 184226
rect 448642 184170 448698 184226
rect 448518 184046 448574 184102
rect 448642 184046 448698 184102
rect 448518 183922 448574 183978
rect 448642 183922 448698 183978
rect 479238 184294 479294 184350
rect 479362 184294 479418 184350
rect 479238 184170 479294 184226
rect 479362 184170 479418 184226
rect 479238 184046 479294 184102
rect 479362 184046 479418 184102
rect 479238 183922 479294 183978
rect 479362 183922 479418 183978
rect 509958 184294 510014 184350
rect 510082 184294 510138 184350
rect 509958 184170 510014 184226
rect 510082 184170 510138 184226
rect 509958 184046 510014 184102
rect 510082 184046 510138 184102
rect 509958 183922 510014 183978
rect 510082 183922 510138 183978
rect 540678 184294 540734 184350
rect 540802 184294 540858 184350
rect 540678 184170 540734 184226
rect 540802 184170 540858 184226
rect 540678 184046 540734 184102
rect 540802 184046 540858 184102
rect 540678 183922 540734 183978
rect 540802 183922 540858 183978
rect 571398 184294 571454 184350
rect 571522 184294 571578 184350
rect 571398 184170 571454 184226
rect 571522 184170 571578 184226
rect 571398 184046 571454 184102
rect 571522 184046 571578 184102
rect 571398 183922 571454 183978
rect 571522 183922 571578 183978
rect 463878 172294 463934 172350
rect 464002 172294 464058 172350
rect 463878 172170 463934 172226
rect 464002 172170 464058 172226
rect 463878 172046 463934 172102
rect 464002 172046 464058 172102
rect 463878 171922 463934 171978
rect 464002 171922 464058 171978
rect 494598 172294 494654 172350
rect 494722 172294 494778 172350
rect 494598 172170 494654 172226
rect 494722 172170 494778 172226
rect 494598 172046 494654 172102
rect 494722 172046 494778 172102
rect 494598 171922 494654 171978
rect 494722 171922 494778 171978
rect 525318 172294 525374 172350
rect 525442 172294 525498 172350
rect 525318 172170 525374 172226
rect 525442 172170 525498 172226
rect 525318 172046 525374 172102
rect 525442 172046 525498 172102
rect 525318 171922 525374 171978
rect 525442 171922 525498 171978
rect 556038 172294 556094 172350
rect 556162 172294 556218 172350
rect 556038 172170 556094 172226
rect 556162 172170 556218 172226
rect 556038 172046 556094 172102
rect 556162 172046 556218 172102
rect 556038 171922 556094 171978
rect 556162 171922 556218 171978
rect 448518 166294 448574 166350
rect 448642 166294 448698 166350
rect 448518 166170 448574 166226
rect 448642 166170 448698 166226
rect 448518 166046 448574 166102
rect 448642 166046 448698 166102
rect 448518 165922 448574 165978
rect 448642 165922 448698 165978
rect 479238 166294 479294 166350
rect 479362 166294 479418 166350
rect 479238 166170 479294 166226
rect 479362 166170 479418 166226
rect 479238 166046 479294 166102
rect 479362 166046 479418 166102
rect 479238 165922 479294 165978
rect 479362 165922 479418 165978
rect 509958 166294 510014 166350
rect 510082 166294 510138 166350
rect 509958 166170 510014 166226
rect 510082 166170 510138 166226
rect 509958 166046 510014 166102
rect 510082 166046 510138 166102
rect 509958 165922 510014 165978
rect 510082 165922 510138 165978
rect 540678 166294 540734 166350
rect 540802 166294 540858 166350
rect 540678 166170 540734 166226
rect 540802 166170 540858 166226
rect 540678 166046 540734 166102
rect 540802 166046 540858 166102
rect 540678 165922 540734 165978
rect 540802 165922 540858 165978
rect 571398 166294 571454 166350
rect 571522 166294 571578 166350
rect 571398 166170 571454 166226
rect 571522 166170 571578 166226
rect 571398 166046 571454 166102
rect 571522 166046 571578 166102
rect 571398 165922 571454 165978
rect 571522 165922 571578 165978
rect 463878 154294 463934 154350
rect 464002 154294 464058 154350
rect 463878 154170 463934 154226
rect 464002 154170 464058 154226
rect 463878 154046 463934 154102
rect 464002 154046 464058 154102
rect 463878 153922 463934 153978
rect 464002 153922 464058 153978
rect 494598 154294 494654 154350
rect 494722 154294 494778 154350
rect 494598 154170 494654 154226
rect 494722 154170 494778 154226
rect 494598 154046 494654 154102
rect 494722 154046 494778 154102
rect 494598 153922 494654 153978
rect 494722 153922 494778 153978
rect 525318 154294 525374 154350
rect 525442 154294 525498 154350
rect 525318 154170 525374 154226
rect 525442 154170 525498 154226
rect 525318 154046 525374 154102
rect 525442 154046 525498 154102
rect 525318 153922 525374 153978
rect 525442 153922 525498 153978
rect 556038 154294 556094 154350
rect 556162 154294 556218 154350
rect 556038 154170 556094 154226
rect 556162 154170 556218 154226
rect 556038 154046 556094 154102
rect 556162 154046 556218 154102
rect 556038 153922 556094 153978
rect 556162 153922 556218 153978
rect 448518 148294 448574 148350
rect 448642 148294 448698 148350
rect 448518 148170 448574 148226
rect 448642 148170 448698 148226
rect 448518 148046 448574 148102
rect 448642 148046 448698 148102
rect 448518 147922 448574 147978
rect 448642 147922 448698 147978
rect 479238 148294 479294 148350
rect 479362 148294 479418 148350
rect 479238 148170 479294 148226
rect 479362 148170 479418 148226
rect 479238 148046 479294 148102
rect 479362 148046 479418 148102
rect 479238 147922 479294 147978
rect 479362 147922 479418 147978
rect 509958 148294 510014 148350
rect 510082 148294 510138 148350
rect 509958 148170 510014 148226
rect 510082 148170 510138 148226
rect 509958 148046 510014 148102
rect 510082 148046 510138 148102
rect 509958 147922 510014 147978
rect 510082 147922 510138 147978
rect 540678 148294 540734 148350
rect 540802 148294 540858 148350
rect 540678 148170 540734 148226
rect 540802 148170 540858 148226
rect 540678 148046 540734 148102
rect 540802 148046 540858 148102
rect 540678 147922 540734 147978
rect 540802 147922 540858 147978
rect 571398 148294 571454 148350
rect 571522 148294 571578 148350
rect 571398 148170 571454 148226
rect 571522 148170 571578 148226
rect 571398 148046 571454 148102
rect 571522 148046 571578 148102
rect 571398 147922 571454 147978
rect 571522 147922 571578 147978
rect 463878 136294 463934 136350
rect 464002 136294 464058 136350
rect 463878 136170 463934 136226
rect 464002 136170 464058 136226
rect 463878 136046 463934 136102
rect 464002 136046 464058 136102
rect 463878 135922 463934 135978
rect 464002 135922 464058 135978
rect 494598 136294 494654 136350
rect 494722 136294 494778 136350
rect 494598 136170 494654 136226
rect 494722 136170 494778 136226
rect 494598 136046 494654 136102
rect 494722 136046 494778 136102
rect 494598 135922 494654 135978
rect 494722 135922 494778 135978
rect 525318 136294 525374 136350
rect 525442 136294 525498 136350
rect 525318 136170 525374 136226
rect 525442 136170 525498 136226
rect 525318 136046 525374 136102
rect 525442 136046 525498 136102
rect 525318 135922 525374 135978
rect 525442 135922 525498 135978
rect 556038 136294 556094 136350
rect 556162 136294 556218 136350
rect 556038 136170 556094 136226
rect 556162 136170 556218 136226
rect 556038 136046 556094 136102
rect 556162 136046 556218 136102
rect 556038 135922 556094 135978
rect 556162 135922 556218 135978
rect 448518 130294 448574 130350
rect 448642 130294 448698 130350
rect 448518 130170 448574 130226
rect 448642 130170 448698 130226
rect 448518 130046 448574 130102
rect 448642 130046 448698 130102
rect 448518 129922 448574 129978
rect 448642 129922 448698 129978
rect 479238 130294 479294 130350
rect 479362 130294 479418 130350
rect 479238 130170 479294 130226
rect 479362 130170 479418 130226
rect 479238 130046 479294 130102
rect 479362 130046 479418 130102
rect 479238 129922 479294 129978
rect 479362 129922 479418 129978
rect 509958 130294 510014 130350
rect 510082 130294 510138 130350
rect 509958 130170 510014 130226
rect 510082 130170 510138 130226
rect 509958 130046 510014 130102
rect 510082 130046 510138 130102
rect 509958 129922 510014 129978
rect 510082 129922 510138 129978
rect 540678 130294 540734 130350
rect 540802 130294 540858 130350
rect 540678 130170 540734 130226
rect 540802 130170 540858 130226
rect 540678 130046 540734 130102
rect 540802 130046 540858 130102
rect 540678 129922 540734 129978
rect 540802 129922 540858 129978
rect 571398 130294 571454 130350
rect 571522 130294 571578 130350
rect 571398 130170 571454 130226
rect 571522 130170 571578 130226
rect 571398 130046 571454 130102
rect 571522 130046 571578 130102
rect 571398 129922 571454 129978
rect 571522 129922 571578 129978
rect 463878 118294 463934 118350
rect 464002 118294 464058 118350
rect 463878 118170 463934 118226
rect 464002 118170 464058 118226
rect 463878 118046 463934 118102
rect 464002 118046 464058 118102
rect 463878 117922 463934 117978
rect 464002 117922 464058 117978
rect 494598 118294 494654 118350
rect 494722 118294 494778 118350
rect 494598 118170 494654 118226
rect 494722 118170 494778 118226
rect 494598 118046 494654 118102
rect 494722 118046 494778 118102
rect 494598 117922 494654 117978
rect 494722 117922 494778 117978
rect 525318 118294 525374 118350
rect 525442 118294 525498 118350
rect 525318 118170 525374 118226
rect 525442 118170 525498 118226
rect 525318 118046 525374 118102
rect 525442 118046 525498 118102
rect 525318 117922 525374 117978
rect 525442 117922 525498 117978
rect 556038 118294 556094 118350
rect 556162 118294 556218 118350
rect 556038 118170 556094 118226
rect 556162 118170 556218 118226
rect 556038 118046 556094 118102
rect 556162 118046 556218 118102
rect 556038 117922 556094 117978
rect 556162 117922 556218 117978
rect 448518 112294 448574 112350
rect 448642 112294 448698 112350
rect 448518 112170 448574 112226
rect 448642 112170 448698 112226
rect 448518 112046 448574 112102
rect 448642 112046 448698 112102
rect 448518 111922 448574 111978
rect 448642 111922 448698 111978
rect 479238 112294 479294 112350
rect 479362 112294 479418 112350
rect 479238 112170 479294 112226
rect 479362 112170 479418 112226
rect 479238 112046 479294 112102
rect 479362 112046 479418 112102
rect 479238 111922 479294 111978
rect 479362 111922 479418 111978
rect 509958 112294 510014 112350
rect 510082 112294 510138 112350
rect 509958 112170 510014 112226
rect 510082 112170 510138 112226
rect 509958 112046 510014 112102
rect 510082 112046 510138 112102
rect 509958 111922 510014 111978
rect 510082 111922 510138 111978
rect 540678 112294 540734 112350
rect 540802 112294 540858 112350
rect 540678 112170 540734 112226
rect 540802 112170 540858 112226
rect 540678 112046 540734 112102
rect 540802 112046 540858 112102
rect 540678 111922 540734 111978
rect 540802 111922 540858 111978
rect 571398 112294 571454 112350
rect 571522 112294 571578 112350
rect 571398 112170 571454 112226
rect 571522 112170 571578 112226
rect 571398 112046 571454 112102
rect 571522 112046 571578 112102
rect 571398 111922 571454 111978
rect 571522 111922 571578 111978
rect 443436 101582 443492 101638
rect 463878 100294 463934 100350
rect 464002 100294 464058 100350
rect 463878 100170 463934 100226
rect 464002 100170 464058 100226
rect 463878 100046 463934 100102
rect 464002 100046 464058 100102
rect 463878 99922 463934 99978
rect 464002 99922 464058 99978
rect 494598 100294 494654 100350
rect 494722 100294 494778 100350
rect 494598 100170 494654 100226
rect 494722 100170 494778 100226
rect 494598 100046 494654 100102
rect 494722 100046 494778 100102
rect 494598 99922 494654 99978
rect 494722 99922 494778 99978
rect 525318 100294 525374 100350
rect 525442 100294 525498 100350
rect 525318 100170 525374 100226
rect 525442 100170 525498 100226
rect 525318 100046 525374 100102
rect 525442 100046 525498 100102
rect 525318 99922 525374 99978
rect 525442 99922 525498 99978
rect 556038 100294 556094 100350
rect 556162 100294 556218 100350
rect 556038 100170 556094 100226
rect 556162 100170 556218 100226
rect 556038 100046 556094 100102
rect 556162 100046 556218 100102
rect 556038 99922 556094 99978
rect 556162 99922 556218 99978
rect 443100 98162 443156 98218
rect 448518 94294 448574 94350
rect 448642 94294 448698 94350
rect 448518 94170 448574 94226
rect 448642 94170 448698 94226
rect 448518 94046 448574 94102
rect 448642 94046 448698 94102
rect 448518 93922 448574 93978
rect 448642 93922 448698 93978
rect 479238 94294 479294 94350
rect 479362 94294 479418 94350
rect 479238 94170 479294 94226
rect 479362 94170 479418 94226
rect 479238 94046 479294 94102
rect 479362 94046 479418 94102
rect 479238 93922 479294 93978
rect 479362 93922 479418 93978
rect 509958 94294 510014 94350
rect 510082 94294 510138 94350
rect 509958 94170 510014 94226
rect 510082 94170 510138 94226
rect 509958 94046 510014 94102
rect 510082 94046 510138 94102
rect 509958 93922 510014 93978
rect 510082 93922 510138 93978
rect 540678 94294 540734 94350
rect 540802 94294 540858 94350
rect 540678 94170 540734 94226
rect 540802 94170 540858 94226
rect 540678 94046 540734 94102
rect 540802 94046 540858 94102
rect 540678 93922 540734 93978
rect 540802 93922 540858 93978
rect 571398 94294 571454 94350
rect 571522 94294 571578 94350
rect 571398 94170 571454 94226
rect 571522 94170 571578 94226
rect 571398 94046 571454 94102
rect 571522 94046 571578 94102
rect 571398 93922 571454 93978
rect 571522 93922 571578 93978
rect 443100 85742 443156 85798
rect 463878 82294 463934 82350
rect 464002 82294 464058 82350
rect 463878 82170 463934 82226
rect 464002 82170 464058 82226
rect 463878 82046 463934 82102
rect 464002 82046 464058 82102
rect 463878 81922 463934 81978
rect 464002 81922 464058 81978
rect 494598 82294 494654 82350
rect 494722 82294 494778 82350
rect 494598 82170 494654 82226
rect 494722 82170 494778 82226
rect 494598 82046 494654 82102
rect 494722 82046 494778 82102
rect 494598 81922 494654 81978
rect 494722 81922 494778 81978
rect 525318 82294 525374 82350
rect 525442 82294 525498 82350
rect 525318 82170 525374 82226
rect 525442 82170 525498 82226
rect 525318 82046 525374 82102
rect 525442 82046 525498 82102
rect 525318 81922 525374 81978
rect 525442 81922 525498 81978
rect 556038 82294 556094 82350
rect 556162 82294 556218 82350
rect 556038 82170 556094 82226
rect 556162 82170 556218 82226
rect 556038 82046 556094 82102
rect 556162 82046 556218 82102
rect 556038 81922 556094 81978
rect 556162 81922 556218 81978
rect 443212 80702 443268 80758
rect 448518 76294 448574 76350
rect 448642 76294 448698 76350
rect 448518 76170 448574 76226
rect 448642 76170 448698 76226
rect 448518 76046 448574 76102
rect 448642 76046 448698 76102
rect 448518 75922 448574 75978
rect 448642 75922 448698 75978
rect 479238 76294 479294 76350
rect 479362 76294 479418 76350
rect 479238 76170 479294 76226
rect 479362 76170 479418 76226
rect 479238 76046 479294 76102
rect 479362 76046 479418 76102
rect 479238 75922 479294 75978
rect 479362 75922 479418 75978
rect 509958 76294 510014 76350
rect 510082 76294 510138 76350
rect 509958 76170 510014 76226
rect 510082 76170 510138 76226
rect 509958 76046 510014 76102
rect 510082 76046 510138 76102
rect 509958 75922 510014 75978
rect 510082 75922 510138 75978
rect 540678 76294 540734 76350
rect 540802 76294 540858 76350
rect 540678 76170 540734 76226
rect 540802 76170 540858 76226
rect 540678 76046 540734 76102
rect 540802 76046 540858 76102
rect 540678 75922 540734 75978
rect 540802 75922 540858 75978
rect 571398 76294 571454 76350
rect 571522 76294 571578 76350
rect 571398 76170 571454 76226
rect 571522 76170 571578 76226
rect 571398 76046 571454 76102
rect 571522 76046 571578 76102
rect 571398 75922 571454 75978
rect 571522 75922 571578 75978
rect 463878 64294 463934 64350
rect 464002 64294 464058 64350
rect 463878 64170 463934 64226
rect 464002 64170 464058 64226
rect 463878 64046 463934 64102
rect 464002 64046 464058 64102
rect 463878 63922 463934 63978
rect 464002 63922 464058 63978
rect 494598 64294 494654 64350
rect 494722 64294 494778 64350
rect 494598 64170 494654 64226
rect 494722 64170 494778 64226
rect 494598 64046 494654 64102
rect 494722 64046 494778 64102
rect 494598 63922 494654 63978
rect 494722 63922 494778 63978
rect 525318 64294 525374 64350
rect 525442 64294 525498 64350
rect 525318 64170 525374 64226
rect 525442 64170 525498 64226
rect 525318 64046 525374 64102
rect 525442 64046 525498 64102
rect 525318 63922 525374 63978
rect 525442 63922 525498 63978
rect 556038 64294 556094 64350
rect 556162 64294 556218 64350
rect 556038 64170 556094 64226
rect 556162 64170 556218 64226
rect 556038 64046 556094 64102
rect 556162 64046 556218 64102
rect 556038 63922 556094 63978
rect 556162 63922 556218 63978
rect 448518 58294 448574 58350
rect 448642 58294 448698 58350
rect 448518 58170 448574 58226
rect 448642 58170 448698 58226
rect 448518 58046 448574 58102
rect 448642 58046 448698 58102
rect 448518 57922 448574 57978
rect 448642 57922 448698 57978
rect 479238 58294 479294 58350
rect 479362 58294 479418 58350
rect 479238 58170 479294 58226
rect 479362 58170 479418 58226
rect 479238 58046 479294 58102
rect 479362 58046 479418 58102
rect 479238 57922 479294 57978
rect 479362 57922 479418 57978
rect 509958 58294 510014 58350
rect 510082 58294 510138 58350
rect 509958 58170 510014 58226
rect 510082 58170 510138 58226
rect 509958 58046 510014 58102
rect 510082 58046 510138 58102
rect 509958 57922 510014 57978
rect 510082 57922 510138 57978
rect 540678 58294 540734 58350
rect 540802 58294 540858 58350
rect 540678 58170 540734 58226
rect 540802 58170 540858 58226
rect 540678 58046 540734 58102
rect 540802 58046 540858 58102
rect 540678 57922 540734 57978
rect 540802 57922 540858 57978
rect 571398 58294 571454 58350
rect 571522 58294 571578 58350
rect 571398 58170 571454 58226
rect 571522 58170 571578 58226
rect 571398 58046 571454 58102
rect 571522 58046 571578 58102
rect 571398 57922 571454 57978
rect 571522 57922 571578 57978
rect 463878 46294 463934 46350
rect 464002 46294 464058 46350
rect 463878 46170 463934 46226
rect 464002 46170 464058 46226
rect 463878 46046 463934 46102
rect 464002 46046 464058 46102
rect 463878 45922 463934 45978
rect 464002 45922 464058 45978
rect 494598 46294 494654 46350
rect 494722 46294 494778 46350
rect 494598 46170 494654 46226
rect 494722 46170 494778 46226
rect 494598 46046 494654 46102
rect 494722 46046 494778 46102
rect 494598 45922 494654 45978
rect 494722 45922 494778 45978
rect 525318 46294 525374 46350
rect 525442 46294 525498 46350
rect 525318 46170 525374 46226
rect 525442 46170 525498 46226
rect 525318 46046 525374 46102
rect 525442 46046 525498 46102
rect 525318 45922 525374 45978
rect 525442 45922 525498 45978
rect 556038 46294 556094 46350
rect 556162 46294 556218 46350
rect 556038 46170 556094 46226
rect 556162 46170 556218 46226
rect 556038 46046 556094 46102
rect 556162 46046 556218 46102
rect 556038 45922 556094 45978
rect 556162 45922 556218 45978
rect 448518 40294 448574 40350
rect 448642 40294 448698 40350
rect 448518 40170 448574 40226
rect 448642 40170 448698 40226
rect 448518 40046 448574 40102
rect 448642 40046 448698 40102
rect 448518 39922 448574 39978
rect 448642 39922 448698 39978
rect 479238 40294 479294 40350
rect 479362 40294 479418 40350
rect 479238 40170 479294 40226
rect 479362 40170 479418 40226
rect 479238 40046 479294 40102
rect 479362 40046 479418 40102
rect 479238 39922 479294 39978
rect 479362 39922 479418 39978
rect 509958 40294 510014 40350
rect 510082 40294 510138 40350
rect 509958 40170 510014 40226
rect 510082 40170 510138 40226
rect 509958 40046 510014 40102
rect 510082 40046 510138 40102
rect 509958 39922 510014 39978
rect 510082 39922 510138 39978
rect 540678 40294 540734 40350
rect 540802 40294 540858 40350
rect 540678 40170 540734 40226
rect 540802 40170 540858 40226
rect 540678 40046 540734 40102
rect 540802 40046 540858 40102
rect 540678 39922 540734 39978
rect 540802 39922 540858 39978
rect 571398 40294 571454 40350
rect 571522 40294 571578 40350
rect 571398 40170 571454 40226
rect 571522 40170 571578 40226
rect 571398 40046 571454 40102
rect 571522 40046 571578 40102
rect 571398 39922 571454 39978
rect 571522 39922 571578 39978
rect 463878 28294 463934 28350
rect 464002 28294 464058 28350
rect 463878 28170 463934 28226
rect 464002 28170 464058 28226
rect 463878 28046 463934 28102
rect 464002 28046 464058 28102
rect 463878 27922 463934 27978
rect 464002 27922 464058 27978
rect 494598 28294 494654 28350
rect 494722 28294 494778 28350
rect 494598 28170 494654 28226
rect 494722 28170 494778 28226
rect 494598 28046 494654 28102
rect 494722 28046 494778 28102
rect 494598 27922 494654 27978
rect 494722 27922 494778 27978
rect 525318 28294 525374 28350
rect 525442 28294 525498 28350
rect 525318 28170 525374 28226
rect 525442 28170 525498 28226
rect 525318 28046 525374 28102
rect 525442 28046 525498 28102
rect 525318 27922 525374 27978
rect 525442 27922 525498 27978
rect 556038 28294 556094 28350
rect 556162 28294 556218 28350
rect 556038 28170 556094 28226
rect 556162 28170 556218 28226
rect 556038 28046 556094 28102
rect 556162 28046 556218 28102
rect 556038 27922 556094 27978
rect 556162 27922 556218 27978
rect 587132 20042 587188 20098
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 479724 7982 479780 8038
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 475916 2762 475972 2818
rect 474012 782 474068 838
rect 485548 644 485604 658
rect 485548 602 485604 644
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 523516 8522 523572 8578
rect 506380 6362 506436 6418
rect 512092 6182 512148 6238
rect 517804 6002 517860 6058
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 531132 9422 531188 9478
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 515900 3122 515956 3178
rect 527324 242 527380 298
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 540652 7802 540708 7858
rect 534940 5822 534996 5878
rect 546364 7622 546420 7678
rect 557788 7442 557844 7498
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 552636 3302 552692 3358
rect 542668 2942 542724 2998
rect 553980 422 554036 478
rect 533036 62 533092 118
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 559692 4742 559748 4798
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 581308 15902 581364 15958
rect 571228 9242 571284 9298
rect 571228 4922 571284 4978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 17816 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 17816 586350
rect -1916 586226 17816 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 17816 586226
rect -1916 586102 17816 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 17816 586102
rect -1916 585978 17816 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 17816 585978
rect -1916 585826 17816 585922
rect 170184 586350 597980 586446
rect 170184 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 170184 586226 597980 586294
rect 170184 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 170184 586102 597980 586170
rect 170184 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 170184 585978 597980 586046
rect 170184 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 170184 585826 597980 585922
rect -1916 580350 17816 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 17816 580350
rect -1916 580226 17816 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 17816 580226
rect -1916 580102 17816 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 17816 580102
rect -1916 579978 17816 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 17816 579978
rect -1916 579826 17816 579922
rect 170184 580350 597980 580446
rect 170184 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect 170184 580226 597980 580294
rect 170184 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect 170184 580102 597980 580170
rect 170184 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect 170184 579978 597980 580046
rect 170184 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect 170184 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 37878 568350
rect 37934 568294 38002 568350
rect 38058 568294 68598 568350
rect 68654 568294 68722 568350
rect 68778 568294 99318 568350
rect 99374 568294 99442 568350
rect 99498 568294 130038 568350
rect 130094 568294 130162 568350
rect 130218 568294 160758 568350
rect 160814 568294 160882 568350
rect 160938 568294 191478 568350
rect 191534 568294 191602 568350
rect 191658 568294 222198 568350
rect 222254 568294 222322 568350
rect 222378 568294 252918 568350
rect 252974 568294 253042 568350
rect 253098 568294 283638 568350
rect 283694 568294 283762 568350
rect 283818 568294 314358 568350
rect 314414 568294 314482 568350
rect 314538 568294 345078 568350
rect 345134 568294 345202 568350
rect 345258 568294 375798 568350
rect 375854 568294 375922 568350
rect 375978 568294 406518 568350
rect 406574 568294 406642 568350
rect 406698 568294 437238 568350
rect 437294 568294 437362 568350
rect 437418 568294 467958 568350
rect 468014 568294 468082 568350
rect 468138 568294 498678 568350
rect 498734 568294 498802 568350
rect 498858 568294 529398 568350
rect 529454 568294 529522 568350
rect 529578 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 37878 568226
rect 37934 568170 38002 568226
rect 38058 568170 68598 568226
rect 68654 568170 68722 568226
rect 68778 568170 99318 568226
rect 99374 568170 99442 568226
rect 99498 568170 130038 568226
rect 130094 568170 130162 568226
rect 130218 568170 160758 568226
rect 160814 568170 160882 568226
rect 160938 568170 191478 568226
rect 191534 568170 191602 568226
rect 191658 568170 222198 568226
rect 222254 568170 222322 568226
rect 222378 568170 252918 568226
rect 252974 568170 253042 568226
rect 253098 568170 283638 568226
rect 283694 568170 283762 568226
rect 283818 568170 314358 568226
rect 314414 568170 314482 568226
rect 314538 568170 345078 568226
rect 345134 568170 345202 568226
rect 345258 568170 375798 568226
rect 375854 568170 375922 568226
rect 375978 568170 406518 568226
rect 406574 568170 406642 568226
rect 406698 568170 437238 568226
rect 437294 568170 437362 568226
rect 437418 568170 467958 568226
rect 468014 568170 468082 568226
rect 468138 568170 498678 568226
rect 498734 568170 498802 568226
rect 498858 568170 529398 568226
rect 529454 568170 529522 568226
rect 529578 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 37878 568102
rect 37934 568046 38002 568102
rect 38058 568046 68598 568102
rect 68654 568046 68722 568102
rect 68778 568046 99318 568102
rect 99374 568046 99442 568102
rect 99498 568046 130038 568102
rect 130094 568046 130162 568102
rect 130218 568046 160758 568102
rect 160814 568046 160882 568102
rect 160938 568046 191478 568102
rect 191534 568046 191602 568102
rect 191658 568046 222198 568102
rect 222254 568046 222322 568102
rect 222378 568046 252918 568102
rect 252974 568046 253042 568102
rect 253098 568046 283638 568102
rect 283694 568046 283762 568102
rect 283818 568046 314358 568102
rect 314414 568046 314482 568102
rect 314538 568046 345078 568102
rect 345134 568046 345202 568102
rect 345258 568046 375798 568102
rect 375854 568046 375922 568102
rect 375978 568046 406518 568102
rect 406574 568046 406642 568102
rect 406698 568046 437238 568102
rect 437294 568046 437362 568102
rect 437418 568046 467958 568102
rect 468014 568046 468082 568102
rect 468138 568046 498678 568102
rect 498734 568046 498802 568102
rect 498858 568046 529398 568102
rect 529454 568046 529522 568102
rect 529578 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 37878 567978
rect 37934 567922 38002 567978
rect 38058 567922 68598 567978
rect 68654 567922 68722 567978
rect 68778 567922 99318 567978
rect 99374 567922 99442 567978
rect 99498 567922 130038 567978
rect 130094 567922 130162 567978
rect 130218 567922 160758 567978
rect 160814 567922 160882 567978
rect 160938 567922 191478 567978
rect 191534 567922 191602 567978
rect 191658 567922 222198 567978
rect 222254 567922 222322 567978
rect 222378 567922 252918 567978
rect 252974 567922 253042 567978
rect 253098 567922 283638 567978
rect 283694 567922 283762 567978
rect 283818 567922 314358 567978
rect 314414 567922 314482 567978
rect 314538 567922 345078 567978
rect 345134 567922 345202 567978
rect 345258 567922 375798 567978
rect 375854 567922 375922 567978
rect 375978 567922 406518 567978
rect 406574 567922 406642 567978
rect 406698 567922 437238 567978
rect 437294 567922 437362 567978
rect 437418 567922 467958 567978
rect 468014 567922 468082 567978
rect 468138 567922 498678 567978
rect 498734 567922 498802 567978
rect 498858 567922 529398 567978
rect 529454 567922 529522 567978
rect 529578 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 22518 562350
rect 22574 562294 22642 562350
rect 22698 562294 53238 562350
rect 53294 562294 53362 562350
rect 53418 562294 83958 562350
rect 84014 562294 84082 562350
rect 84138 562294 114678 562350
rect 114734 562294 114802 562350
rect 114858 562294 145398 562350
rect 145454 562294 145522 562350
rect 145578 562294 176118 562350
rect 176174 562294 176242 562350
rect 176298 562294 206838 562350
rect 206894 562294 206962 562350
rect 207018 562294 237558 562350
rect 237614 562294 237682 562350
rect 237738 562294 268278 562350
rect 268334 562294 268402 562350
rect 268458 562294 298998 562350
rect 299054 562294 299122 562350
rect 299178 562294 329718 562350
rect 329774 562294 329842 562350
rect 329898 562294 360438 562350
rect 360494 562294 360562 562350
rect 360618 562294 391158 562350
rect 391214 562294 391282 562350
rect 391338 562294 421878 562350
rect 421934 562294 422002 562350
rect 422058 562294 452598 562350
rect 452654 562294 452722 562350
rect 452778 562294 483318 562350
rect 483374 562294 483442 562350
rect 483498 562294 514038 562350
rect 514094 562294 514162 562350
rect 514218 562294 544758 562350
rect 544814 562294 544882 562350
rect 544938 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 22518 562226
rect 22574 562170 22642 562226
rect 22698 562170 53238 562226
rect 53294 562170 53362 562226
rect 53418 562170 83958 562226
rect 84014 562170 84082 562226
rect 84138 562170 114678 562226
rect 114734 562170 114802 562226
rect 114858 562170 145398 562226
rect 145454 562170 145522 562226
rect 145578 562170 176118 562226
rect 176174 562170 176242 562226
rect 176298 562170 206838 562226
rect 206894 562170 206962 562226
rect 207018 562170 237558 562226
rect 237614 562170 237682 562226
rect 237738 562170 268278 562226
rect 268334 562170 268402 562226
rect 268458 562170 298998 562226
rect 299054 562170 299122 562226
rect 299178 562170 329718 562226
rect 329774 562170 329842 562226
rect 329898 562170 360438 562226
rect 360494 562170 360562 562226
rect 360618 562170 391158 562226
rect 391214 562170 391282 562226
rect 391338 562170 421878 562226
rect 421934 562170 422002 562226
rect 422058 562170 452598 562226
rect 452654 562170 452722 562226
rect 452778 562170 483318 562226
rect 483374 562170 483442 562226
rect 483498 562170 514038 562226
rect 514094 562170 514162 562226
rect 514218 562170 544758 562226
rect 544814 562170 544882 562226
rect 544938 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 22518 562102
rect 22574 562046 22642 562102
rect 22698 562046 53238 562102
rect 53294 562046 53362 562102
rect 53418 562046 83958 562102
rect 84014 562046 84082 562102
rect 84138 562046 114678 562102
rect 114734 562046 114802 562102
rect 114858 562046 145398 562102
rect 145454 562046 145522 562102
rect 145578 562046 176118 562102
rect 176174 562046 176242 562102
rect 176298 562046 206838 562102
rect 206894 562046 206962 562102
rect 207018 562046 237558 562102
rect 237614 562046 237682 562102
rect 237738 562046 268278 562102
rect 268334 562046 268402 562102
rect 268458 562046 298998 562102
rect 299054 562046 299122 562102
rect 299178 562046 329718 562102
rect 329774 562046 329842 562102
rect 329898 562046 360438 562102
rect 360494 562046 360562 562102
rect 360618 562046 391158 562102
rect 391214 562046 391282 562102
rect 391338 562046 421878 562102
rect 421934 562046 422002 562102
rect 422058 562046 452598 562102
rect 452654 562046 452722 562102
rect 452778 562046 483318 562102
rect 483374 562046 483442 562102
rect 483498 562046 514038 562102
rect 514094 562046 514162 562102
rect 514218 562046 544758 562102
rect 544814 562046 544882 562102
rect 544938 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 22518 561978
rect 22574 561922 22642 561978
rect 22698 561922 53238 561978
rect 53294 561922 53362 561978
rect 53418 561922 83958 561978
rect 84014 561922 84082 561978
rect 84138 561922 114678 561978
rect 114734 561922 114802 561978
rect 114858 561922 145398 561978
rect 145454 561922 145522 561978
rect 145578 561922 176118 561978
rect 176174 561922 176242 561978
rect 176298 561922 206838 561978
rect 206894 561922 206962 561978
rect 207018 561922 237558 561978
rect 237614 561922 237682 561978
rect 237738 561922 268278 561978
rect 268334 561922 268402 561978
rect 268458 561922 298998 561978
rect 299054 561922 299122 561978
rect 299178 561922 329718 561978
rect 329774 561922 329842 561978
rect 329898 561922 360438 561978
rect 360494 561922 360562 561978
rect 360618 561922 391158 561978
rect 391214 561922 391282 561978
rect 391338 561922 421878 561978
rect 421934 561922 422002 561978
rect 422058 561922 452598 561978
rect 452654 561922 452722 561978
rect 452778 561922 483318 561978
rect 483374 561922 483442 561978
rect 483498 561922 514038 561978
rect 514094 561922 514162 561978
rect 514218 561922 544758 561978
rect 544814 561922 544882 561978
rect 544938 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 37878 550350
rect 37934 550294 38002 550350
rect 38058 550294 68598 550350
rect 68654 550294 68722 550350
rect 68778 550294 99318 550350
rect 99374 550294 99442 550350
rect 99498 550294 130038 550350
rect 130094 550294 130162 550350
rect 130218 550294 160758 550350
rect 160814 550294 160882 550350
rect 160938 550294 191478 550350
rect 191534 550294 191602 550350
rect 191658 550294 222198 550350
rect 222254 550294 222322 550350
rect 222378 550294 252918 550350
rect 252974 550294 253042 550350
rect 253098 550294 283638 550350
rect 283694 550294 283762 550350
rect 283818 550294 314358 550350
rect 314414 550294 314482 550350
rect 314538 550294 345078 550350
rect 345134 550294 345202 550350
rect 345258 550294 375798 550350
rect 375854 550294 375922 550350
rect 375978 550294 406518 550350
rect 406574 550294 406642 550350
rect 406698 550294 437238 550350
rect 437294 550294 437362 550350
rect 437418 550294 467958 550350
rect 468014 550294 468082 550350
rect 468138 550294 498678 550350
rect 498734 550294 498802 550350
rect 498858 550294 529398 550350
rect 529454 550294 529522 550350
rect 529578 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 37878 550226
rect 37934 550170 38002 550226
rect 38058 550170 68598 550226
rect 68654 550170 68722 550226
rect 68778 550170 99318 550226
rect 99374 550170 99442 550226
rect 99498 550170 130038 550226
rect 130094 550170 130162 550226
rect 130218 550170 160758 550226
rect 160814 550170 160882 550226
rect 160938 550170 191478 550226
rect 191534 550170 191602 550226
rect 191658 550170 222198 550226
rect 222254 550170 222322 550226
rect 222378 550170 252918 550226
rect 252974 550170 253042 550226
rect 253098 550170 283638 550226
rect 283694 550170 283762 550226
rect 283818 550170 314358 550226
rect 314414 550170 314482 550226
rect 314538 550170 345078 550226
rect 345134 550170 345202 550226
rect 345258 550170 375798 550226
rect 375854 550170 375922 550226
rect 375978 550170 406518 550226
rect 406574 550170 406642 550226
rect 406698 550170 437238 550226
rect 437294 550170 437362 550226
rect 437418 550170 467958 550226
rect 468014 550170 468082 550226
rect 468138 550170 498678 550226
rect 498734 550170 498802 550226
rect 498858 550170 529398 550226
rect 529454 550170 529522 550226
rect 529578 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 37878 550102
rect 37934 550046 38002 550102
rect 38058 550046 68598 550102
rect 68654 550046 68722 550102
rect 68778 550046 99318 550102
rect 99374 550046 99442 550102
rect 99498 550046 130038 550102
rect 130094 550046 130162 550102
rect 130218 550046 160758 550102
rect 160814 550046 160882 550102
rect 160938 550046 191478 550102
rect 191534 550046 191602 550102
rect 191658 550046 222198 550102
rect 222254 550046 222322 550102
rect 222378 550046 252918 550102
rect 252974 550046 253042 550102
rect 253098 550046 283638 550102
rect 283694 550046 283762 550102
rect 283818 550046 314358 550102
rect 314414 550046 314482 550102
rect 314538 550046 345078 550102
rect 345134 550046 345202 550102
rect 345258 550046 375798 550102
rect 375854 550046 375922 550102
rect 375978 550046 406518 550102
rect 406574 550046 406642 550102
rect 406698 550046 437238 550102
rect 437294 550046 437362 550102
rect 437418 550046 467958 550102
rect 468014 550046 468082 550102
rect 468138 550046 498678 550102
rect 498734 550046 498802 550102
rect 498858 550046 529398 550102
rect 529454 550046 529522 550102
rect 529578 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 37878 549978
rect 37934 549922 38002 549978
rect 38058 549922 68598 549978
rect 68654 549922 68722 549978
rect 68778 549922 99318 549978
rect 99374 549922 99442 549978
rect 99498 549922 130038 549978
rect 130094 549922 130162 549978
rect 130218 549922 160758 549978
rect 160814 549922 160882 549978
rect 160938 549922 191478 549978
rect 191534 549922 191602 549978
rect 191658 549922 222198 549978
rect 222254 549922 222322 549978
rect 222378 549922 252918 549978
rect 252974 549922 253042 549978
rect 253098 549922 283638 549978
rect 283694 549922 283762 549978
rect 283818 549922 314358 549978
rect 314414 549922 314482 549978
rect 314538 549922 345078 549978
rect 345134 549922 345202 549978
rect 345258 549922 375798 549978
rect 375854 549922 375922 549978
rect 375978 549922 406518 549978
rect 406574 549922 406642 549978
rect 406698 549922 437238 549978
rect 437294 549922 437362 549978
rect 437418 549922 467958 549978
rect 468014 549922 468082 549978
rect 468138 549922 498678 549978
rect 498734 549922 498802 549978
rect 498858 549922 529398 549978
rect 529454 549922 529522 549978
rect 529578 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 22518 544350
rect 22574 544294 22642 544350
rect 22698 544294 53238 544350
rect 53294 544294 53362 544350
rect 53418 544294 83958 544350
rect 84014 544294 84082 544350
rect 84138 544294 114678 544350
rect 114734 544294 114802 544350
rect 114858 544294 145398 544350
rect 145454 544294 145522 544350
rect 145578 544294 176118 544350
rect 176174 544294 176242 544350
rect 176298 544294 206838 544350
rect 206894 544294 206962 544350
rect 207018 544294 237558 544350
rect 237614 544294 237682 544350
rect 237738 544294 268278 544350
rect 268334 544294 268402 544350
rect 268458 544294 298998 544350
rect 299054 544294 299122 544350
rect 299178 544294 329718 544350
rect 329774 544294 329842 544350
rect 329898 544294 360438 544350
rect 360494 544294 360562 544350
rect 360618 544294 391158 544350
rect 391214 544294 391282 544350
rect 391338 544294 421878 544350
rect 421934 544294 422002 544350
rect 422058 544294 452598 544350
rect 452654 544294 452722 544350
rect 452778 544294 483318 544350
rect 483374 544294 483442 544350
rect 483498 544294 514038 544350
rect 514094 544294 514162 544350
rect 514218 544294 544758 544350
rect 544814 544294 544882 544350
rect 544938 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 22518 544226
rect 22574 544170 22642 544226
rect 22698 544170 53238 544226
rect 53294 544170 53362 544226
rect 53418 544170 83958 544226
rect 84014 544170 84082 544226
rect 84138 544170 114678 544226
rect 114734 544170 114802 544226
rect 114858 544170 145398 544226
rect 145454 544170 145522 544226
rect 145578 544170 176118 544226
rect 176174 544170 176242 544226
rect 176298 544170 206838 544226
rect 206894 544170 206962 544226
rect 207018 544170 237558 544226
rect 237614 544170 237682 544226
rect 237738 544170 268278 544226
rect 268334 544170 268402 544226
rect 268458 544170 298998 544226
rect 299054 544170 299122 544226
rect 299178 544170 329718 544226
rect 329774 544170 329842 544226
rect 329898 544170 360438 544226
rect 360494 544170 360562 544226
rect 360618 544170 391158 544226
rect 391214 544170 391282 544226
rect 391338 544170 421878 544226
rect 421934 544170 422002 544226
rect 422058 544170 452598 544226
rect 452654 544170 452722 544226
rect 452778 544170 483318 544226
rect 483374 544170 483442 544226
rect 483498 544170 514038 544226
rect 514094 544170 514162 544226
rect 514218 544170 544758 544226
rect 544814 544170 544882 544226
rect 544938 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 22518 544102
rect 22574 544046 22642 544102
rect 22698 544046 53238 544102
rect 53294 544046 53362 544102
rect 53418 544046 83958 544102
rect 84014 544046 84082 544102
rect 84138 544046 114678 544102
rect 114734 544046 114802 544102
rect 114858 544046 145398 544102
rect 145454 544046 145522 544102
rect 145578 544046 176118 544102
rect 176174 544046 176242 544102
rect 176298 544046 206838 544102
rect 206894 544046 206962 544102
rect 207018 544046 237558 544102
rect 237614 544046 237682 544102
rect 237738 544046 268278 544102
rect 268334 544046 268402 544102
rect 268458 544046 298998 544102
rect 299054 544046 299122 544102
rect 299178 544046 329718 544102
rect 329774 544046 329842 544102
rect 329898 544046 360438 544102
rect 360494 544046 360562 544102
rect 360618 544046 391158 544102
rect 391214 544046 391282 544102
rect 391338 544046 421878 544102
rect 421934 544046 422002 544102
rect 422058 544046 452598 544102
rect 452654 544046 452722 544102
rect 452778 544046 483318 544102
rect 483374 544046 483442 544102
rect 483498 544046 514038 544102
rect 514094 544046 514162 544102
rect 514218 544046 544758 544102
rect 544814 544046 544882 544102
rect 544938 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 22518 543978
rect 22574 543922 22642 543978
rect 22698 543922 53238 543978
rect 53294 543922 53362 543978
rect 53418 543922 83958 543978
rect 84014 543922 84082 543978
rect 84138 543922 114678 543978
rect 114734 543922 114802 543978
rect 114858 543922 145398 543978
rect 145454 543922 145522 543978
rect 145578 543922 176118 543978
rect 176174 543922 176242 543978
rect 176298 543922 206838 543978
rect 206894 543922 206962 543978
rect 207018 543922 237558 543978
rect 237614 543922 237682 543978
rect 237738 543922 268278 543978
rect 268334 543922 268402 543978
rect 268458 543922 298998 543978
rect 299054 543922 299122 543978
rect 299178 543922 329718 543978
rect 329774 543922 329842 543978
rect 329898 543922 360438 543978
rect 360494 543922 360562 543978
rect 360618 543922 391158 543978
rect 391214 543922 391282 543978
rect 391338 543922 421878 543978
rect 421934 543922 422002 543978
rect 422058 543922 452598 543978
rect 452654 543922 452722 543978
rect 452778 543922 483318 543978
rect 483374 543922 483442 543978
rect 483498 543922 514038 543978
rect 514094 543922 514162 543978
rect 514218 543922 544758 543978
rect 544814 543922 544882 543978
rect 544938 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 37878 532350
rect 37934 532294 38002 532350
rect 38058 532294 68598 532350
rect 68654 532294 68722 532350
rect 68778 532294 99318 532350
rect 99374 532294 99442 532350
rect 99498 532294 130038 532350
rect 130094 532294 130162 532350
rect 130218 532294 160758 532350
rect 160814 532294 160882 532350
rect 160938 532294 191478 532350
rect 191534 532294 191602 532350
rect 191658 532294 222198 532350
rect 222254 532294 222322 532350
rect 222378 532294 252918 532350
rect 252974 532294 253042 532350
rect 253098 532294 283638 532350
rect 283694 532294 283762 532350
rect 283818 532294 314358 532350
rect 314414 532294 314482 532350
rect 314538 532294 345078 532350
rect 345134 532294 345202 532350
rect 345258 532294 375798 532350
rect 375854 532294 375922 532350
rect 375978 532294 406518 532350
rect 406574 532294 406642 532350
rect 406698 532294 437238 532350
rect 437294 532294 437362 532350
rect 437418 532294 467958 532350
rect 468014 532294 468082 532350
rect 468138 532294 498678 532350
rect 498734 532294 498802 532350
rect 498858 532294 529398 532350
rect 529454 532294 529522 532350
rect 529578 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 37878 532226
rect 37934 532170 38002 532226
rect 38058 532170 68598 532226
rect 68654 532170 68722 532226
rect 68778 532170 99318 532226
rect 99374 532170 99442 532226
rect 99498 532170 130038 532226
rect 130094 532170 130162 532226
rect 130218 532170 160758 532226
rect 160814 532170 160882 532226
rect 160938 532170 191478 532226
rect 191534 532170 191602 532226
rect 191658 532170 222198 532226
rect 222254 532170 222322 532226
rect 222378 532170 252918 532226
rect 252974 532170 253042 532226
rect 253098 532170 283638 532226
rect 283694 532170 283762 532226
rect 283818 532170 314358 532226
rect 314414 532170 314482 532226
rect 314538 532170 345078 532226
rect 345134 532170 345202 532226
rect 345258 532170 375798 532226
rect 375854 532170 375922 532226
rect 375978 532170 406518 532226
rect 406574 532170 406642 532226
rect 406698 532170 437238 532226
rect 437294 532170 437362 532226
rect 437418 532170 467958 532226
rect 468014 532170 468082 532226
rect 468138 532170 498678 532226
rect 498734 532170 498802 532226
rect 498858 532170 529398 532226
rect 529454 532170 529522 532226
rect 529578 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 37878 532102
rect 37934 532046 38002 532102
rect 38058 532046 68598 532102
rect 68654 532046 68722 532102
rect 68778 532046 99318 532102
rect 99374 532046 99442 532102
rect 99498 532046 130038 532102
rect 130094 532046 130162 532102
rect 130218 532046 160758 532102
rect 160814 532046 160882 532102
rect 160938 532046 191478 532102
rect 191534 532046 191602 532102
rect 191658 532046 222198 532102
rect 222254 532046 222322 532102
rect 222378 532046 252918 532102
rect 252974 532046 253042 532102
rect 253098 532046 283638 532102
rect 283694 532046 283762 532102
rect 283818 532046 314358 532102
rect 314414 532046 314482 532102
rect 314538 532046 345078 532102
rect 345134 532046 345202 532102
rect 345258 532046 375798 532102
rect 375854 532046 375922 532102
rect 375978 532046 406518 532102
rect 406574 532046 406642 532102
rect 406698 532046 437238 532102
rect 437294 532046 437362 532102
rect 437418 532046 467958 532102
rect 468014 532046 468082 532102
rect 468138 532046 498678 532102
rect 498734 532046 498802 532102
rect 498858 532046 529398 532102
rect 529454 532046 529522 532102
rect 529578 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 37878 531978
rect 37934 531922 38002 531978
rect 38058 531922 68598 531978
rect 68654 531922 68722 531978
rect 68778 531922 99318 531978
rect 99374 531922 99442 531978
rect 99498 531922 130038 531978
rect 130094 531922 130162 531978
rect 130218 531922 160758 531978
rect 160814 531922 160882 531978
rect 160938 531922 191478 531978
rect 191534 531922 191602 531978
rect 191658 531922 222198 531978
rect 222254 531922 222322 531978
rect 222378 531922 252918 531978
rect 252974 531922 253042 531978
rect 253098 531922 283638 531978
rect 283694 531922 283762 531978
rect 283818 531922 314358 531978
rect 314414 531922 314482 531978
rect 314538 531922 345078 531978
rect 345134 531922 345202 531978
rect 345258 531922 375798 531978
rect 375854 531922 375922 531978
rect 375978 531922 406518 531978
rect 406574 531922 406642 531978
rect 406698 531922 437238 531978
rect 437294 531922 437362 531978
rect 437418 531922 467958 531978
rect 468014 531922 468082 531978
rect 468138 531922 498678 531978
rect 498734 531922 498802 531978
rect 498858 531922 529398 531978
rect 529454 531922 529522 531978
rect 529578 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 22518 526350
rect 22574 526294 22642 526350
rect 22698 526294 53238 526350
rect 53294 526294 53362 526350
rect 53418 526294 83958 526350
rect 84014 526294 84082 526350
rect 84138 526294 114678 526350
rect 114734 526294 114802 526350
rect 114858 526294 145398 526350
rect 145454 526294 145522 526350
rect 145578 526294 176118 526350
rect 176174 526294 176242 526350
rect 176298 526294 206838 526350
rect 206894 526294 206962 526350
rect 207018 526294 237558 526350
rect 237614 526294 237682 526350
rect 237738 526294 268278 526350
rect 268334 526294 268402 526350
rect 268458 526294 298998 526350
rect 299054 526294 299122 526350
rect 299178 526294 329718 526350
rect 329774 526294 329842 526350
rect 329898 526294 360438 526350
rect 360494 526294 360562 526350
rect 360618 526294 391158 526350
rect 391214 526294 391282 526350
rect 391338 526294 421878 526350
rect 421934 526294 422002 526350
rect 422058 526294 452598 526350
rect 452654 526294 452722 526350
rect 452778 526294 483318 526350
rect 483374 526294 483442 526350
rect 483498 526294 514038 526350
rect 514094 526294 514162 526350
rect 514218 526294 544758 526350
rect 544814 526294 544882 526350
rect 544938 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 22518 526226
rect 22574 526170 22642 526226
rect 22698 526170 53238 526226
rect 53294 526170 53362 526226
rect 53418 526170 83958 526226
rect 84014 526170 84082 526226
rect 84138 526170 114678 526226
rect 114734 526170 114802 526226
rect 114858 526170 145398 526226
rect 145454 526170 145522 526226
rect 145578 526170 176118 526226
rect 176174 526170 176242 526226
rect 176298 526170 206838 526226
rect 206894 526170 206962 526226
rect 207018 526170 237558 526226
rect 237614 526170 237682 526226
rect 237738 526170 268278 526226
rect 268334 526170 268402 526226
rect 268458 526170 298998 526226
rect 299054 526170 299122 526226
rect 299178 526170 329718 526226
rect 329774 526170 329842 526226
rect 329898 526170 360438 526226
rect 360494 526170 360562 526226
rect 360618 526170 391158 526226
rect 391214 526170 391282 526226
rect 391338 526170 421878 526226
rect 421934 526170 422002 526226
rect 422058 526170 452598 526226
rect 452654 526170 452722 526226
rect 452778 526170 483318 526226
rect 483374 526170 483442 526226
rect 483498 526170 514038 526226
rect 514094 526170 514162 526226
rect 514218 526170 544758 526226
rect 544814 526170 544882 526226
rect 544938 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 22518 526102
rect 22574 526046 22642 526102
rect 22698 526046 53238 526102
rect 53294 526046 53362 526102
rect 53418 526046 83958 526102
rect 84014 526046 84082 526102
rect 84138 526046 114678 526102
rect 114734 526046 114802 526102
rect 114858 526046 145398 526102
rect 145454 526046 145522 526102
rect 145578 526046 176118 526102
rect 176174 526046 176242 526102
rect 176298 526046 206838 526102
rect 206894 526046 206962 526102
rect 207018 526046 237558 526102
rect 237614 526046 237682 526102
rect 237738 526046 268278 526102
rect 268334 526046 268402 526102
rect 268458 526046 298998 526102
rect 299054 526046 299122 526102
rect 299178 526046 329718 526102
rect 329774 526046 329842 526102
rect 329898 526046 360438 526102
rect 360494 526046 360562 526102
rect 360618 526046 391158 526102
rect 391214 526046 391282 526102
rect 391338 526046 421878 526102
rect 421934 526046 422002 526102
rect 422058 526046 452598 526102
rect 452654 526046 452722 526102
rect 452778 526046 483318 526102
rect 483374 526046 483442 526102
rect 483498 526046 514038 526102
rect 514094 526046 514162 526102
rect 514218 526046 544758 526102
rect 544814 526046 544882 526102
rect 544938 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 22518 525978
rect 22574 525922 22642 525978
rect 22698 525922 53238 525978
rect 53294 525922 53362 525978
rect 53418 525922 83958 525978
rect 84014 525922 84082 525978
rect 84138 525922 114678 525978
rect 114734 525922 114802 525978
rect 114858 525922 145398 525978
rect 145454 525922 145522 525978
rect 145578 525922 176118 525978
rect 176174 525922 176242 525978
rect 176298 525922 206838 525978
rect 206894 525922 206962 525978
rect 207018 525922 237558 525978
rect 237614 525922 237682 525978
rect 237738 525922 268278 525978
rect 268334 525922 268402 525978
rect 268458 525922 298998 525978
rect 299054 525922 299122 525978
rect 299178 525922 329718 525978
rect 329774 525922 329842 525978
rect 329898 525922 360438 525978
rect 360494 525922 360562 525978
rect 360618 525922 391158 525978
rect 391214 525922 391282 525978
rect 391338 525922 421878 525978
rect 421934 525922 422002 525978
rect 422058 525922 452598 525978
rect 452654 525922 452722 525978
rect 452778 525922 483318 525978
rect 483374 525922 483442 525978
rect 483498 525922 514038 525978
rect 514094 525922 514162 525978
rect 514218 525922 544758 525978
rect 544814 525922 544882 525978
rect 544938 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 37878 514350
rect 37934 514294 38002 514350
rect 38058 514294 68598 514350
rect 68654 514294 68722 514350
rect 68778 514294 99318 514350
rect 99374 514294 99442 514350
rect 99498 514294 130038 514350
rect 130094 514294 130162 514350
rect 130218 514294 160758 514350
rect 160814 514294 160882 514350
rect 160938 514294 191478 514350
rect 191534 514294 191602 514350
rect 191658 514294 222198 514350
rect 222254 514294 222322 514350
rect 222378 514294 252918 514350
rect 252974 514294 253042 514350
rect 253098 514294 283638 514350
rect 283694 514294 283762 514350
rect 283818 514294 314358 514350
rect 314414 514294 314482 514350
rect 314538 514294 345078 514350
rect 345134 514294 345202 514350
rect 345258 514294 375798 514350
rect 375854 514294 375922 514350
rect 375978 514294 406518 514350
rect 406574 514294 406642 514350
rect 406698 514294 437238 514350
rect 437294 514294 437362 514350
rect 437418 514294 467958 514350
rect 468014 514294 468082 514350
rect 468138 514294 498678 514350
rect 498734 514294 498802 514350
rect 498858 514294 529398 514350
rect 529454 514294 529522 514350
rect 529578 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 37878 514226
rect 37934 514170 38002 514226
rect 38058 514170 68598 514226
rect 68654 514170 68722 514226
rect 68778 514170 99318 514226
rect 99374 514170 99442 514226
rect 99498 514170 130038 514226
rect 130094 514170 130162 514226
rect 130218 514170 160758 514226
rect 160814 514170 160882 514226
rect 160938 514170 191478 514226
rect 191534 514170 191602 514226
rect 191658 514170 222198 514226
rect 222254 514170 222322 514226
rect 222378 514170 252918 514226
rect 252974 514170 253042 514226
rect 253098 514170 283638 514226
rect 283694 514170 283762 514226
rect 283818 514170 314358 514226
rect 314414 514170 314482 514226
rect 314538 514170 345078 514226
rect 345134 514170 345202 514226
rect 345258 514170 375798 514226
rect 375854 514170 375922 514226
rect 375978 514170 406518 514226
rect 406574 514170 406642 514226
rect 406698 514170 437238 514226
rect 437294 514170 437362 514226
rect 437418 514170 467958 514226
rect 468014 514170 468082 514226
rect 468138 514170 498678 514226
rect 498734 514170 498802 514226
rect 498858 514170 529398 514226
rect 529454 514170 529522 514226
rect 529578 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 37878 514102
rect 37934 514046 38002 514102
rect 38058 514046 68598 514102
rect 68654 514046 68722 514102
rect 68778 514046 99318 514102
rect 99374 514046 99442 514102
rect 99498 514046 130038 514102
rect 130094 514046 130162 514102
rect 130218 514046 160758 514102
rect 160814 514046 160882 514102
rect 160938 514046 191478 514102
rect 191534 514046 191602 514102
rect 191658 514046 222198 514102
rect 222254 514046 222322 514102
rect 222378 514046 252918 514102
rect 252974 514046 253042 514102
rect 253098 514046 283638 514102
rect 283694 514046 283762 514102
rect 283818 514046 314358 514102
rect 314414 514046 314482 514102
rect 314538 514046 345078 514102
rect 345134 514046 345202 514102
rect 345258 514046 375798 514102
rect 375854 514046 375922 514102
rect 375978 514046 406518 514102
rect 406574 514046 406642 514102
rect 406698 514046 437238 514102
rect 437294 514046 437362 514102
rect 437418 514046 467958 514102
rect 468014 514046 468082 514102
rect 468138 514046 498678 514102
rect 498734 514046 498802 514102
rect 498858 514046 529398 514102
rect 529454 514046 529522 514102
rect 529578 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 37878 513978
rect 37934 513922 38002 513978
rect 38058 513922 68598 513978
rect 68654 513922 68722 513978
rect 68778 513922 99318 513978
rect 99374 513922 99442 513978
rect 99498 513922 130038 513978
rect 130094 513922 130162 513978
rect 130218 513922 160758 513978
rect 160814 513922 160882 513978
rect 160938 513922 191478 513978
rect 191534 513922 191602 513978
rect 191658 513922 222198 513978
rect 222254 513922 222322 513978
rect 222378 513922 252918 513978
rect 252974 513922 253042 513978
rect 253098 513922 283638 513978
rect 283694 513922 283762 513978
rect 283818 513922 314358 513978
rect 314414 513922 314482 513978
rect 314538 513922 345078 513978
rect 345134 513922 345202 513978
rect 345258 513922 375798 513978
rect 375854 513922 375922 513978
rect 375978 513922 406518 513978
rect 406574 513922 406642 513978
rect 406698 513922 437238 513978
rect 437294 513922 437362 513978
rect 437418 513922 467958 513978
rect 468014 513922 468082 513978
rect 468138 513922 498678 513978
rect 498734 513922 498802 513978
rect 498858 513922 529398 513978
rect 529454 513922 529522 513978
rect 529578 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 22518 508350
rect 22574 508294 22642 508350
rect 22698 508294 53238 508350
rect 53294 508294 53362 508350
rect 53418 508294 83958 508350
rect 84014 508294 84082 508350
rect 84138 508294 114678 508350
rect 114734 508294 114802 508350
rect 114858 508294 145398 508350
rect 145454 508294 145522 508350
rect 145578 508294 176118 508350
rect 176174 508294 176242 508350
rect 176298 508294 206838 508350
rect 206894 508294 206962 508350
rect 207018 508294 237558 508350
rect 237614 508294 237682 508350
rect 237738 508294 268278 508350
rect 268334 508294 268402 508350
rect 268458 508294 298998 508350
rect 299054 508294 299122 508350
rect 299178 508294 329718 508350
rect 329774 508294 329842 508350
rect 329898 508294 360438 508350
rect 360494 508294 360562 508350
rect 360618 508294 391158 508350
rect 391214 508294 391282 508350
rect 391338 508294 421878 508350
rect 421934 508294 422002 508350
rect 422058 508294 452598 508350
rect 452654 508294 452722 508350
rect 452778 508294 483318 508350
rect 483374 508294 483442 508350
rect 483498 508294 514038 508350
rect 514094 508294 514162 508350
rect 514218 508294 544758 508350
rect 544814 508294 544882 508350
rect 544938 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 22518 508226
rect 22574 508170 22642 508226
rect 22698 508170 53238 508226
rect 53294 508170 53362 508226
rect 53418 508170 83958 508226
rect 84014 508170 84082 508226
rect 84138 508170 114678 508226
rect 114734 508170 114802 508226
rect 114858 508170 145398 508226
rect 145454 508170 145522 508226
rect 145578 508170 176118 508226
rect 176174 508170 176242 508226
rect 176298 508170 206838 508226
rect 206894 508170 206962 508226
rect 207018 508170 237558 508226
rect 237614 508170 237682 508226
rect 237738 508170 268278 508226
rect 268334 508170 268402 508226
rect 268458 508170 298998 508226
rect 299054 508170 299122 508226
rect 299178 508170 329718 508226
rect 329774 508170 329842 508226
rect 329898 508170 360438 508226
rect 360494 508170 360562 508226
rect 360618 508170 391158 508226
rect 391214 508170 391282 508226
rect 391338 508170 421878 508226
rect 421934 508170 422002 508226
rect 422058 508170 452598 508226
rect 452654 508170 452722 508226
rect 452778 508170 483318 508226
rect 483374 508170 483442 508226
rect 483498 508170 514038 508226
rect 514094 508170 514162 508226
rect 514218 508170 544758 508226
rect 544814 508170 544882 508226
rect 544938 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 22518 508102
rect 22574 508046 22642 508102
rect 22698 508046 53238 508102
rect 53294 508046 53362 508102
rect 53418 508046 83958 508102
rect 84014 508046 84082 508102
rect 84138 508046 114678 508102
rect 114734 508046 114802 508102
rect 114858 508046 145398 508102
rect 145454 508046 145522 508102
rect 145578 508046 176118 508102
rect 176174 508046 176242 508102
rect 176298 508046 206838 508102
rect 206894 508046 206962 508102
rect 207018 508046 237558 508102
rect 237614 508046 237682 508102
rect 237738 508046 268278 508102
rect 268334 508046 268402 508102
rect 268458 508046 298998 508102
rect 299054 508046 299122 508102
rect 299178 508046 329718 508102
rect 329774 508046 329842 508102
rect 329898 508046 360438 508102
rect 360494 508046 360562 508102
rect 360618 508046 391158 508102
rect 391214 508046 391282 508102
rect 391338 508046 421878 508102
rect 421934 508046 422002 508102
rect 422058 508046 452598 508102
rect 452654 508046 452722 508102
rect 452778 508046 483318 508102
rect 483374 508046 483442 508102
rect 483498 508046 514038 508102
rect 514094 508046 514162 508102
rect 514218 508046 544758 508102
rect 544814 508046 544882 508102
rect 544938 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 22518 507978
rect 22574 507922 22642 507978
rect 22698 507922 53238 507978
rect 53294 507922 53362 507978
rect 53418 507922 83958 507978
rect 84014 507922 84082 507978
rect 84138 507922 114678 507978
rect 114734 507922 114802 507978
rect 114858 507922 145398 507978
rect 145454 507922 145522 507978
rect 145578 507922 176118 507978
rect 176174 507922 176242 507978
rect 176298 507922 206838 507978
rect 206894 507922 206962 507978
rect 207018 507922 237558 507978
rect 237614 507922 237682 507978
rect 237738 507922 268278 507978
rect 268334 507922 268402 507978
rect 268458 507922 298998 507978
rect 299054 507922 299122 507978
rect 299178 507922 329718 507978
rect 329774 507922 329842 507978
rect 329898 507922 360438 507978
rect 360494 507922 360562 507978
rect 360618 507922 391158 507978
rect 391214 507922 391282 507978
rect 391338 507922 421878 507978
rect 421934 507922 422002 507978
rect 422058 507922 452598 507978
rect 452654 507922 452722 507978
rect 452778 507922 483318 507978
rect 483374 507922 483442 507978
rect 483498 507922 514038 507978
rect 514094 507922 514162 507978
rect 514218 507922 544758 507978
rect 544814 507922 544882 507978
rect 544938 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 37878 496350
rect 37934 496294 38002 496350
rect 38058 496294 68598 496350
rect 68654 496294 68722 496350
rect 68778 496294 99318 496350
rect 99374 496294 99442 496350
rect 99498 496294 130038 496350
rect 130094 496294 130162 496350
rect 130218 496294 160758 496350
rect 160814 496294 160882 496350
rect 160938 496294 191478 496350
rect 191534 496294 191602 496350
rect 191658 496294 222198 496350
rect 222254 496294 222322 496350
rect 222378 496294 252918 496350
rect 252974 496294 253042 496350
rect 253098 496294 283638 496350
rect 283694 496294 283762 496350
rect 283818 496294 314358 496350
rect 314414 496294 314482 496350
rect 314538 496294 345078 496350
rect 345134 496294 345202 496350
rect 345258 496294 375798 496350
rect 375854 496294 375922 496350
rect 375978 496294 406518 496350
rect 406574 496294 406642 496350
rect 406698 496294 437238 496350
rect 437294 496294 437362 496350
rect 437418 496294 467958 496350
rect 468014 496294 468082 496350
rect 468138 496294 498678 496350
rect 498734 496294 498802 496350
rect 498858 496294 529398 496350
rect 529454 496294 529522 496350
rect 529578 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 37878 496226
rect 37934 496170 38002 496226
rect 38058 496170 68598 496226
rect 68654 496170 68722 496226
rect 68778 496170 99318 496226
rect 99374 496170 99442 496226
rect 99498 496170 130038 496226
rect 130094 496170 130162 496226
rect 130218 496170 160758 496226
rect 160814 496170 160882 496226
rect 160938 496170 191478 496226
rect 191534 496170 191602 496226
rect 191658 496170 222198 496226
rect 222254 496170 222322 496226
rect 222378 496170 252918 496226
rect 252974 496170 253042 496226
rect 253098 496170 283638 496226
rect 283694 496170 283762 496226
rect 283818 496170 314358 496226
rect 314414 496170 314482 496226
rect 314538 496170 345078 496226
rect 345134 496170 345202 496226
rect 345258 496170 375798 496226
rect 375854 496170 375922 496226
rect 375978 496170 406518 496226
rect 406574 496170 406642 496226
rect 406698 496170 437238 496226
rect 437294 496170 437362 496226
rect 437418 496170 467958 496226
rect 468014 496170 468082 496226
rect 468138 496170 498678 496226
rect 498734 496170 498802 496226
rect 498858 496170 529398 496226
rect 529454 496170 529522 496226
rect 529578 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 37878 496102
rect 37934 496046 38002 496102
rect 38058 496046 68598 496102
rect 68654 496046 68722 496102
rect 68778 496046 99318 496102
rect 99374 496046 99442 496102
rect 99498 496046 130038 496102
rect 130094 496046 130162 496102
rect 130218 496046 160758 496102
rect 160814 496046 160882 496102
rect 160938 496046 191478 496102
rect 191534 496046 191602 496102
rect 191658 496046 222198 496102
rect 222254 496046 222322 496102
rect 222378 496046 252918 496102
rect 252974 496046 253042 496102
rect 253098 496046 283638 496102
rect 283694 496046 283762 496102
rect 283818 496046 314358 496102
rect 314414 496046 314482 496102
rect 314538 496046 345078 496102
rect 345134 496046 345202 496102
rect 345258 496046 375798 496102
rect 375854 496046 375922 496102
rect 375978 496046 406518 496102
rect 406574 496046 406642 496102
rect 406698 496046 437238 496102
rect 437294 496046 437362 496102
rect 437418 496046 467958 496102
rect 468014 496046 468082 496102
rect 468138 496046 498678 496102
rect 498734 496046 498802 496102
rect 498858 496046 529398 496102
rect 529454 496046 529522 496102
rect 529578 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 37878 495978
rect 37934 495922 38002 495978
rect 38058 495922 68598 495978
rect 68654 495922 68722 495978
rect 68778 495922 99318 495978
rect 99374 495922 99442 495978
rect 99498 495922 130038 495978
rect 130094 495922 130162 495978
rect 130218 495922 160758 495978
rect 160814 495922 160882 495978
rect 160938 495922 191478 495978
rect 191534 495922 191602 495978
rect 191658 495922 222198 495978
rect 222254 495922 222322 495978
rect 222378 495922 252918 495978
rect 252974 495922 253042 495978
rect 253098 495922 283638 495978
rect 283694 495922 283762 495978
rect 283818 495922 314358 495978
rect 314414 495922 314482 495978
rect 314538 495922 345078 495978
rect 345134 495922 345202 495978
rect 345258 495922 375798 495978
rect 375854 495922 375922 495978
rect 375978 495922 406518 495978
rect 406574 495922 406642 495978
rect 406698 495922 437238 495978
rect 437294 495922 437362 495978
rect 437418 495922 467958 495978
rect 468014 495922 468082 495978
rect 468138 495922 498678 495978
rect 498734 495922 498802 495978
rect 498858 495922 529398 495978
rect 529454 495922 529522 495978
rect 529578 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 22518 490350
rect 22574 490294 22642 490350
rect 22698 490294 53238 490350
rect 53294 490294 53362 490350
rect 53418 490294 83958 490350
rect 84014 490294 84082 490350
rect 84138 490294 114678 490350
rect 114734 490294 114802 490350
rect 114858 490294 145398 490350
rect 145454 490294 145522 490350
rect 145578 490294 176118 490350
rect 176174 490294 176242 490350
rect 176298 490294 206838 490350
rect 206894 490294 206962 490350
rect 207018 490294 237558 490350
rect 237614 490294 237682 490350
rect 237738 490294 268278 490350
rect 268334 490294 268402 490350
rect 268458 490294 298998 490350
rect 299054 490294 299122 490350
rect 299178 490294 329718 490350
rect 329774 490294 329842 490350
rect 329898 490294 360438 490350
rect 360494 490294 360562 490350
rect 360618 490294 391158 490350
rect 391214 490294 391282 490350
rect 391338 490294 421878 490350
rect 421934 490294 422002 490350
rect 422058 490294 452598 490350
rect 452654 490294 452722 490350
rect 452778 490294 483318 490350
rect 483374 490294 483442 490350
rect 483498 490294 514038 490350
rect 514094 490294 514162 490350
rect 514218 490294 544758 490350
rect 544814 490294 544882 490350
rect 544938 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 22518 490226
rect 22574 490170 22642 490226
rect 22698 490170 53238 490226
rect 53294 490170 53362 490226
rect 53418 490170 83958 490226
rect 84014 490170 84082 490226
rect 84138 490170 114678 490226
rect 114734 490170 114802 490226
rect 114858 490170 145398 490226
rect 145454 490170 145522 490226
rect 145578 490170 176118 490226
rect 176174 490170 176242 490226
rect 176298 490170 206838 490226
rect 206894 490170 206962 490226
rect 207018 490170 237558 490226
rect 237614 490170 237682 490226
rect 237738 490170 268278 490226
rect 268334 490170 268402 490226
rect 268458 490170 298998 490226
rect 299054 490170 299122 490226
rect 299178 490170 329718 490226
rect 329774 490170 329842 490226
rect 329898 490170 360438 490226
rect 360494 490170 360562 490226
rect 360618 490170 391158 490226
rect 391214 490170 391282 490226
rect 391338 490170 421878 490226
rect 421934 490170 422002 490226
rect 422058 490170 452598 490226
rect 452654 490170 452722 490226
rect 452778 490170 483318 490226
rect 483374 490170 483442 490226
rect 483498 490170 514038 490226
rect 514094 490170 514162 490226
rect 514218 490170 544758 490226
rect 544814 490170 544882 490226
rect 544938 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 22518 490102
rect 22574 490046 22642 490102
rect 22698 490046 53238 490102
rect 53294 490046 53362 490102
rect 53418 490046 83958 490102
rect 84014 490046 84082 490102
rect 84138 490046 114678 490102
rect 114734 490046 114802 490102
rect 114858 490046 145398 490102
rect 145454 490046 145522 490102
rect 145578 490046 176118 490102
rect 176174 490046 176242 490102
rect 176298 490046 206838 490102
rect 206894 490046 206962 490102
rect 207018 490046 237558 490102
rect 237614 490046 237682 490102
rect 237738 490046 268278 490102
rect 268334 490046 268402 490102
rect 268458 490046 298998 490102
rect 299054 490046 299122 490102
rect 299178 490046 329718 490102
rect 329774 490046 329842 490102
rect 329898 490046 360438 490102
rect 360494 490046 360562 490102
rect 360618 490046 391158 490102
rect 391214 490046 391282 490102
rect 391338 490046 421878 490102
rect 421934 490046 422002 490102
rect 422058 490046 452598 490102
rect 452654 490046 452722 490102
rect 452778 490046 483318 490102
rect 483374 490046 483442 490102
rect 483498 490046 514038 490102
rect 514094 490046 514162 490102
rect 514218 490046 544758 490102
rect 544814 490046 544882 490102
rect 544938 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 22518 489978
rect 22574 489922 22642 489978
rect 22698 489922 53238 489978
rect 53294 489922 53362 489978
rect 53418 489922 83958 489978
rect 84014 489922 84082 489978
rect 84138 489922 114678 489978
rect 114734 489922 114802 489978
rect 114858 489922 145398 489978
rect 145454 489922 145522 489978
rect 145578 489922 176118 489978
rect 176174 489922 176242 489978
rect 176298 489922 206838 489978
rect 206894 489922 206962 489978
rect 207018 489922 237558 489978
rect 237614 489922 237682 489978
rect 237738 489922 268278 489978
rect 268334 489922 268402 489978
rect 268458 489922 298998 489978
rect 299054 489922 299122 489978
rect 299178 489922 329718 489978
rect 329774 489922 329842 489978
rect 329898 489922 360438 489978
rect 360494 489922 360562 489978
rect 360618 489922 391158 489978
rect 391214 489922 391282 489978
rect 391338 489922 421878 489978
rect 421934 489922 422002 489978
rect 422058 489922 452598 489978
rect 452654 489922 452722 489978
rect 452778 489922 483318 489978
rect 483374 489922 483442 489978
rect 483498 489922 514038 489978
rect 514094 489922 514162 489978
rect 514218 489922 544758 489978
rect 544814 489922 544882 489978
rect 544938 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 37878 478350
rect 37934 478294 38002 478350
rect 38058 478294 68598 478350
rect 68654 478294 68722 478350
rect 68778 478294 99318 478350
rect 99374 478294 99442 478350
rect 99498 478294 130038 478350
rect 130094 478294 130162 478350
rect 130218 478294 160758 478350
rect 160814 478294 160882 478350
rect 160938 478294 191478 478350
rect 191534 478294 191602 478350
rect 191658 478294 222198 478350
rect 222254 478294 222322 478350
rect 222378 478294 252918 478350
rect 252974 478294 253042 478350
rect 253098 478294 283638 478350
rect 283694 478294 283762 478350
rect 283818 478294 314358 478350
rect 314414 478294 314482 478350
rect 314538 478294 345078 478350
rect 345134 478294 345202 478350
rect 345258 478294 375798 478350
rect 375854 478294 375922 478350
rect 375978 478294 406518 478350
rect 406574 478294 406642 478350
rect 406698 478294 437238 478350
rect 437294 478294 437362 478350
rect 437418 478294 467958 478350
rect 468014 478294 468082 478350
rect 468138 478294 498678 478350
rect 498734 478294 498802 478350
rect 498858 478294 529398 478350
rect 529454 478294 529522 478350
rect 529578 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 37878 478226
rect 37934 478170 38002 478226
rect 38058 478170 68598 478226
rect 68654 478170 68722 478226
rect 68778 478170 99318 478226
rect 99374 478170 99442 478226
rect 99498 478170 130038 478226
rect 130094 478170 130162 478226
rect 130218 478170 160758 478226
rect 160814 478170 160882 478226
rect 160938 478170 191478 478226
rect 191534 478170 191602 478226
rect 191658 478170 222198 478226
rect 222254 478170 222322 478226
rect 222378 478170 252918 478226
rect 252974 478170 253042 478226
rect 253098 478170 283638 478226
rect 283694 478170 283762 478226
rect 283818 478170 314358 478226
rect 314414 478170 314482 478226
rect 314538 478170 345078 478226
rect 345134 478170 345202 478226
rect 345258 478170 375798 478226
rect 375854 478170 375922 478226
rect 375978 478170 406518 478226
rect 406574 478170 406642 478226
rect 406698 478170 437238 478226
rect 437294 478170 437362 478226
rect 437418 478170 467958 478226
rect 468014 478170 468082 478226
rect 468138 478170 498678 478226
rect 498734 478170 498802 478226
rect 498858 478170 529398 478226
rect 529454 478170 529522 478226
rect 529578 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 37878 478102
rect 37934 478046 38002 478102
rect 38058 478046 68598 478102
rect 68654 478046 68722 478102
rect 68778 478046 99318 478102
rect 99374 478046 99442 478102
rect 99498 478046 130038 478102
rect 130094 478046 130162 478102
rect 130218 478046 160758 478102
rect 160814 478046 160882 478102
rect 160938 478046 191478 478102
rect 191534 478046 191602 478102
rect 191658 478046 222198 478102
rect 222254 478046 222322 478102
rect 222378 478046 252918 478102
rect 252974 478046 253042 478102
rect 253098 478046 283638 478102
rect 283694 478046 283762 478102
rect 283818 478046 314358 478102
rect 314414 478046 314482 478102
rect 314538 478046 345078 478102
rect 345134 478046 345202 478102
rect 345258 478046 375798 478102
rect 375854 478046 375922 478102
rect 375978 478046 406518 478102
rect 406574 478046 406642 478102
rect 406698 478046 437238 478102
rect 437294 478046 437362 478102
rect 437418 478046 467958 478102
rect 468014 478046 468082 478102
rect 468138 478046 498678 478102
rect 498734 478046 498802 478102
rect 498858 478046 529398 478102
rect 529454 478046 529522 478102
rect 529578 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 37878 477978
rect 37934 477922 38002 477978
rect 38058 477922 68598 477978
rect 68654 477922 68722 477978
rect 68778 477922 99318 477978
rect 99374 477922 99442 477978
rect 99498 477922 130038 477978
rect 130094 477922 130162 477978
rect 130218 477922 160758 477978
rect 160814 477922 160882 477978
rect 160938 477922 191478 477978
rect 191534 477922 191602 477978
rect 191658 477922 222198 477978
rect 222254 477922 222322 477978
rect 222378 477922 252918 477978
rect 252974 477922 253042 477978
rect 253098 477922 283638 477978
rect 283694 477922 283762 477978
rect 283818 477922 314358 477978
rect 314414 477922 314482 477978
rect 314538 477922 345078 477978
rect 345134 477922 345202 477978
rect 345258 477922 375798 477978
rect 375854 477922 375922 477978
rect 375978 477922 406518 477978
rect 406574 477922 406642 477978
rect 406698 477922 437238 477978
rect 437294 477922 437362 477978
rect 437418 477922 467958 477978
rect 468014 477922 468082 477978
rect 468138 477922 498678 477978
rect 498734 477922 498802 477978
rect 498858 477922 529398 477978
rect 529454 477922 529522 477978
rect 529578 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 22518 472350
rect 22574 472294 22642 472350
rect 22698 472294 53238 472350
rect 53294 472294 53362 472350
rect 53418 472294 83958 472350
rect 84014 472294 84082 472350
rect 84138 472294 114678 472350
rect 114734 472294 114802 472350
rect 114858 472294 145398 472350
rect 145454 472294 145522 472350
rect 145578 472294 176118 472350
rect 176174 472294 176242 472350
rect 176298 472294 206838 472350
rect 206894 472294 206962 472350
rect 207018 472294 237558 472350
rect 237614 472294 237682 472350
rect 237738 472294 268278 472350
rect 268334 472294 268402 472350
rect 268458 472294 298998 472350
rect 299054 472294 299122 472350
rect 299178 472294 329718 472350
rect 329774 472294 329842 472350
rect 329898 472294 360438 472350
rect 360494 472294 360562 472350
rect 360618 472294 391158 472350
rect 391214 472294 391282 472350
rect 391338 472294 421878 472350
rect 421934 472294 422002 472350
rect 422058 472294 452598 472350
rect 452654 472294 452722 472350
rect 452778 472294 483318 472350
rect 483374 472294 483442 472350
rect 483498 472294 514038 472350
rect 514094 472294 514162 472350
rect 514218 472294 544758 472350
rect 544814 472294 544882 472350
rect 544938 472294 558474 472350
rect 558530 472294 558598 472350
rect 558654 472294 558722 472350
rect 558778 472294 558846 472350
rect 558902 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 22518 472226
rect 22574 472170 22642 472226
rect 22698 472170 53238 472226
rect 53294 472170 53362 472226
rect 53418 472170 83958 472226
rect 84014 472170 84082 472226
rect 84138 472170 114678 472226
rect 114734 472170 114802 472226
rect 114858 472170 145398 472226
rect 145454 472170 145522 472226
rect 145578 472170 176118 472226
rect 176174 472170 176242 472226
rect 176298 472170 206838 472226
rect 206894 472170 206962 472226
rect 207018 472170 237558 472226
rect 237614 472170 237682 472226
rect 237738 472170 268278 472226
rect 268334 472170 268402 472226
rect 268458 472170 298998 472226
rect 299054 472170 299122 472226
rect 299178 472170 329718 472226
rect 329774 472170 329842 472226
rect 329898 472170 360438 472226
rect 360494 472170 360562 472226
rect 360618 472170 391158 472226
rect 391214 472170 391282 472226
rect 391338 472170 421878 472226
rect 421934 472170 422002 472226
rect 422058 472170 452598 472226
rect 452654 472170 452722 472226
rect 452778 472170 483318 472226
rect 483374 472170 483442 472226
rect 483498 472170 514038 472226
rect 514094 472170 514162 472226
rect 514218 472170 544758 472226
rect 544814 472170 544882 472226
rect 544938 472170 558474 472226
rect 558530 472170 558598 472226
rect 558654 472170 558722 472226
rect 558778 472170 558846 472226
rect 558902 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 22518 472102
rect 22574 472046 22642 472102
rect 22698 472046 53238 472102
rect 53294 472046 53362 472102
rect 53418 472046 83958 472102
rect 84014 472046 84082 472102
rect 84138 472046 114678 472102
rect 114734 472046 114802 472102
rect 114858 472046 145398 472102
rect 145454 472046 145522 472102
rect 145578 472046 176118 472102
rect 176174 472046 176242 472102
rect 176298 472046 206838 472102
rect 206894 472046 206962 472102
rect 207018 472046 237558 472102
rect 237614 472046 237682 472102
rect 237738 472046 268278 472102
rect 268334 472046 268402 472102
rect 268458 472046 298998 472102
rect 299054 472046 299122 472102
rect 299178 472046 329718 472102
rect 329774 472046 329842 472102
rect 329898 472046 360438 472102
rect 360494 472046 360562 472102
rect 360618 472046 391158 472102
rect 391214 472046 391282 472102
rect 391338 472046 421878 472102
rect 421934 472046 422002 472102
rect 422058 472046 452598 472102
rect 452654 472046 452722 472102
rect 452778 472046 483318 472102
rect 483374 472046 483442 472102
rect 483498 472046 514038 472102
rect 514094 472046 514162 472102
rect 514218 472046 544758 472102
rect 544814 472046 544882 472102
rect 544938 472046 558474 472102
rect 558530 472046 558598 472102
rect 558654 472046 558722 472102
rect 558778 472046 558846 472102
rect 558902 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 22518 471978
rect 22574 471922 22642 471978
rect 22698 471922 53238 471978
rect 53294 471922 53362 471978
rect 53418 471922 83958 471978
rect 84014 471922 84082 471978
rect 84138 471922 114678 471978
rect 114734 471922 114802 471978
rect 114858 471922 145398 471978
rect 145454 471922 145522 471978
rect 145578 471922 176118 471978
rect 176174 471922 176242 471978
rect 176298 471922 206838 471978
rect 206894 471922 206962 471978
rect 207018 471922 237558 471978
rect 237614 471922 237682 471978
rect 237738 471922 268278 471978
rect 268334 471922 268402 471978
rect 268458 471922 298998 471978
rect 299054 471922 299122 471978
rect 299178 471922 329718 471978
rect 329774 471922 329842 471978
rect 329898 471922 360438 471978
rect 360494 471922 360562 471978
rect 360618 471922 391158 471978
rect 391214 471922 391282 471978
rect 391338 471922 421878 471978
rect 421934 471922 422002 471978
rect 422058 471922 452598 471978
rect 452654 471922 452722 471978
rect 452778 471922 483318 471978
rect 483374 471922 483442 471978
rect 483498 471922 514038 471978
rect 514094 471922 514162 471978
rect 514218 471922 544758 471978
rect 544814 471922 544882 471978
rect 544938 471922 558474 471978
rect 558530 471922 558598 471978
rect 558654 471922 558722 471978
rect 558778 471922 558846 471978
rect 558902 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 37878 460350
rect 37934 460294 38002 460350
rect 38058 460294 68598 460350
rect 68654 460294 68722 460350
rect 68778 460294 99318 460350
rect 99374 460294 99442 460350
rect 99498 460294 130038 460350
rect 130094 460294 130162 460350
rect 130218 460294 160758 460350
rect 160814 460294 160882 460350
rect 160938 460294 191478 460350
rect 191534 460294 191602 460350
rect 191658 460294 222198 460350
rect 222254 460294 222322 460350
rect 222378 460294 252918 460350
rect 252974 460294 253042 460350
rect 253098 460294 283638 460350
rect 283694 460294 283762 460350
rect 283818 460294 314358 460350
rect 314414 460294 314482 460350
rect 314538 460294 345078 460350
rect 345134 460294 345202 460350
rect 345258 460294 375798 460350
rect 375854 460294 375922 460350
rect 375978 460294 406518 460350
rect 406574 460294 406642 460350
rect 406698 460294 437238 460350
rect 437294 460294 437362 460350
rect 437418 460294 467958 460350
rect 468014 460294 468082 460350
rect 468138 460294 498678 460350
rect 498734 460294 498802 460350
rect 498858 460294 529398 460350
rect 529454 460294 529522 460350
rect 529578 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 37878 460226
rect 37934 460170 38002 460226
rect 38058 460170 68598 460226
rect 68654 460170 68722 460226
rect 68778 460170 99318 460226
rect 99374 460170 99442 460226
rect 99498 460170 130038 460226
rect 130094 460170 130162 460226
rect 130218 460170 160758 460226
rect 160814 460170 160882 460226
rect 160938 460170 191478 460226
rect 191534 460170 191602 460226
rect 191658 460170 222198 460226
rect 222254 460170 222322 460226
rect 222378 460170 252918 460226
rect 252974 460170 253042 460226
rect 253098 460170 283638 460226
rect 283694 460170 283762 460226
rect 283818 460170 314358 460226
rect 314414 460170 314482 460226
rect 314538 460170 345078 460226
rect 345134 460170 345202 460226
rect 345258 460170 375798 460226
rect 375854 460170 375922 460226
rect 375978 460170 406518 460226
rect 406574 460170 406642 460226
rect 406698 460170 437238 460226
rect 437294 460170 437362 460226
rect 437418 460170 467958 460226
rect 468014 460170 468082 460226
rect 468138 460170 498678 460226
rect 498734 460170 498802 460226
rect 498858 460170 529398 460226
rect 529454 460170 529522 460226
rect 529578 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 37878 460102
rect 37934 460046 38002 460102
rect 38058 460046 68598 460102
rect 68654 460046 68722 460102
rect 68778 460046 99318 460102
rect 99374 460046 99442 460102
rect 99498 460046 130038 460102
rect 130094 460046 130162 460102
rect 130218 460046 160758 460102
rect 160814 460046 160882 460102
rect 160938 460046 191478 460102
rect 191534 460046 191602 460102
rect 191658 460046 222198 460102
rect 222254 460046 222322 460102
rect 222378 460046 252918 460102
rect 252974 460046 253042 460102
rect 253098 460046 283638 460102
rect 283694 460046 283762 460102
rect 283818 460046 314358 460102
rect 314414 460046 314482 460102
rect 314538 460046 345078 460102
rect 345134 460046 345202 460102
rect 345258 460046 375798 460102
rect 375854 460046 375922 460102
rect 375978 460046 406518 460102
rect 406574 460046 406642 460102
rect 406698 460046 437238 460102
rect 437294 460046 437362 460102
rect 437418 460046 467958 460102
rect 468014 460046 468082 460102
rect 468138 460046 498678 460102
rect 498734 460046 498802 460102
rect 498858 460046 529398 460102
rect 529454 460046 529522 460102
rect 529578 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 37878 459978
rect 37934 459922 38002 459978
rect 38058 459922 68598 459978
rect 68654 459922 68722 459978
rect 68778 459922 99318 459978
rect 99374 459922 99442 459978
rect 99498 459922 130038 459978
rect 130094 459922 130162 459978
rect 130218 459922 160758 459978
rect 160814 459922 160882 459978
rect 160938 459922 191478 459978
rect 191534 459922 191602 459978
rect 191658 459922 222198 459978
rect 222254 459922 222322 459978
rect 222378 459922 252918 459978
rect 252974 459922 253042 459978
rect 253098 459922 283638 459978
rect 283694 459922 283762 459978
rect 283818 459922 314358 459978
rect 314414 459922 314482 459978
rect 314538 459922 345078 459978
rect 345134 459922 345202 459978
rect 345258 459922 375798 459978
rect 375854 459922 375922 459978
rect 375978 459922 406518 459978
rect 406574 459922 406642 459978
rect 406698 459922 437238 459978
rect 437294 459922 437362 459978
rect 437418 459922 467958 459978
rect 468014 459922 468082 459978
rect 468138 459922 498678 459978
rect 498734 459922 498802 459978
rect 498858 459922 529398 459978
rect 529454 459922 529522 459978
rect 529578 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 22518 454350
rect 22574 454294 22642 454350
rect 22698 454294 53238 454350
rect 53294 454294 53362 454350
rect 53418 454294 83958 454350
rect 84014 454294 84082 454350
rect 84138 454294 114678 454350
rect 114734 454294 114802 454350
rect 114858 454294 145398 454350
rect 145454 454294 145522 454350
rect 145578 454294 176118 454350
rect 176174 454294 176242 454350
rect 176298 454294 206838 454350
rect 206894 454294 206962 454350
rect 207018 454294 237558 454350
rect 237614 454294 237682 454350
rect 237738 454294 268278 454350
rect 268334 454294 268402 454350
rect 268458 454294 298998 454350
rect 299054 454294 299122 454350
rect 299178 454294 329718 454350
rect 329774 454294 329842 454350
rect 329898 454294 360438 454350
rect 360494 454294 360562 454350
rect 360618 454294 391158 454350
rect 391214 454294 391282 454350
rect 391338 454294 421878 454350
rect 421934 454294 422002 454350
rect 422058 454294 452598 454350
rect 452654 454294 452722 454350
rect 452778 454294 483318 454350
rect 483374 454294 483442 454350
rect 483498 454294 514038 454350
rect 514094 454294 514162 454350
rect 514218 454294 544758 454350
rect 544814 454294 544882 454350
rect 544938 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 22518 454226
rect 22574 454170 22642 454226
rect 22698 454170 53238 454226
rect 53294 454170 53362 454226
rect 53418 454170 83958 454226
rect 84014 454170 84082 454226
rect 84138 454170 114678 454226
rect 114734 454170 114802 454226
rect 114858 454170 145398 454226
rect 145454 454170 145522 454226
rect 145578 454170 176118 454226
rect 176174 454170 176242 454226
rect 176298 454170 206838 454226
rect 206894 454170 206962 454226
rect 207018 454170 237558 454226
rect 237614 454170 237682 454226
rect 237738 454170 268278 454226
rect 268334 454170 268402 454226
rect 268458 454170 298998 454226
rect 299054 454170 299122 454226
rect 299178 454170 329718 454226
rect 329774 454170 329842 454226
rect 329898 454170 360438 454226
rect 360494 454170 360562 454226
rect 360618 454170 391158 454226
rect 391214 454170 391282 454226
rect 391338 454170 421878 454226
rect 421934 454170 422002 454226
rect 422058 454170 452598 454226
rect 452654 454170 452722 454226
rect 452778 454170 483318 454226
rect 483374 454170 483442 454226
rect 483498 454170 514038 454226
rect 514094 454170 514162 454226
rect 514218 454170 544758 454226
rect 544814 454170 544882 454226
rect 544938 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 22518 454102
rect 22574 454046 22642 454102
rect 22698 454046 53238 454102
rect 53294 454046 53362 454102
rect 53418 454046 83958 454102
rect 84014 454046 84082 454102
rect 84138 454046 114678 454102
rect 114734 454046 114802 454102
rect 114858 454046 145398 454102
rect 145454 454046 145522 454102
rect 145578 454046 176118 454102
rect 176174 454046 176242 454102
rect 176298 454046 206838 454102
rect 206894 454046 206962 454102
rect 207018 454046 237558 454102
rect 237614 454046 237682 454102
rect 237738 454046 268278 454102
rect 268334 454046 268402 454102
rect 268458 454046 298998 454102
rect 299054 454046 299122 454102
rect 299178 454046 329718 454102
rect 329774 454046 329842 454102
rect 329898 454046 360438 454102
rect 360494 454046 360562 454102
rect 360618 454046 391158 454102
rect 391214 454046 391282 454102
rect 391338 454046 421878 454102
rect 421934 454046 422002 454102
rect 422058 454046 452598 454102
rect 452654 454046 452722 454102
rect 452778 454046 483318 454102
rect 483374 454046 483442 454102
rect 483498 454046 514038 454102
rect 514094 454046 514162 454102
rect 514218 454046 544758 454102
rect 544814 454046 544882 454102
rect 544938 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 22518 453978
rect 22574 453922 22642 453978
rect 22698 453922 53238 453978
rect 53294 453922 53362 453978
rect 53418 453922 83958 453978
rect 84014 453922 84082 453978
rect 84138 453922 114678 453978
rect 114734 453922 114802 453978
rect 114858 453922 145398 453978
rect 145454 453922 145522 453978
rect 145578 453922 176118 453978
rect 176174 453922 176242 453978
rect 176298 453922 206838 453978
rect 206894 453922 206962 453978
rect 207018 453922 237558 453978
rect 237614 453922 237682 453978
rect 237738 453922 268278 453978
rect 268334 453922 268402 453978
rect 268458 453922 298998 453978
rect 299054 453922 299122 453978
rect 299178 453922 329718 453978
rect 329774 453922 329842 453978
rect 329898 453922 360438 453978
rect 360494 453922 360562 453978
rect 360618 453922 391158 453978
rect 391214 453922 391282 453978
rect 391338 453922 421878 453978
rect 421934 453922 422002 453978
rect 422058 453922 452598 453978
rect 452654 453922 452722 453978
rect 452778 453922 483318 453978
rect 483374 453922 483442 453978
rect 483498 453922 514038 453978
rect 514094 453922 514162 453978
rect 514218 453922 544758 453978
rect 544814 453922 544882 453978
rect 544938 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 37878 442350
rect 37934 442294 38002 442350
rect 38058 442294 68598 442350
rect 68654 442294 68722 442350
rect 68778 442294 99318 442350
rect 99374 442294 99442 442350
rect 99498 442294 130038 442350
rect 130094 442294 130162 442350
rect 130218 442294 160758 442350
rect 160814 442294 160882 442350
rect 160938 442294 191478 442350
rect 191534 442294 191602 442350
rect 191658 442294 222198 442350
rect 222254 442294 222322 442350
rect 222378 442294 252918 442350
rect 252974 442294 253042 442350
rect 253098 442294 283638 442350
rect 283694 442294 283762 442350
rect 283818 442294 314358 442350
rect 314414 442294 314482 442350
rect 314538 442294 345078 442350
rect 345134 442294 345202 442350
rect 345258 442294 375798 442350
rect 375854 442294 375922 442350
rect 375978 442294 406518 442350
rect 406574 442294 406642 442350
rect 406698 442294 437238 442350
rect 437294 442294 437362 442350
rect 437418 442294 467958 442350
rect 468014 442294 468082 442350
rect 468138 442294 498678 442350
rect 498734 442294 498802 442350
rect 498858 442294 529398 442350
rect 529454 442294 529522 442350
rect 529578 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 37878 442226
rect 37934 442170 38002 442226
rect 38058 442170 68598 442226
rect 68654 442170 68722 442226
rect 68778 442170 99318 442226
rect 99374 442170 99442 442226
rect 99498 442170 130038 442226
rect 130094 442170 130162 442226
rect 130218 442170 160758 442226
rect 160814 442170 160882 442226
rect 160938 442170 191478 442226
rect 191534 442170 191602 442226
rect 191658 442170 222198 442226
rect 222254 442170 222322 442226
rect 222378 442170 252918 442226
rect 252974 442170 253042 442226
rect 253098 442170 283638 442226
rect 283694 442170 283762 442226
rect 283818 442170 314358 442226
rect 314414 442170 314482 442226
rect 314538 442170 345078 442226
rect 345134 442170 345202 442226
rect 345258 442170 375798 442226
rect 375854 442170 375922 442226
rect 375978 442170 406518 442226
rect 406574 442170 406642 442226
rect 406698 442170 437238 442226
rect 437294 442170 437362 442226
rect 437418 442170 467958 442226
rect 468014 442170 468082 442226
rect 468138 442170 498678 442226
rect 498734 442170 498802 442226
rect 498858 442170 529398 442226
rect 529454 442170 529522 442226
rect 529578 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 37878 442102
rect 37934 442046 38002 442102
rect 38058 442046 68598 442102
rect 68654 442046 68722 442102
rect 68778 442046 99318 442102
rect 99374 442046 99442 442102
rect 99498 442046 130038 442102
rect 130094 442046 130162 442102
rect 130218 442046 160758 442102
rect 160814 442046 160882 442102
rect 160938 442046 191478 442102
rect 191534 442046 191602 442102
rect 191658 442046 222198 442102
rect 222254 442046 222322 442102
rect 222378 442046 252918 442102
rect 252974 442046 253042 442102
rect 253098 442046 283638 442102
rect 283694 442046 283762 442102
rect 283818 442046 314358 442102
rect 314414 442046 314482 442102
rect 314538 442046 345078 442102
rect 345134 442046 345202 442102
rect 345258 442046 375798 442102
rect 375854 442046 375922 442102
rect 375978 442046 406518 442102
rect 406574 442046 406642 442102
rect 406698 442046 437238 442102
rect 437294 442046 437362 442102
rect 437418 442046 467958 442102
rect 468014 442046 468082 442102
rect 468138 442046 498678 442102
rect 498734 442046 498802 442102
rect 498858 442046 529398 442102
rect 529454 442046 529522 442102
rect 529578 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 37878 441978
rect 37934 441922 38002 441978
rect 38058 441922 68598 441978
rect 68654 441922 68722 441978
rect 68778 441922 99318 441978
rect 99374 441922 99442 441978
rect 99498 441922 130038 441978
rect 130094 441922 130162 441978
rect 130218 441922 160758 441978
rect 160814 441922 160882 441978
rect 160938 441922 191478 441978
rect 191534 441922 191602 441978
rect 191658 441922 222198 441978
rect 222254 441922 222322 441978
rect 222378 441922 252918 441978
rect 252974 441922 253042 441978
rect 253098 441922 283638 441978
rect 283694 441922 283762 441978
rect 283818 441922 314358 441978
rect 314414 441922 314482 441978
rect 314538 441922 345078 441978
rect 345134 441922 345202 441978
rect 345258 441922 375798 441978
rect 375854 441922 375922 441978
rect 375978 441922 406518 441978
rect 406574 441922 406642 441978
rect 406698 441922 437238 441978
rect 437294 441922 437362 441978
rect 437418 441922 467958 441978
rect 468014 441922 468082 441978
rect 468138 441922 498678 441978
rect 498734 441922 498802 441978
rect 498858 441922 529398 441978
rect 529454 441922 529522 441978
rect 529578 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 22518 436350
rect 22574 436294 22642 436350
rect 22698 436294 53238 436350
rect 53294 436294 53362 436350
rect 53418 436294 83958 436350
rect 84014 436294 84082 436350
rect 84138 436294 114678 436350
rect 114734 436294 114802 436350
rect 114858 436294 145398 436350
rect 145454 436294 145522 436350
rect 145578 436294 176118 436350
rect 176174 436294 176242 436350
rect 176298 436294 206838 436350
rect 206894 436294 206962 436350
rect 207018 436294 237558 436350
rect 237614 436294 237682 436350
rect 237738 436294 268278 436350
rect 268334 436294 268402 436350
rect 268458 436294 298998 436350
rect 299054 436294 299122 436350
rect 299178 436294 329718 436350
rect 329774 436294 329842 436350
rect 329898 436294 360438 436350
rect 360494 436294 360562 436350
rect 360618 436294 391158 436350
rect 391214 436294 391282 436350
rect 391338 436294 421878 436350
rect 421934 436294 422002 436350
rect 422058 436294 452598 436350
rect 452654 436294 452722 436350
rect 452778 436294 483318 436350
rect 483374 436294 483442 436350
rect 483498 436294 514038 436350
rect 514094 436294 514162 436350
rect 514218 436294 544758 436350
rect 544814 436294 544882 436350
rect 544938 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 22518 436226
rect 22574 436170 22642 436226
rect 22698 436170 53238 436226
rect 53294 436170 53362 436226
rect 53418 436170 83958 436226
rect 84014 436170 84082 436226
rect 84138 436170 114678 436226
rect 114734 436170 114802 436226
rect 114858 436170 145398 436226
rect 145454 436170 145522 436226
rect 145578 436170 176118 436226
rect 176174 436170 176242 436226
rect 176298 436170 206838 436226
rect 206894 436170 206962 436226
rect 207018 436170 237558 436226
rect 237614 436170 237682 436226
rect 237738 436170 268278 436226
rect 268334 436170 268402 436226
rect 268458 436170 298998 436226
rect 299054 436170 299122 436226
rect 299178 436170 329718 436226
rect 329774 436170 329842 436226
rect 329898 436170 360438 436226
rect 360494 436170 360562 436226
rect 360618 436170 391158 436226
rect 391214 436170 391282 436226
rect 391338 436170 421878 436226
rect 421934 436170 422002 436226
rect 422058 436170 452598 436226
rect 452654 436170 452722 436226
rect 452778 436170 483318 436226
rect 483374 436170 483442 436226
rect 483498 436170 514038 436226
rect 514094 436170 514162 436226
rect 514218 436170 544758 436226
rect 544814 436170 544882 436226
rect 544938 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 22518 436102
rect 22574 436046 22642 436102
rect 22698 436046 53238 436102
rect 53294 436046 53362 436102
rect 53418 436046 83958 436102
rect 84014 436046 84082 436102
rect 84138 436046 114678 436102
rect 114734 436046 114802 436102
rect 114858 436046 145398 436102
rect 145454 436046 145522 436102
rect 145578 436046 176118 436102
rect 176174 436046 176242 436102
rect 176298 436046 206838 436102
rect 206894 436046 206962 436102
rect 207018 436046 237558 436102
rect 237614 436046 237682 436102
rect 237738 436046 268278 436102
rect 268334 436046 268402 436102
rect 268458 436046 298998 436102
rect 299054 436046 299122 436102
rect 299178 436046 329718 436102
rect 329774 436046 329842 436102
rect 329898 436046 360438 436102
rect 360494 436046 360562 436102
rect 360618 436046 391158 436102
rect 391214 436046 391282 436102
rect 391338 436046 421878 436102
rect 421934 436046 422002 436102
rect 422058 436046 452598 436102
rect 452654 436046 452722 436102
rect 452778 436046 483318 436102
rect 483374 436046 483442 436102
rect 483498 436046 514038 436102
rect 514094 436046 514162 436102
rect 514218 436046 544758 436102
rect 544814 436046 544882 436102
rect 544938 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 22518 435978
rect 22574 435922 22642 435978
rect 22698 435922 53238 435978
rect 53294 435922 53362 435978
rect 53418 435922 83958 435978
rect 84014 435922 84082 435978
rect 84138 435922 114678 435978
rect 114734 435922 114802 435978
rect 114858 435922 145398 435978
rect 145454 435922 145522 435978
rect 145578 435922 176118 435978
rect 176174 435922 176242 435978
rect 176298 435922 206838 435978
rect 206894 435922 206962 435978
rect 207018 435922 237558 435978
rect 237614 435922 237682 435978
rect 237738 435922 268278 435978
rect 268334 435922 268402 435978
rect 268458 435922 298998 435978
rect 299054 435922 299122 435978
rect 299178 435922 329718 435978
rect 329774 435922 329842 435978
rect 329898 435922 360438 435978
rect 360494 435922 360562 435978
rect 360618 435922 391158 435978
rect 391214 435922 391282 435978
rect 391338 435922 421878 435978
rect 421934 435922 422002 435978
rect 422058 435922 452598 435978
rect 452654 435922 452722 435978
rect 452778 435922 483318 435978
rect 483374 435922 483442 435978
rect 483498 435922 514038 435978
rect 514094 435922 514162 435978
rect 514218 435922 544758 435978
rect 544814 435922 544882 435978
rect 544938 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 37878 424350
rect 37934 424294 38002 424350
rect 38058 424294 68598 424350
rect 68654 424294 68722 424350
rect 68778 424294 99318 424350
rect 99374 424294 99442 424350
rect 99498 424294 130038 424350
rect 130094 424294 130162 424350
rect 130218 424294 160758 424350
rect 160814 424294 160882 424350
rect 160938 424294 191478 424350
rect 191534 424294 191602 424350
rect 191658 424294 222198 424350
rect 222254 424294 222322 424350
rect 222378 424294 252918 424350
rect 252974 424294 253042 424350
rect 253098 424294 283638 424350
rect 283694 424294 283762 424350
rect 283818 424294 314358 424350
rect 314414 424294 314482 424350
rect 314538 424294 345078 424350
rect 345134 424294 345202 424350
rect 345258 424294 375798 424350
rect 375854 424294 375922 424350
rect 375978 424294 406518 424350
rect 406574 424294 406642 424350
rect 406698 424294 437238 424350
rect 437294 424294 437362 424350
rect 437418 424294 467958 424350
rect 468014 424294 468082 424350
rect 468138 424294 498678 424350
rect 498734 424294 498802 424350
rect 498858 424294 529398 424350
rect 529454 424294 529522 424350
rect 529578 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 37878 424226
rect 37934 424170 38002 424226
rect 38058 424170 68598 424226
rect 68654 424170 68722 424226
rect 68778 424170 99318 424226
rect 99374 424170 99442 424226
rect 99498 424170 130038 424226
rect 130094 424170 130162 424226
rect 130218 424170 160758 424226
rect 160814 424170 160882 424226
rect 160938 424170 191478 424226
rect 191534 424170 191602 424226
rect 191658 424170 222198 424226
rect 222254 424170 222322 424226
rect 222378 424170 252918 424226
rect 252974 424170 253042 424226
rect 253098 424170 283638 424226
rect 283694 424170 283762 424226
rect 283818 424170 314358 424226
rect 314414 424170 314482 424226
rect 314538 424170 345078 424226
rect 345134 424170 345202 424226
rect 345258 424170 375798 424226
rect 375854 424170 375922 424226
rect 375978 424170 406518 424226
rect 406574 424170 406642 424226
rect 406698 424170 437238 424226
rect 437294 424170 437362 424226
rect 437418 424170 467958 424226
rect 468014 424170 468082 424226
rect 468138 424170 498678 424226
rect 498734 424170 498802 424226
rect 498858 424170 529398 424226
rect 529454 424170 529522 424226
rect 529578 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 37878 424102
rect 37934 424046 38002 424102
rect 38058 424046 68598 424102
rect 68654 424046 68722 424102
rect 68778 424046 99318 424102
rect 99374 424046 99442 424102
rect 99498 424046 130038 424102
rect 130094 424046 130162 424102
rect 130218 424046 160758 424102
rect 160814 424046 160882 424102
rect 160938 424046 191478 424102
rect 191534 424046 191602 424102
rect 191658 424046 222198 424102
rect 222254 424046 222322 424102
rect 222378 424046 252918 424102
rect 252974 424046 253042 424102
rect 253098 424046 283638 424102
rect 283694 424046 283762 424102
rect 283818 424046 314358 424102
rect 314414 424046 314482 424102
rect 314538 424046 345078 424102
rect 345134 424046 345202 424102
rect 345258 424046 375798 424102
rect 375854 424046 375922 424102
rect 375978 424046 406518 424102
rect 406574 424046 406642 424102
rect 406698 424046 437238 424102
rect 437294 424046 437362 424102
rect 437418 424046 467958 424102
rect 468014 424046 468082 424102
rect 468138 424046 498678 424102
rect 498734 424046 498802 424102
rect 498858 424046 529398 424102
rect 529454 424046 529522 424102
rect 529578 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 37878 423978
rect 37934 423922 38002 423978
rect 38058 423922 68598 423978
rect 68654 423922 68722 423978
rect 68778 423922 99318 423978
rect 99374 423922 99442 423978
rect 99498 423922 130038 423978
rect 130094 423922 130162 423978
rect 130218 423922 160758 423978
rect 160814 423922 160882 423978
rect 160938 423922 191478 423978
rect 191534 423922 191602 423978
rect 191658 423922 222198 423978
rect 222254 423922 222322 423978
rect 222378 423922 252918 423978
rect 252974 423922 253042 423978
rect 253098 423922 283638 423978
rect 283694 423922 283762 423978
rect 283818 423922 314358 423978
rect 314414 423922 314482 423978
rect 314538 423922 345078 423978
rect 345134 423922 345202 423978
rect 345258 423922 375798 423978
rect 375854 423922 375922 423978
rect 375978 423922 406518 423978
rect 406574 423922 406642 423978
rect 406698 423922 437238 423978
rect 437294 423922 437362 423978
rect 437418 423922 467958 423978
rect 468014 423922 468082 423978
rect 468138 423922 498678 423978
rect 498734 423922 498802 423978
rect 498858 423922 529398 423978
rect 529454 423922 529522 423978
rect 529578 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 22518 418350
rect 22574 418294 22642 418350
rect 22698 418294 53238 418350
rect 53294 418294 53362 418350
rect 53418 418294 83958 418350
rect 84014 418294 84082 418350
rect 84138 418294 114678 418350
rect 114734 418294 114802 418350
rect 114858 418294 145398 418350
rect 145454 418294 145522 418350
rect 145578 418294 176118 418350
rect 176174 418294 176242 418350
rect 176298 418294 206838 418350
rect 206894 418294 206962 418350
rect 207018 418294 237558 418350
rect 237614 418294 237682 418350
rect 237738 418294 268278 418350
rect 268334 418294 268402 418350
rect 268458 418294 298998 418350
rect 299054 418294 299122 418350
rect 299178 418294 329718 418350
rect 329774 418294 329842 418350
rect 329898 418294 360438 418350
rect 360494 418294 360562 418350
rect 360618 418294 391158 418350
rect 391214 418294 391282 418350
rect 391338 418294 421878 418350
rect 421934 418294 422002 418350
rect 422058 418294 452598 418350
rect 452654 418294 452722 418350
rect 452778 418294 483318 418350
rect 483374 418294 483442 418350
rect 483498 418294 514038 418350
rect 514094 418294 514162 418350
rect 514218 418294 544758 418350
rect 544814 418294 544882 418350
rect 544938 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 22518 418226
rect 22574 418170 22642 418226
rect 22698 418170 53238 418226
rect 53294 418170 53362 418226
rect 53418 418170 83958 418226
rect 84014 418170 84082 418226
rect 84138 418170 114678 418226
rect 114734 418170 114802 418226
rect 114858 418170 145398 418226
rect 145454 418170 145522 418226
rect 145578 418170 176118 418226
rect 176174 418170 176242 418226
rect 176298 418170 206838 418226
rect 206894 418170 206962 418226
rect 207018 418170 237558 418226
rect 237614 418170 237682 418226
rect 237738 418170 268278 418226
rect 268334 418170 268402 418226
rect 268458 418170 298998 418226
rect 299054 418170 299122 418226
rect 299178 418170 329718 418226
rect 329774 418170 329842 418226
rect 329898 418170 360438 418226
rect 360494 418170 360562 418226
rect 360618 418170 391158 418226
rect 391214 418170 391282 418226
rect 391338 418170 421878 418226
rect 421934 418170 422002 418226
rect 422058 418170 452598 418226
rect 452654 418170 452722 418226
rect 452778 418170 483318 418226
rect 483374 418170 483442 418226
rect 483498 418170 514038 418226
rect 514094 418170 514162 418226
rect 514218 418170 544758 418226
rect 544814 418170 544882 418226
rect 544938 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 22518 418102
rect 22574 418046 22642 418102
rect 22698 418046 53238 418102
rect 53294 418046 53362 418102
rect 53418 418046 83958 418102
rect 84014 418046 84082 418102
rect 84138 418046 114678 418102
rect 114734 418046 114802 418102
rect 114858 418046 145398 418102
rect 145454 418046 145522 418102
rect 145578 418046 176118 418102
rect 176174 418046 176242 418102
rect 176298 418046 206838 418102
rect 206894 418046 206962 418102
rect 207018 418046 237558 418102
rect 237614 418046 237682 418102
rect 237738 418046 268278 418102
rect 268334 418046 268402 418102
rect 268458 418046 298998 418102
rect 299054 418046 299122 418102
rect 299178 418046 329718 418102
rect 329774 418046 329842 418102
rect 329898 418046 360438 418102
rect 360494 418046 360562 418102
rect 360618 418046 391158 418102
rect 391214 418046 391282 418102
rect 391338 418046 421878 418102
rect 421934 418046 422002 418102
rect 422058 418046 452598 418102
rect 452654 418046 452722 418102
rect 452778 418046 483318 418102
rect 483374 418046 483442 418102
rect 483498 418046 514038 418102
rect 514094 418046 514162 418102
rect 514218 418046 544758 418102
rect 544814 418046 544882 418102
rect 544938 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 22518 417978
rect 22574 417922 22642 417978
rect 22698 417922 53238 417978
rect 53294 417922 53362 417978
rect 53418 417922 83958 417978
rect 84014 417922 84082 417978
rect 84138 417922 114678 417978
rect 114734 417922 114802 417978
rect 114858 417922 145398 417978
rect 145454 417922 145522 417978
rect 145578 417922 176118 417978
rect 176174 417922 176242 417978
rect 176298 417922 206838 417978
rect 206894 417922 206962 417978
rect 207018 417922 237558 417978
rect 237614 417922 237682 417978
rect 237738 417922 268278 417978
rect 268334 417922 268402 417978
rect 268458 417922 298998 417978
rect 299054 417922 299122 417978
rect 299178 417922 329718 417978
rect 329774 417922 329842 417978
rect 329898 417922 360438 417978
rect 360494 417922 360562 417978
rect 360618 417922 391158 417978
rect 391214 417922 391282 417978
rect 391338 417922 421878 417978
rect 421934 417922 422002 417978
rect 422058 417922 452598 417978
rect 452654 417922 452722 417978
rect 452778 417922 483318 417978
rect 483374 417922 483442 417978
rect 483498 417922 514038 417978
rect 514094 417922 514162 417978
rect 514218 417922 544758 417978
rect 544814 417922 544882 417978
rect 544938 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 37878 406350
rect 37934 406294 38002 406350
rect 38058 406294 68598 406350
rect 68654 406294 68722 406350
rect 68778 406294 99318 406350
rect 99374 406294 99442 406350
rect 99498 406294 130038 406350
rect 130094 406294 130162 406350
rect 130218 406294 160758 406350
rect 160814 406294 160882 406350
rect 160938 406294 191478 406350
rect 191534 406294 191602 406350
rect 191658 406294 222198 406350
rect 222254 406294 222322 406350
rect 222378 406294 252918 406350
rect 252974 406294 253042 406350
rect 253098 406294 283638 406350
rect 283694 406294 283762 406350
rect 283818 406294 314358 406350
rect 314414 406294 314482 406350
rect 314538 406294 345078 406350
rect 345134 406294 345202 406350
rect 345258 406294 375798 406350
rect 375854 406294 375922 406350
rect 375978 406294 406518 406350
rect 406574 406294 406642 406350
rect 406698 406294 437238 406350
rect 437294 406294 437362 406350
rect 437418 406294 467958 406350
rect 468014 406294 468082 406350
rect 468138 406294 498678 406350
rect 498734 406294 498802 406350
rect 498858 406294 529398 406350
rect 529454 406294 529522 406350
rect 529578 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 37878 406226
rect 37934 406170 38002 406226
rect 38058 406170 68598 406226
rect 68654 406170 68722 406226
rect 68778 406170 99318 406226
rect 99374 406170 99442 406226
rect 99498 406170 130038 406226
rect 130094 406170 130162 406226
rect 130218 406170 160758 406226
rect 160814 406170 160882 406226
rect 160938 406170 191478 406226
rect 191534 406170 191602 406226
rect 191658 406170 222198 406226
rect 222254 406170 222322 406226
rect 222378 406170 252918 406226
rect 252974 406170 253042 406226
rect 253098 406170 283638 406226
rect 283694 406170 283762 406226
rect 283818 406170 314358 406226
rect 314414 406170 314482 406226
rect 314538 406170 345078 406226
rect 345134 406170 345202 406226
rect 345258 406170 375798 406226
rect 375854 406170 375922 406226
rect 375978 406170 406518 406226
rect 406574 406170 406642 406226
rect 406698 406170 437238 406226
rect 437294 406170 437362 406226
rect 437418 406170 467958 406226
rect 468014 406170 468082 406226
rect 468138 406170 498678 406226
rect 498734 406170 498802 406226
rect 498858 406170 529398 406226
rect 529454 406170 529522 406226
rect 529578 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 37878 406102
rect 37934 406046 38002 406102
rect 38058 406046 68598 406102
rect 68654 406046 68722 406102
rect 68778 406046 99318 406102
rect 99374 406046 99442 406102
rect 99498 406046 130038 406102
rect 130094 406046 130162 406102
rect 130218 406046 160758 406102
rect 160814 406046 160882 406102
rect 160938 406046 191478 406102
rect 191534 406046 191602 406102
rect 191658 406046 222198 406102
rect 222254 406046 222322 406102
rect 222378 406046 252918 406102
rect 252974 406046 253042 406102
rect 253098 406046 283638 406102
rect 283694 406046 283762 406102
rect 283818 406046 314358 406102
rect 314414 406046 314482 406102
rect 314538 406046 345078 406102
rect 345134 406046 345202 406102
rect 345258 406046 375798 406102
rect 375854 406046 375922 406102
rect 375978 406046 406518 406102
rect 406574 406046 406642 406102
rect 406698 406046 437238 406102
rect 437294 406046 437362 406102
rect 437418 406046 467958 406102
rect 468014 406046 468082 406102
rect 468138 406046 498678 406102
rect 498734 406046 498802 406102
rect 498858 406046 529398 406102
rect 529454 406046 529522 406102
rect 529578 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 37878 405978
rect 37934 405922 38002 405978
rect 38058 405922 68598 405978
rect 68654 405922 68722 405978
rect 68778 405922 99318 405978
rect 99374 405922 99442 405978
rect 99498 405922 130038 405978
rect 130094 405922 130162 405978
rect 130218 405922 160758 405978
rect 160814 405922 160882 405978
rect 160938 405922 191478 405978
rect 191534 405922 191602 405978
rect 191658 405922 222198 405978
rect 222254 405922 222322 405978
rect 222378 405922 252918 405978
rect 252974 405922 253042 405978
rect 253098 405922 283638 405978
rect 283694 405922 283762 405978
rect 283818 405922 314358 405978
rect 314414 405922 314482 405978
rect 314538 405922 345078 405978
rect 345134 405922 345202 405978
rect 345258 405922 375798 405978
rect 375854 405922 375922 405978
rect 375978 405922 406518 405978
rect 406574 405922 406642 405978
rect 406698 405922 437238 405978
rect 437294 405922 437362 405978
rect 437418 405922 467958 405978
rect 468014 405922 468082 405978
rect 468138 405922 498678 405978
rect 498734 405922 498802 405978
rect 498858 405922 529398 405978
rect 529454 405922 529522 405978
rect 529578 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 22518 400350
rect 22574 400294 22642 400350
rect 22698 400294 53238 400350
rect 53294 400294 53362 400350
rect 53418 400294 83958 400350
rect 84014 400294 84082 400350
rect 84138 400294 114678 400350
rect 114734 400294 114802 400350
rect 114858 400294 145398 400350
rect 145454 400294 145522 400350
rect 145578 400294 176118 400350
rect 176174 400294 176242 400350
rect 176298 400294 206838 400350
rect 206894 400294 206962 400350
rect 207018 400294 237558 400350
rect 237614 400294 237682 400350
rect 237738 400294 268278 400350
rect 268334 400294 268402 400350
rect 268458 400294 298998 400350
rect 299054 400294 299122 400350
rect 299178 400294 329718 400350
rect 329774 400294 329842 400350
rect 329898 400294 360438 400350
rect 360494 400294 360562 400350
rect 360618 400294 391158 400350
rect 391214 400294 391282 400350
rect 391338 400294 421878 400350
rect 421934 400294 422002 400350
rect 422058 400294 452598 400350
rect 452654 400294 452722 400350
rect 452778 400294 483318 400350
rect 483374 400294 483442 400350
rect 483498 400294 514038 400350
rect 514094 400294 514162 400350
rect 514218 400294 544758 400350
rect 544814 400294 544882 400350
rect 544938 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 22518 400226
rect 22574 400170 22642 400226
rect 22698 400170 53238 400226
rect 53294 400170 53362 400226
rect 53418 400170 83958 400226
rect 84014 400170 84082 400226
rect 84138 400170 114678 400226
rect 114734 400170 114802 400226
rect 114858 400170 145398 400226
rect 145454 400170 145522 400226
rect 145578 400170 176118 400226
rect 176174 400170 176242 400226
rect 176298 400170 206838 400226
rect 206894 400170 206962 400226
rect 207018 400170 237558 400226
rect 237614 400170 237682 400226
rect 237738 400170 268278 400226
rect 268334 400170 268402 400226
rect 268458 400170 298998 400226
rect 299054 400170 299122 400226
rect 299178 400170 329718 400226
rect 329774 400170 329842 400226
rect 329898 400170 360438 400226
rect 360494 400170 360562 400226
rect 360618 400170 391158 400226
rect 391214 400170 391282 400226
rect 391338 400170 421878 400226
rect 421934 400170 422002 400226
rect 422058 400170 452598 400226
rect 452654 400170 452722 400226
rect 452778 400170 483318 400226
rect 483374 400170 483442 400226
rect 483498 400170 514038 400226
rect 514094 400170 514162 400226
rect 514218 400170 544758 400226
rect 544814 400170 544882 400226
rect 544938 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 22518 400102
rect 22574 400046 22642 400102
rect 22698 400046 53238 400102
rect 53294 400046 53362 400102
rect 53418 400046 83958 400102
rect 84014 400046 84082 400102
rect 84138 400046 114678 400102
rect 114734 400046 114802 400102
rect 114858 400046 145398 400102
rect 145454 400046 145522 400102
rect 145578 400046 176118 400102
rect 176174 400046 176242 400102
rect 176298 400046 206838 400102
rect 206894 400046 206962 400102
rect 207018 400046 237558 400102
rect 237614 400046 237682 400102
rect 237738 400046 268278 400102
rect 268334 400046 268402 400102
rect 268458 400046 298998 400102
rect 299054 400046 299122 400102
rect 299178 400046 329718 400102
rect 329774 400046 329842 400102
rect 329898 400046 360438 400102
rect 360494 400046 360562 400102
rect 360618 400046 391158 400102
rect 391214 400046 391282 400102
rect 391338 400046 421878 400102
rect 421934 400046 422002 400102
rect 422058 400046 452598 400102
rect 452654 400046 452722 400102
rect 452778 400046 483318 400102
rect 483374 400046 483442 400102
rect 483498 400046 514038 400102
rect 514094 400046 514162 400102
rect 514218 400046 544758 400102
rect 544814 400046 544882 400102
rect 544938 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 22518 399978
rect 22574 399922 22642 399978
rect 22698 399922 53238 399978
rect 53294 399922 53362 399978
rect 53418 399922 83958 399978
rect 84014 399922 84082 399978
rect 84138 399922 114678 399978
rect 114734 399922 114802 399978
rect 114858 399922 145398 399978
rect 145454 399922 145522 399978
rect 145578 399922 176118 399978
rect 176174 399922 176242 399978
rect 176298 399922 206838 399978
rect 206894 399922 206962 399978
rect 207018 399922 237558 399978
rect 237614 399922 237682 399978
rect 237738 399922 268278 399978
rect 268334 399922 268402 399978
rect 268458 399922 298998 399978
rect 299054 399922 299122 399978
rect 299178 399922 329718 399978
rect 329774 399922 329842 399978
rect 329898 399922 360438 399978
rect 360494 399922 360562 399978
rect 360618 399922 391158 399978
rect 391214 399922 391282 399978
rect 391338 399922 421878 399978
rect 421934 399922 422002 399978
rect 422058 399922 452598 399978
rect 452654 399922 452722 399978
rect 452778 399922 483318 399978
rect 483374 399922 483442 399978
rect 483498 399922 514038 399978
rect 514094 399922 514162 399978
rect 514218 399922 544758 399978
rect 544814 399922 544882 399978
rect 544938 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 443084 392518 548116 392534
rect 443084 392462 443100 392518
rect 443156 392462 548044 392518
rect 548100 392462 548116 392518
rect 443084 392446 548116 392462
rect 439948 392338 590900 392354
rect 439948 392282 439964 392338
rect 440020 392282 590828 392338
rect 590884 392282 590900 392338
rect 439948 392266 590900 392282
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 37782 370350
rect 37838 370294 37906 370350
rect 37962 370294 68502 370350
rect 68558 370294 68626 370350
rect 68682 370294 99222 370350
rect 99278 370294 99346 370350
rect 99402 370294 129942 370350
rect 129998 370294 130066 370350
rect 130122 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193878 370350
rect 193934 370294 194002 370350
rect 194058 370294 224598 370350
rect 224654 370294 224722 370350
rect 224778 370294 255318 370350
rect 255374 370294 255442 370350
rect 255498 370294 286038 370350
rect 286094 370294 286162 370350
rect 286218 370294 316758 370350
rect 316814 370294 316882 370350
rect 316938 370294 347478 370350
rect 347534 370294 347602 370350
rect 347658 370294 378198 370350
rect 378254 370294 378322 370350
rect 378378 370294 408918 370350
rect 408974 370294 409042 370350
rect 409098 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 463878 370350
rect 463934 370294 464002 370350
rect 464058 370294 494598 370350
rect 494654 370294 494722 370350
rect 494778 370294 525318 370350
rect 525374 370294 525442 370350
rect 525498 370294 556038 370350
rect 556094 370294 556162 370350
rect 556218 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 37782 370226
rect 37838 370170 37906 370226
rect 37962 370170 68502 370226
rect 68558 370170 68626 370226
rect 68682 370170 99222 370226
rect 99278 370170 99346 370226
rect 99402 370170 129942 370226
rect 129998 370170 130066 370226
rect 130122 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193878 370226
rect 193934 370170 194002 370226
rect 194058 370170 224598 370226
rect 224654 370170 224722 370226
rect 224778 370170 255318 370226
rect 255374 370170 255442 370226
rect 255498 370170 286038 370226
rect 286094 370170 286162 370226
rect 286218 370170 316758 370226
rect 316814 370170 316882 370226
rect 316938 370170 347478 370226
rect 347534 370170 347602 370226
rect 347658 370170 378198 370226
rect 378254 370170 378322 370226
rect 378378 370170 408918 370226
rect 408974 370170 409042 370226
rect 409098 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 463878 370226
rect 463934 370170 464002 370226
rect 464058 370170 494598 370226
rect 494654 370170 494722 370226
rect 494778 370170 525318 370226
rect 525374 370170 525442 370226
rect 525498 370170 556038 370226
rect 556094 370170 556162 370226
rect 556218 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 37782 370102
rect 37838 370046 37906 370102
rect 37962 370046 68502 370102
rect 68558 370046 68626 370102
rect 68682 370046 99222 370102
rect 99278 370046 99346 370102
rect 99402 370046 129942 370102
rect 129998 370046 130066 370102
rect 130122 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193878 370102
rect 193934 370046 194002 370102
rect 194058 370046 224598 370102
rect 224654 370046 224722 370102
rect 224778 370046 255318 370102
rect 255374 370046 255442 370102
rect 255498 370046 286038 370102
rect 286094 370046 286162 370102
rect 286218 370046 316758 370102
rect 316814 370046 316882 370102
rect 316938 370046 347478 370102
rect 347534 370046 347602 370102
rect 347658 370046 378198 370102
rect 378254 370046 378322 370102
rect 378378 370046 408918 370102
rect 408974 370046 409042 370102
rect 409098 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 463878 370102
rect 463934 370046 464002 370102
rect 464058 370046 494598 370102
rect 494654 370046 494722 370102
rect 494778 370046 525318 370102
rect 525374 370046 525442 370102
rect 525498 370046 556038 370102
rect 556094 370046 556162 370102
rect 556218 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 37782 369978
rect 37838 369922 37906 369978
rect 37962 369922 68502 369978
rect 68558 369922 68626 369978
rect 68682 369922 99222 369978
rect 99278 369922 99346 369978
rect 99402 369922 129942 369978
rect 129998 369922 130066 369978
rect 130122 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193878 369978
rect 193934 369922 194002 369978
rect 194058 369922 224598 369978
rect 224654 369922 224722 369978
rect 224778 369922 255318 369978
rect 255374 369922 255442 369978
rect 255498 369922 286038 369978
rect 286094 369922 286162 369978
rect 286218 369922 316758 369978
rect 316814 369922 316882 369978
rect 316938 369922 347478 369978
rect 347534 369922 347602 369978
rect 347658 369922 378198 369978
rect 378254 369922 378322 369978
rect 378378 369922 408918 369978
rect 408974 369922 409042 369978
rect 409098 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 463878 369978
rect 463934 369922 464002 369978
rect 464058 369922 494598 369978
rect 494654 369922 494722 369978
rect 494778 369922 525318 369978
rect 525374 369922 525442 369978
rect 525498 369922 556038 369978
rect 556094 369922 556162 369978
rect 556218 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 22422 364350
rect 22478 364294 22546 364350
rect 22602 364294 53142 364350
rect 53198 364294 53266 364350
rect 53322 364294 83862 364350
rect 83918 364294 83986 364350
rect 84042 364294 114582 364350
rect 114638 364294 114706 364350
rect 114762 364294 145302 364350
rect 145358 364294 145426 364350
rect 145482 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 178518 364350
rect 178574 364294 178642 364350
rect 178698 364294 209238 364350
rect 209294 364294 209362 364350
rect 209418 364294 239958 364350
rect 240014 364294 240082 364350
rect 240138 364294 270678 364350
rect 270734 364294 270802 364350
rect 270858 364294 301398 364350
rect 301454 364294 301522 364350
rect 301578 364294 332118 364350
rect 332174 364294 332242 364350
rect 332298 364294 362838 364350
rect 362894 364294 362962 364350
rect 363018 364294 393558 364350
rect 393614 364294 393682 364350
rect 393738 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 448518 364350
rect 448574 364294 448642 364350
rect 448698 364294 479238 364350
rect 479294 364294 479362 364350
rect 479418 364294 509958 364350
rect 510014 364294 510082 364350
rect 510138 364294 540678 364350
rect 540734 364294 540802 364350
rect 540858 364294 571398 364350
rect 571454 364294 571522 364350
rect 571578 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 22422 364226
rect 22478 364170 22546 364226
rect 22602 364170 53142 364226
rect 53198 364170 53266 364226
rect 53322 364170 83862 364226
rect 83918 364170 83986 364226
rect 84042 364170 114582 364226
rect 114638 364170 114706 364226
rect 114762 364170 145302 364226
rect 145358 364170 145426 364226
rect 145482 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 178518 364226
rect 178574 364170 178642 364226
rect 178698 364170 209238 364226
rect 209294 364170 209362 364226
rect 209418 364170 239958 364226
rect 240014 364170 240082 364226
rect 240138 364170 270678 364226
rect 270734 364170 270802 364226
rect 270858 364170 301398 364226
rect 301454 364170 301522 364226
rect 301578 364170 332118 364226
rect 332174 364170 332242 364226
rect 332298 364170 362838 364226
rect 362894 364170 362962 364226
rect 363018 364170 393558 364226
rect 393614 364170 393682 364226
rect 393738 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 448518 364226
rect 448574 364170 448642 364226
rect 448698 364170 479238 364226
rect 479294 364170 479362 364226
rect 479418 364170 509958 364226
rect 510014 364170 510082 364226
rect 510138 364170 540678 364226
rect 540734 364170 540802 364226
rect 540858 364170 571398 364226
rect 571454 364170 571522 364226
rect 571578 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 22422 364102
rect 22478 364046 22546 364102
rect 22602 364046 53142 364102
rect 53198 364046 53266 364102
rect 53322 364046 83862 364102
rect 83918 364046 83986 364102
rect 84042 364046 114582 364102
rect 114638 364046 114706 364102
rect 114762 364046 145302 364102
rect 145358 364046 145426 364102
rect 145482 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 178518 364102
rect 178574 364046 178642 364102
rect 178698 364046 209238 364102
rect 209294 364046 209362 364102
rect 209418 364046 239958 364102
rect 240014 364046 240082 364102
rect 240138 364046 270678 364102
rect 270734 364046 270802 364102
rect 270858 364046 301398 364102
rect 301454 364046 301522 364102
rect 301578 364046 332118 364102
rect 332174 364046 332242 364102
rect 332298 364046 362838 364102
rect 362894 364046 362962 364102
rect 363018 364046 393558 364102
rect 393614 364046 393682 364102
rect 393738 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 448518 364102
rect 448574 364046 448642 364102
rect 448698 364046 479238 364102
rect 479294 364046 479362 364102
rect 479418 364046 509958 364102
rect 510014 364046 510082 364102
rect 510138 364046 540678 364102
rect 540734 364046 540802 364102
rect 540858 364046 571398 364102
rect 571454 364046 571522 364102
rect 571578 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 22422 363978
rect 22478 363922 22546 363978
rect 22602 363922 53142 363978
rect 53198 363922 53266 363978
rect 53322 363922 83862 363978
rect 83918 363922 83986 363978
rect 84042 363922 114582 363978
rect 114638 363922 114706 363978
rect 114762 363922 145302 363978
rect 145358 363922 145426 363978
rect 145482 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 178518 363978
rect 178574 363922 178642 363978
rect 178698 363922 209238 363978
rect 209294 363922 209362 363978
rect 209418 363922 239958 363978
rect 240014 363922 240082 363978
rect 240138 363922 270678 363978
rect 270734 363922 270802 363978
rect 270858 363922 301398 363978
rect 301454 363922 301522 363978
rect 301578 363922 332118 363978
rect 332174 363922 332242 363978
rect 332298 363922 362838 363978
rect 362894 363922 362962 363978
rect 363018 363922 393558 363978
rect 393614 363922 393682 363978
rect 393738 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 448518 363978
rect 448574 363922 448642 363978
rect 448698 363922 479238 363978
rect 479294 363922 479362 363978
rect 479418 363922 509958 363978
rect 510014 363922 510082 363978
rect 510138 363922 540678 363978
rect 540734 363922 540802 363978
rect 540858 363922 571398 363978
rect 571454 363922 571522 363978
rect 571578 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 37782 352350
rect 37838 352294 37906 352350
rect 37962 352294 68502 352350
rect 68558 352294 68626 352350
rect 68682 352294 99222 352350
rect 99278 352294 99346 352350
rect 99402 352294 129942 352350
rect 129998 352294 130066 352350
rect 130122 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 193878 352350
rect 193934 352294 194002 352350
rect 194058 352294 224598 352350
rect 224654 352294 224722 352350
rect 224778 352294 255318 352350
rect 255374 352294 255442 352350
rect 255498 352294 286038 352350
rect 286094 352294 286162 352350
rect 286218 352294 316758 352350
rect 316814 352294 316882 352350
rect 316938 352294 347478 352350
rect 347534 352294 347602 352350
rect 347658 352294 378198 352350
rect 378254 352294 378322 352350
rect 378378 352294 408918 352350
rect 408974 352294 409042 352350
rect 409098 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 463878 352350
rect 463934 352294 464002 352350
rect 464058 352294 494598 352350
rect 494654 352294 494722 352350
rect 494778 352294 525318 352350
rect 525374 352294 525442 352350
rect 525498 352294 556038 352350
rect 556094 352294 556162 352350
rect 556218 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 37782 352226
rect 37838 352170 37906 352226
rect 37962 352170 68502 352226
rect 68558 352170 68626 352226
rect 68682 352170 99222 352226
rect 99278 352170 99346 352226
rect 99402 352170 129942 352226
rect 129998 352170 130066 352226
rect 130122 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 193878 352226
rect 193934 352170 194002 352226
rect 194058 352170 224598 352226
rect 224654 352170 224722 352226
rect 224778 352170 255318 352226
rect 255374 352170 255442 352226
rect 255498 352170 286038 352226
rect 286094 352170 286162 352226
rect 286218 352170 316758 352226
rect 316814 352170 316882 352226
rect 316938 352170 347478 352226
rect 347534 352170 347602 352226
rect 347658 352170 378198 352226
rect 378254 352170 378322 352226
rect 378378 352170 408918 352226
rect 408974 352170 409042 352226
rect 409098 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 463878 352226
rect 463934 352170 464002 352226
rect 464058 352170 494598 352226
rect 494654 352170 494722 352226
rect 494778 352170 525318 352226
rect 525374 352170 525442 352226
rect 525498 352170 556038 352226
rect 556094 352170 556162 352226
rect 556218 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 37782 352102
rect 37838 352046 37906 352102
rect 37962 352046 68502 352102
rect 68558 352046 68626 352102
rect 68682 352046 99222 352102
rect 99278 352046 99346 352102
rect 99402 352046 129942 352102
rect 129998 352046 130066 352102
rect 130122 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 193878 352102
rect 193934 352046 194002 352102
rect 194058 352046 224598 352102
rect 224654 352046 224722 352102
rect 224778 352046 255318 352102
rect 255374 352046 255442 352102
rect 255498 352046 286038 352102
rect 286094 352046 286162 352102
rect 286218 352046 316758 352102
rect 316814 352046 316882 352102
rect 316938 352046 347478 352102
rect 347534 352046 347602 352102
rect 347658 352046 378198 352102
rect 378254 352046 378322 352102
rect 378378 352046 408918 352102
rect 408974 352046 409042 352102
rect 409098 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 463878 352102
rect 463934 352046 464002 352102
rect 464058 352046 494598 352102
rect 494654 352046 494722 352102
rect 494778 352046 525318 352102
rect 525374 352046 525442 352102
rect 525498 352046 556038 352102
rect 556094 352046 556162 352102
rect 556218 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 37782 351978
rect 37838 351922 37906 351978
rect 37962 351922 68502 351978
rect 68558 351922 68626 351978
rect 68682 351922 99222 351978
rect 99278 351922 99346 351978
rect 99402 351922 129942 351978
rect 129998 351922 130066 351978
rect 130122 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 193878 351978
rect 193934 351922 194002 351978
rect 194058 351922 224598 351978
rect 224654 351922 224722 351978
rect 224778 351922 255318 351978
rect 255374 351922 255442 351978
rect 255498 351922 286038 351978
rect 286094 351922 286162 351978
rect 286218 351922 316758 351978
rect 316814 351922 316882 351978
rect 316938 351922 347478 351978
rect 347534 351922 347602 351978
rect 347658 351922 378198 351978
rect 378254 351922 378322 351978
rect 378378 351922 408918 351978
rect 408974 351922 409042 351978
rect 409098 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 463878 351978
rect 463934 351922 464002 351978
rect 464058 351922 494598 351978
rect 494654 351922 494722 351978
rect 494778 351922 525318 351978
rect 525374 351922 525442 351978
rect 525498 351922 556038 351978
rect 556094 351922 556162 351978
rect 556218 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 22422 346350
rect 22478 346294 22546 346350
rect 22602 346294 53142 346350
rect 53198 346294 53266 346350
rect 53322 346294 83862 346350
rect 83918 346294 83986 346350
rect 84042 346294 114582 346350
rect 114638 346294 114706 346350
rect 114762 346294 145302 346350
rect 145358 346294 145426 346350
rect 145482 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 178518 346350
rect 178574 346294 178642 346350
rect 178698 346294 209238 346350
rect 209294 346294 209362 346350
rect 209418 346294 239958 346350
rect 240014 346294 240082 346350
rect 240138 346294 270678 346350
rect 270734 346294 270802 346350
rect 270858 346294 301398 346350
rect 301454 346294 301522 346350
rect 301578 346294 332118 346350
rect 332174 346294 332242 346350
rect 332298 346294 362838 346350
rect 362894 346294 362962 346350
rect 363018 346294 393558 346350
rect 393614 346294 393682 346350
rect 393738 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 448518 346350
rect 448574 346294 448642 346350
rect 448698 346294 479238 346350
rect 479294 346294 479362 346350
rect 479418 346294 509958 346350
rect 510014 346294 510082 346350
rect 510138 346294 540678 346350
rect 540734 346294 540802 346350
rect 540858 346294 571398 346350
rect 571454 346294 571522 346350
rect 571578 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 22422 346226
rect 22478 346170 22546 346226
rect 22602 346170 53142 346226
rect 53198 346170 53266 346226
rect 53322 346170 83862 346226
rect 83918 346170 83986 346226
rect 84042 346170 114582 346226
rect 114638 346170 114706 346226
rect 114762 346170 145302 346226
rect 145358 346170 145426 346226
rect 145482 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 178518 346226
rect 178574 346170 178642 346226
rect 178698 346170 209238 346226
rect 209294 346170 209362 346226
rect 209418 346170 239958 346226
rect 240014 346170 240082 346226
rect 240138 346170 270678 346226
rect 270734 346170 270802 346226
rect 270858 346170 301398 346226
rect 301454 346170 301522 346226
rect 301578 346170 332118 346226
rect 332174 346170 332242 346226
rect 332298 346170 362838 346226
rect 362894 346170 362962 346226
rect 363018 346170 393558 346226
rect 393614 346170 393682 346226
rect 393738 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 448518 346226
rect 448574 346170 448642 346226
rect 448698 346170 479238 346226
rect 479294 346170 479362 346226
rect 479418 346170 509958 346226
rect 510014 346170 510082 346226
rect 510138 346170 540678 346226
rect 540734 346170 540802 346226
rect 540858 346170 571398 346226
rect 571454 346170 571522 346226
rect 571578 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 22422 346102
rect 22478 346046 22546 346102
rect 22602 346046 53142 346102
rect 53198 346046 53266 346102
rect 53322 346046 83862 346102
rect 83918 346046 83986 346102
rect 84042 346046 114582 346102
rect 114638 346046 114706 346102
rect 114762 346046 145302 346102
rect 145358 346046 145426 346102
rect 145482 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 178518 346102
rect 178574 346046 178642 346102
rect 178698 346046 209238 346102
rect 209294 346046 209362 346102
rect 209418 346046 239958 346102
rect 240014 346046 240082 346102
rect 240138 346046 270678 346102
rect 270734 346046 270802 346102
rect 270858 346046 301398 346102
rect 301454 346046 301522 346102
rect 301578 346046 332118 346102
rect 332174 346046 332242 346102
rect 332298 346046 362838 346102
rect 362894 346046 362962 346102
rect 363018 346046 393558 346102
rect 393614 346046 393682 346102
rect 393738 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 448518 346102
rect 448574 346046 448642 346102
rect 448698 346046 479238 346102
rect 479294 346046 479362 346102
rect 479418 346046 509958 346102
rect 510014 346046 510082 346102
rect 510138 346046 540678 346102
rect 540734 346046 540802 346102
rect 540858 346046 571398 346102
rect 571454 346046 571522 346102
rect 571578 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 22422 345978
rect 22478 345922 22546 345978
rect 22602 345922 53142 345978
rect 53198 345922 53266 345978
rect 53322 345922 83862 345978
rect 83918 345922 83986 345978
rect 84042 345922 114582 345978
rect 114638 345922 114706 345978
rect 114762 345922 145302 345978
rect 145358 345922 145426 345978
rect 145482 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 178518 345978
rect 178574 345922 178642 345978
rect 178698 345922 209238 345978
rect 209294 345922 209362 345978
rect 209418 345922 239958 345978
rect 240014 345922 240082 345978
rect 240138 345922 270678 345978
rect 270734 345922 270802 345978
rect 270858 345922 301398 345978
rect 301454 345922 301522 345978
rect 301578 345922 332118 345978
rect 332174 345922 332242 345978
rect 332298 345922 362838 345978
rect 362894 345922 362962 345978
rect 363018 345922 393558 345978
rect 393614 345922 393682 345978
rect 393738 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 448518 345978
rect 448574 345922 448642 345978
rect 448698 345922 479238 345978
rect 479294 345922 479362 345978
rect 479418 345922 509958 345978
rect 510014 345922 510082 345978
rect 510138 345922 540678 345978
rect 540734 345922 540802 345978
rect 540858 345922 571398 345978
rect 571454 345922 571522 345978
rect 571578 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 37782 334350
rect 37838 334294 37906 334350
rect 37962 334294 68502 334350
rect 68558 334294 68626 334350
rect 68682 334294 99222 334350
rect 99278 334294 99346 334350
rect 99402 334294 129942 334350
rect 129998 334294 130066 334350
rect 130122 334294 162834 334350
rect 162890 334294 162958 334350
rect 163014 334294 163082 334350
rect 163138 334294 163206 334350
rect 163262 334294 193878 334350
rect 193934 334294 194002 334350
rect 194058 334294 224598 334350
rect 224654 334294 224722 334350
rect 224778 334294 255318 334350
rect 255374 334294 255442 334350
rect 255498 334294 286038 334350
rect 286094 334294 286162 334350
rect 286218 334294 316758 334350
rect 316814 334294 316882 334350
rect 316938 334294 347478 334350
rect 347534 334294 347602 334350
rect 347658 334294 378198 334350
rect 378254 334294 378322 334350
rect 378378 334294 408918 334350
rect 408974 334294 409042 334350
rect 409098 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 463878 334350
rect 463934 334294 464002 334350
rect 464058 334294 494598 334350
rect 494654 334294 494722 334350
rect 494778 334294 525318 334350
rect 525374 334294 525442 334350
rect 525498 334294 556038 334350
rect 556094 334294 556162 334350
rect 556218 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 37782 334226
rect 37838 334170 37906 334226
rect 37962 334170 68502 334226
rect 68558 334170 68626 334226
rect 68682 334170 99222 334226
rect 99278 334170 99346 334226
rect 99402 334170 129942 334226
rect 129998 334170 130066 334226
rect 130122 334170 162834 334226
rect 162890 334170 162958 334226
rect 163014 334170 163082 334226
rect 163138 334170 163206 334226
rect 163262 334170 193878 334226
rect 193934 334170 194002 334226
rect 194058 334170 224598 334226
rect 224654 334170 224722 334226
rect 224778 334170 255318 334226
rect 255374 334170 255442 334226
rect 255498 334170 286038 334226
rect 286094 334170 286162 334226
rect 286218 334170 316758 334226
rect 316814 334170 316882 334226
rect 316938 334170 347478 334226
rect 347534 334170 347602 334226
rect 347658 334170 378198 334226
rect 378254 334170 378322 334226
rect 378378 334170 408918 334226
rect 408974 334170 409042 334226
rect 409098 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 463878 334226
rect 463934 334170 464002 334226
rect 464058 334170 494598 334226
rect 494654 334170 494722 334226
rect 494778 334170 525318 334226
rect 525374 334170 525442 334226
rect 525498 334170 556038 334226
rect 556094 334170 556162 334226
rect 556218 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 37782 334102
rect 37838 334046 37906 334102
rect 37962 334046 68502 334102
rect 68558 334046 68626 334102
rect 68682 334046 99222 334102
rect 99278 334046 99346 334102
rect 99402 334046 129942 334102
rect 129998 334046 130066 334102
rect 130122 334046 162834 334102
rect 162890 334046 162958 334102
rect 163014 334046 163082 334102
rect 163138 334046 163206 334102
rect 163262 334046 193878 334102
rect 193934 334046 194002 334102
rect 194058 334046 224598 334102
rect 224654 334046 224722 334102
rect 224778 334046 255318 334102
rect 255374 334046 255442 334102
rect 255498 334046 286038 334102
rect 286094 334046 286162 334102
rect 286218 334046 316758 334102
rect 316814 334046 316882 334102
rect 316938 334046 347478 334102
rect 347534 334046 347602 334102
rect 347658 334046 378198 334102
rect 378254 334046 378322 334102
rect 378378 334046 408918 334102
rect 408974 334046 409042 334102
rect 409098 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 463878 334102
rect 463934 334046 464002 334102
rect 464058 334046 494598 334102
rect 494654 334046 494722 334102
rect 494778 334046 525318 334102
rect 525374 334046 525442 334102
rect 525498 334046 556038 334102
rect 556094 334046 556162 334102
rect 556218 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 37782 333978
rect 37838 333922 37906 333978
rect 37962 333922 68502 333978
rect 68558 333922 68626 333978
rect 68682 333922 99222 333978
rect 99278 333922 99346 333978
rect 99402 333922 129942 333978
rect 129998 333922 130066 333978
rect 130122 333922 162834 333978
rect 162890 333922 162958 333978
rect 163014 333922 163082 333978
rect 163138 333922 163206 333978
rect 163262 333922 193878 333978
rect 193934 333922 194002 333978
rect 194058 333922 224598 333978
rect 224654 333922 224722 333978
rect 224778 333922 255318 333978
rect 255374 333922 255442 333978
rect 255498 333922 286038 333978
rect 286094 333922 286162 333978
rect 286218 333922 316758 333978
rect 316814 333922 316882 333978
rect 316938 333922 347478 333978
rect 347534 333922 347602 333978
rect 347658 333922 378198 333978
rect 378254 333922 378322 333978
rect 378378 333922 408918 333978
rect 408974 333922 409042 333978
rect 409098 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 463878 333978
rect 463934 333922 464002 333978
rect 464058 333922 494598 333978
rect 494654 333922 494722 333978
rect 494778 333922 525318 333978
rect 525374 333922 525442 333978
rect 525498 333922 556038 333978
rect 556094 333922 556162 333978
rect 556218 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 22422 328350
rect 22478 328294 22546 328350
rect 22602 328294 53142 328350
rect 53198 328294 53266 328350
rect 53322 328294 83862 328350
rect 83918 328294 83986 328350
rect 84042 328294 114582 328350
rect 114638 328294 114706 328350
rect 114762 328294 145302 328350
rect 145358 328294 145426 328350
rect 145482 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 178518 328350
rect 178574 328294 178642 328350
rect 178698 328294 209238 328350
rect 209294 328294 209362 328350
rect 209418 328294 239958 328350
rect 240014 328294 240082 328350
rect 240138 328294 270678 328350
rect 270734 328294 270802 328350
rect 270858 328294 301398 328350
rect 301454 328294 301522 328350
rect 301578 328294 332118 328350
rect 332174 328294 332242 328350
rect 332298 328294 362838 328350
rect 362894 328294 362962 328350
rect 363018 328294 393558 328350
rect 393614 328294 393682 328350
rect 393738 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 448518 328350
rect 448574 328294 448642 328350
rect 448698 328294 479238 328350
rect 479294 328294 479362 328350
rect 479418 328294 509958 328350
rect 510014 328294 510082 328350
rect 510138 328294 540678 328350
rect 540734 328294 540802 328350
rect 540858 328294 571398 328350
rect 571454 328294 571522 328350
rect 571578 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 22422 328226
rect 22478 328170 22546 328226
rect 22602 328170 53142 328226
rect 53198 328170 53266 328226
rect 53322 328170 83862 328226
rect 83918 328170 83986 328226
rect 84042 328170 114582 328226
rect 114638 328170 114706 328226
rect 114762 328170 145302 328226
rect 145358 328170 145426 328226
rect 145482 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 178518 328226
rect 178574 328170 178642 328226
rect 178698 328170 209238 328226
rect 209294 328170 209362 328226
rect 209418 328170 239958 328226
rect 240014 328170 240082 328226
rect 240138 328170 270678 328226
rect 270734 328170 270802 328226
rect 270858 328170 301398 328226
rect 301454 328170 301522 328226
rect 301578 328170 332118 328226
rect 332174 328170 332242 328226
rect 332298 328170 362838 328226
rect 362894 328170 362962 328226
rect 363018 328170 393558 328226
rect 393614 328170 393682 328226
rect 393738 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 448518 328226
rect 448574 328170 448642 328226
rect 448698 328170 479238 328226
rect 479294 328170 479362 328226
rect 479418 328170 509958 328226
rect 510014 328170 510082 328226
rect 510138 328170 540678 328226
rect 540734 328170 540802 328226
rect 540858 328170 571398 328226
rect 571454 328170 571522 328226
rect 571578 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 22422 328102
rect 22478 328046 22546 328102
rect 22602 328046 53142 328102
rect 53198 328046 53266 328102
rect 53322 328046 83862 328102
rect 83918 328046 83986 328102
rect 84042 328046 114582 328102
rect 114638 328046 114706 328102
rect 114762 328046 145302 328102
rect 145358 328046 145426 328102
rect 145482 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 178518 328102
rect 178574 328046 178642 328102
rect 178698 328046 209238 328102
rect 209294 328046 209362 328102
rect 209418 328046 239958 328102
rect 240014 328046 240082 328102
rect 240138 328046 270678 328102
rect 270734 328046 270802 328102
rect 270858 328046 301398 328102
rect 301454 328046 301522 328102
rect 301578 328046 332118 328102
rect 332174 328046 332242 328102
rect 332298 328046 362838 328102
rect 362894 328046 362962 328102
rect 363018 328046 393558 328102
rect 393614 328046 393682 328102
rect 393738 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 448518 328102
rect 448574 328046 448642 328102
rect 448698 328046 479238 328102
rect 479294 328046 479362 328102
rect 479418 328046 509958 328102
rect 510014 328046 510082 328102
rect 510138 328046 540678 328102
rect 540734 328046 540802 328102
rect 540858 328046 571398 328102
rect 571454 328046 571522 328102
rect 571578 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 22422 327978
rect 22478 327922 22546 327978
rect 22602 327922 53142 327978
rect 53198 327922 53266 327978
rect 53322 327922 83862 327978
rect 83918 327922 83986 327978
rect 84042 327922 114582 327978
rect 114638 327922 114706 327978
rect 114762 327922 145302 327978
rect 145358 327922 145426 327978
rect 145482 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 178518 327978
rect 178574 327922 178642 327978
rect 178698 327922 209238 327978
rect 209294 327922 209362 327978
rect 209418 327922 239958 327978
rect 240014 327922 240082 327978
rect 240138 327922 270678 327978
rect 270734 327922 270802 327978
rect 270858 327922 301398 327978
rect 301454 327922 301522 327978
rect 301578 327922 332118 327978
rect 332174 327922 332242 327978
rect 332298 327922 362838 327978
rect 362894 327922 362962 327978
rect 363018 327922 393558 327978
rect 393614 327922 393682 327978
rect 393738 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 448518 327978
rect 448574 327922 448642 327978
rect 448698 327922 479238 327978
rect 479294 327922 479362 327978
rect 479418 327922 509958 327978
rect 510014 327922 510082 327978
rect 510138 327922 540678 327978
rect 540734 327922 540802 327978
rect 540858 327922 571398 327978
rect 571454 327922 571522 327978
rect 571578 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 37782 316350
rect 37838 316294 37906 316350
rect 37962 316294 68502 316350
rect 68558 316294 68626 316350
rect 68682 316294 99222 316350
rect 99278 316294 99346 316350
rect 99402 316294 129942 316350
rect 129998 316294 130066 316350
rect 130122 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 193878 316350
rect 193934 316294 194002 316350
rect 194058 316294 224598 316350
rect 224654 316294 224722 316350
rect 224778 316294 255318 316350
rect 255374 316294 255442 316350
rect 255498 316294 286038 316350
rect 286094 316294 286162 316350
rect 286218 316294 316758 316350
rect 316814 316294 316882 316350
rect 316938 316294 347478 316350
rect 347534 316294 347602 316350
rect 347658 316294 378198 316350
rect 378254 316294 378322 316350
rect 378378 316294 408918 316350
rect 408974 316294 409042 316350
rect 409098 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 463878 316350
rect 463934 316294 464002 316350
rect 464058 316294 494598 316350
rect 494654 316294 494722 316350
rect 494778 316294 525318 316350
rect 525374 316294 525442 316350
rect 525498 316294 556038 316350
rect 556094 316294 556162 316350
rect 556218 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 37782 316226
rect 37838 316170 37906 316226
rect 37962 316170 68502 316226
rect 68558 316170 68626 316226
rect 68682 316170 99222 316226
rect 99278 316170 99346 316226
rect 99402 316170 129942 316226
rect 129998 316170 130066 316226
rect 130122 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 193878 316226
rect 193934 316170 194002 316226
rect 194058 316170 224598 316226
rect 224654 316170 224722 316226
rect 224778 316170 255318 316226
rect 255374 316170 255442 316226
rect 255498 316170 286038 316226
rect 286094 316170 286162 316226
rect 286218 316170 316758 316226
rect 316814 316170 316882 316226
rect 316938 316170 347478 316226
rect 347534 316170 347602 316226
rect 347658 316170 378198 316226
rect 378254 316170 378322 316226
rect 378378 316170 408918 316226
rect 408974 316170 409042 316226
rect 409098 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 463878 316226
rect 463934 316170 464002 316226
rect 464058 316170 494598 316226
rect 494654 316170 494722 316226
rect 494778 316170 525318 316226
rect 525374 316170 525442 316226
rect 525498 316170 556038 316226
rect 556094 316170 556162 316226
rect 556218 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 37782 316102
rect 37838 316046 37906 316102
rect 37962 316046 68502 316102
rect 68558 316046 68626 316102
rect 68682 316046 99222 316102
rect 99278 316046 99346 316102
rect 99402 316046 129942 316102
rect 129998 316046 130066 316102
rect 130122 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 193878 316102
rect 193934 316046 194002 316102
rect 194058 316046 224598 316102
rect 224654 316046 224722 316102
rect 224778 316046 255318 316102
rect 255374 316046 255442 316102
rect 255498 316046 286038 316102
rect 286094 316046 286162 316102
rect 286218 316046 316758 316102
rect 316814 316046 316882 316102
rect 316938 316046 347478 316102
rect 347534 316046 347602 316102
rect 347658 316046 378198 316102
rect 378254 316046 378322 316102
rect 378378 316046 408918 316102
rect 408974 316046 409042 316102
rect 409098 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 463878 316102
rect 463934 316046 464002 316102
rect 464058 316046 494598 316102
rect 494654 316046 494722 316102
rect 494778 316046 525318 316102
rect 525374 316046 525442 316102
rect 525498 316046 556038 316102
rect 556094 316046 556162 316102
rect 556218 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 37782 315978
rect 37838 315922 37906 315978
rect 37962 315922 68502 315978
rect 68558 315922 68626 315978
rect 68682 315922 99222 315978
rect 99278 315922 99346 315978
rect 99402 315922 129942 315978
rect 129998 315922 130066 315978
rect 130122 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 193878 315978
rect 193934 315922 194002 315978
rect 194058 315922 224598 315978
rect 224654 315922 224722 315978
rect 224778 315922 255318 315978
rect 255374 315922 255442 315978
rect 255498 315922 286038 315978
rect 286094 315922 286162 315978
rect 286218 315922 316758 315978
rect 316814 315922 316882 315978
rect 316938 315922 347478 315978
rect 347534 315922 347602 315978
rect 347658 315922 378198 315978
rect 378254 315922 378322 315978
rect 378378 315922 408918 315978
rect 408974 315922 409042 315978
rect 409098 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 463878 315978
rect 463934 315922 464002 315978
rect 464058 315922 494598 315978
rect 494654 315922 494722 315978
rect 494778 315922 525318 315978
rect 525374 315922 525442 315978
rect 525498 315922 556038 315978
rect 556094 315922 556162 315978
rect 556218 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 22422 310350
rect 22478 310294 22546 310350
rect 22602 310294 53142 310350
rect 53198 310294 53266 310350
rect 53322 310294 83862 310350
rect 83918 310294 83986 310350
rect 84042 310294 114582 310350
rect 114638 310294 114706 310350
rect 114762 310294 145302 310350
rect 145358 310294 145426 310350
rect 145482 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 448518 310350
rect 448574 310294 448642 310350
rect 448698 310294 479238 310350
rect 479294 310294 479362 310350
rect 479418 310294 509958 310350
rect 510014 310294 510082 310350
rect 510138 310294 540678 310350
rect 540734 310294 540802 310350
rect 540858 310294 571398 310350
rect 571454 310294 571522 310350
rect 571578 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 22422 310226
rect 22478 310170 22546 310226
rect 22602 310170 53142 310226
rect 53198 310170 53266 310226
rect 53322 310170 83862 310226
rect 83918 310170 83986 310226
rect 84042 310170 114582 310226
rect 114638 310170 114706 310226
rect 114762 310170 145302 310226
rect 145358 310170 145426 310226
rect 145482 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 448518 310226
rect 448574 310170 448642 310226
rect 448698 310170 479238 310226
rect 479294 310170 479362 310226
rect 479418 310170 509958 310226
rect 510014 310170 510082 310226
rect 510138 310170 540678 310226
rect 540734 310170 540802 310226
rect 540858 310170 571398 310226
rect 571454 310170 571522 310226
rect 571578 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 22422 310102
rect 22478 310046 22546 310102
rect 22602 310046 53142 310102
rect 53198 310046 53266 310102
rect 53322 310046 83862 310102
rect 83918 310046 83986 310102
rect 84042 310046 114582 310102
rect 114638 310046 114706 310102
rect 114762 310046 145302 310102
rect 145358 310046 145426 310102
rect 145482 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 448518 310102
rect 448574 310046 448642 310102
rect 448698 310046 479238 310102
rect 479294 310046 479362 310102
rect 479418 310046 509958 310102
rect 510014 310046 510082 310102
rect 510138 310046 540678 310102
rect 540734 310046 540802 310102
rect 540858 310046 571398 310102
rect 571454 310046 571522 310102
rect 571578 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 22422 309978
rect 22478 309922 22546 309978
rect 22602 309922 53142 309978
rect 53198 309922 53266 309978
rect 53322 309922 83862 309978
rect 83918 309922 83986 309978
rect 84042 309922 114582 309978
rect 114638 309922 114706 309978
rect 114762 309922 145302 309978
rect 145358 309922 145426 309978
rect 145482 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 448518 309978
rect 448574 309922 448642 309978
rect 448698 309922 479238 309978
rect 479294 309922 479362 309978
rect 479418 309922 509958 309978
rect 510014 309922 510082 309978
rect 510138 309922 540678 309978
rect 540734 309922 540802 309978
rect 540858 309922 571398 309978
rect 571454 309922 571522 309978
rect 571578 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect 310812 305038 327812 305054
rect 310812 304982 310828 305038
rect 310884 304982 327740 305038
rect 327796 304982 327812 305038
rect 310812 304966 327812 304982
rect 336460 305038 355924 305054
rect 336460 304982 336476 305038
rect 336532 304982 355852 305038
rect 355908 304982 355924 305038
rect 336460 304966 355924 304982
rect 324140 304858 344724 304874
rect 324140 304802 324156 304858
rect 324212 304802 344652 304858
rect 344708 304802 344724 304858
rect 324140 304786 344724 304802
rect 357740 304858 376532 304874
rect 357740 304802 357756 304858
rect 357812 304802 376460 304858
rect 376516 304802 376532 304858
rect 357740 304786 376532 304802
rect 381036 304858 401620 304874
rect 381036 304802 381052 304858
rect 381108 304802 401548 304858
rect 401604 304802 401620 304858
rect 381036 304786 401620 304802
rect 342508 304318 357828 304334
rect 342508 304262 342524 304318
rect 342580 304262 357756 304318
rect 357812 304262 357828 304318
rect 342508 304246 357828 304262
rect 173836 304138 272260 304154
rect 173836 304082 173852 304138
rect 173908 304082 272188 304138
rect 272244 304082 272260 304138
rect 173836 304066 272260 304082
rect 330412 304138 351444 304154
rect 330412 304082 330428 304138
rect 330484 304082 351372 304138
rect 351428 304082 351444 304138
rect 330412 304066 351444 304082
rect 352364 304138 372500 304154
rect 352364 304082 352380 304138
rect 352436 304082 372428 304138
rect 372484 304082 372500 304138
rect 352364 304066 372500 304082
rect 342956 303958 363540 303974
rect 342956 303902 342972 303958
rect 343028 303902 363468 303958
rect 363524 303902 363540 303958
rect 342956 303886 363540 303902
rect 369388 303958 389972 303974
rect 369388 303902 369404 303958
rect 369460 303902 389900 303958
rect 389956 303902 389972 303958
rect 369388 303886 389972 303902
rect 330860 303778 347860 303794
rect 330860 303722 330876 303778
rect 330932 303722 347788 303778
rect 347844 303722 347860 303778
rect 330860 303706 347860 303722
rect 379580 303778 398484 303794
rect 379580 303722 379596 303778
rect 379652 303722 398412 303778
rect 398468 303722 398484 303778
rect 379580 303706 398484 303722
rect 336012 303598 351108 303614
rect 336012 303542 336028 303598
rect 336084 303542 351036 303598
rect 351092 303542 351108 303598
rect 336012 303526 351108 303542
rect 360876 303598 381460 303614
rect 360876 303542 360892 303598
rect 360948 303542 381388 303598
rect 381444 303542 381460 303598
rect 360876 303526 381460 303542
rect 324588 303418 342708 303434
rect 324588 303362 324604 303418
rect 324660 303362 342636 303418
rect 342692 303362 342708 303418
rect 324588 303346 342708 303362
rect 309132 303238 324564 303254
rect 309132 303182 309148 303238
rect 309204 303182 324492 303238
rect 324548 303182 324564 303238
rect 309132 303166 324564 303182
rect 327276 303238 344500 303254
rect 327276 303182 327292 303238
rect 327348 303182 344428 303238
rect 344484 303182 344500 303238
rect 327276 303166 344500 303182
rect 362668 303238 379780 303254
rect 362668 303182 362684 303238
rect 362740 303182 379708 303238
rect 379764 303182 379780 303238
rect 362668 303166 379780 303182
rect 394476 303238 415060 303254
rect 394476 303182 394492 303238
rect 394548 303182 414988 303238
rect 415044 303182 415060 303238
rect 394476 303166 415060 303182
rect 318988 302518 332628 302534
rect 318988 302462 319004 302518
rect 319060 302462 332556 302518
rect 332612 302462 332628 302518
rect 318988 302446 332628 302462
rect 320780 302338 329940 302354
rect 320780 302282 320796 302338
rect 320852 302282 329868 302338
rect 329924 302282 329940 302338
rect 320780 302266 329940 302282
rect 364572 302338 374628 302354
rect 364572 302282 364588 302338
rect 364644 302282 374556 302338
rect 374612 302282 374628 302338
rect 364572 302266 374628 302282
rect 320668 302158 329492 302174
rect 320668 302102 320684 302158
rect 320740 302102 329420 302158
rect 329476 302102 329492 302158
rect 320668 302086 329492 302102
rect 393132 302158 399828 302174
rect 393132 302102 393148 302158
rect 393204 302102 399756 302158
rect 399812 302102 399828 302158
rect 393132 302086 399828 302102
rect 374316 301798 394900 301814
rect 374316 301742 374332 301798
rect 374388 301742 394828 301798
rect 394884 301742 394900 301798
rect 374316 301726 394900 301742
rect 228716 301618 315156 301634
rect 228716 301562 228732 301618
rect 228788 301562 315084 301618
rect 315140 301562 315156 301618
rect 228716 301546 315156 301562
rect 344300 301618 364884 301634
rect 344300 301562 344316 301618
rect 344372 301562 364812 301618
rect 364868 301562 364884 301618
rect 344300 301546 364884 301562
rect 367596 301618 388180 301634
rect 367596 301562 367612 301618
rect 367668 301562 388108 301618
rect 388164 301562 388180 301618
rect 367596 301546 388180 301562
rect 229164 301438 318404 301454
rect 229164 301382 229180 301438
rect 229236 301382 318332 301438
rect 318388 301382 318404 301438
rect 229164 301366 318404 301382
rect 218412 301258 310676 301274
rect 218412 301202 218428 301258
rect 218484 301202 310604 301258
rect 310660 301202 310676 301258
rect 218412 301186 310676 301202
rect 310812 301258 434436 301274
rect 310812 301202 310828 301258
rect 310884 301202 434364 301258
rect 434420 301202 434436 301258
rect 310812 301186 434436 301202
rect 260524 301078 423572 301094
rect 260524 301022 260540 301078
rect 260596 301022 423500 301078
rect 423556 301022 423572 301078
rect 260524 301006 423572 301022
rect 242156 300898 437908 300914
rect 242156 300842 242172 300898
rect 242228 300842 437836 300898
rect 437892 300842 437908 300898
rect 242156 300826 437908 300842
rect 237676 300178 442836 300194
rect 237676 300122 237692 300178
rect 237748 300122 442764 300178
rect 442820 300122 442836 300178
rect 237676 300106 442836 300122
rect 217964 299998 431860 300014
rect 217964 299942 217980 299998
rect 218036 299942 431788 299998
rect 431844 299942 431860 299998
rect 217964 299926 431860 299942
rect 223340 299818 436900 299834
rect 223340 299762 223356 299818
rect 223412 299762 436828 299818
rect 436884 299762 436900 299818
rect 223340 299746 436900 299762
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 37782 298350
rect 37838 298294 37906 298350
rect 37962 298294 68502 298350
rect 68558 298294 68626 298350
rect 68682 298294 99222 298350
rect 99278 298294 99346 298350
rect 99402 298294 129942 298350
rect 129998 298294 130066 298350
rect 130122 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 285714 298350
rect 285770 298294 285838 298350
rect 285894 298294 285962 298350
rect 286018 298294 286086 298350
rect 286142 298294 316434 298350
rect 316490 298294 316558 298350
rect 316614 298294 316682 298350
rect 316738 298294 316806 298350
rect 316862 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 463878 298350
rect 463934 298294 464002 298350
rect 464058 298294 494598 298350
rect 494654 298294 494722 298350
rect 494778 298294 525318 298350
rect 525374 298294 525442 298350
rect 525498 298294 556038 298350
rect 556094 298294 556162 298350
rect 556218 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 37782 298226
rect 37838 298170 37906 298226
rect 37962 298170 68502 298226
rect 68558 298170 68626 298226
rect 68682 298170 99222 298226
rect 99278 298170 99346 298226
rect 99402 298170 129942 298226
rect 129998 298170 130066 298226
rect 130122 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 285714 298226
rect 285770 298170 285838 298226
rect 285894 298170 285962 298226
rect 286018 298170 286086 298226
rect 286142 298170 316434 298226
rect 316490 298170 316558 298226
rect 316614 298170 316682 298226
rect 316738 298170 316806 298226
rect 316862 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 463878 298226
rect 463934 298170 464002 298226
rect 464058 298170 494598 298226
rect 494654 298170 494722 298226
rect 494778 298170 525318 298226
rect 525374 298170 525442 298226
rect 525498 298170 556038 298226
rect 556094 298170 556162 298226
rect 556218 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 37782 298102
rect 37838 298046 37906 298102
rect 37962 298046 68502 298102
rect 68558 298046 68626 298102
rect 68682 298046 99222 298102
rect 99278 298046 99346 298102
rect 99402 298046 129942 298102
rect 129998 298046 130066 298102
rect 130122 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 285714 298102
rect 285770 298046 285838 298102
rect 285894 298046 285962 298102
rect 286018 298046 286086 298102
rect 286142 298046 316434 298102
rect 316490 298046 316558 298102
rect 316614 298046 316682 298102
rect 316738 298046 316806 298102
rect 316862 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 463878 298102
rect 463934 298046 464002 298102
rect 464058 298046 494598 298102
rect 494654 298046 494722 298102
rect 494778 298046 525318 298102
rect 525374 298046 525442 298102
rect 525498 298046 556038 298102
rect 556094 298046 556162 298102
rect 556218 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 37782 297978
rect 37838 297922 37906 297978
rect 37962 297922 68502 297978
rect 68558 297922 68626 297978
rect 68682 297922 99222 297978
rect 99278 297922 99346 297978
rect 99402 297922 129942 297978
rect 129998 297922 130066 297978
rect 130122 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 285714 297978
rect 285770 297922 285838 297978
rect 285894 297922 285962 297978
rect 286018 297922 286086 297978
rect 286142 297922 316434 297978
rect 316490 297922 316558 297978
rect 316614 297922 316682 297978
rect 316738 297922 316806 297978
rect 316862 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 463878 297978
rect 463934 297922 464002 297978
rect 464058 297922 494598 297978
rect 494654 297922 494722 297978
rect 494778 297922 525318 297978
rect 525374 297922 525442 297978
rect 525498 297922 556038 297978
rect 556094 297922 556162 297978
rect 556218 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 22422 292350
rect 22478 292294 22546 292350
rect 22602 292294 53142 292350
rect 53198 292294 53266 292350
rect 53322 292294 83862 292350
rect 83918 292294 83986 292350
rect 84042 292294 114582 292350
rect 114638 292294 114706 292350
rect 114762 292294 145302 292350
rect 145358 292294 145426 292350
rect 145482 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 178518 292350
rect 178574 292294 178642 292350
rect 178698 292294 209238 292350
rect 209294 292294 209362 292350
rect 209418 292294 239958 292350
rect 240014 292294 240082 292350
rect 240138 292294 270678 292350
rect 270734 292294 270802 292350
rect 270858 292294 281994 292350
rect 282050 292294 282118 292350
rect 282174 292294 282242 292350
rect 282298 292294 282366 292350
rect 282422 292294 312714 292350
rect 312770 292294 312838 292350
rect 312894 292294 312962 292350
rect 313018 292294 313086 292350
rect 313142 292294 324518 292350
rect 324574 292294 324642 292350
rect 324698 292294 355238 292350
rect 355294 292294 355362 292350
rect 355418 292294 385958 292350
rect 386014 292294 386082 292350
rect 386138 292294 416678 292350
rect 416734 292294 416802 292350
rect 416858 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 448518 292350
rect 448574 292294 448642 292350
rect 448698 292294 479238 292350
rect 479294 292294 479362 292350
rect 479418 292294 509958 292350
rect 510014 292294 510082 292350
rect 510138 292294 540678 292350
rect 540734 292294 540802 292350
rect 540858 292294 571398 292350
rect 571454 292294 571522 292350
rect 571578 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 22422 292226
rect 22478 292170 22546 292226
rect 22602 292170 53142 292226
rect 53198 292170 53266 292226
rect 53322 292170 83862 292226
rect 83918 292170 83986 292226
rect 84042 292170 114582 292226
rect 114638 292170 114706 292226
rect 114762 292170 145302 292226
rect 145358 292170 145426 292226
rect 145482 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 178518 292226
rect 178574 292170 178642 292226
rect 178698 292170 209238 292226
rect 209294 292170 209362 292226
rect 209418 292170 239958 292226
rect 240014 292170 240082 292226
rect 240138 292170 270678 292226
rect 270734 292170 270802 292226
rect 270858 292170 281994 292226
rect 282050 292170 282118 292226
rect 282174 292170 282242 292226
rect 282298 292170 282366 292226
rect 282422 292170 312714 292226
rect 312770 292170 312838 292226
rect 312894 292170 312962 292226
rect 313018 292170 313086 292226
rect 313142 292170 324518 292226
rect 324574 292170 324642 292226
rect 324698 292170 355238 292226
rect 355294 292170 355362 292226
rect 355418 292170 385958 292226
rect 386014 292170 386082 292226
rect 386138 292170 416678 292226
rect 416734 292170 416802 292226
rect 416858 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 448518 292226
rect 448574 292170 448642 292226
rect 448698 292170 479238 292226
rect 479294 292170 479362 292226
rect 479418 292170 509958 292226
rect 510014 292170 510082 292226
rect 510138 292170 540678 292226
rect 540734 292170 540802 292226
rect 540858 292170 571398 292226
rect 571454 292170 571522 292226
rect 571578 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 22422 292102
rect 22478 292046 22546 292102
rect 22602 292046 53142 292102
rect 53198 292046 53266 292102
rect 53322 292046 83862 292102
rect 83918 292046 83986 292102
rect 84042 292046 114582 292102
rect 114638 292046 114706 292102
rect 114762 292046 145302 292102
rect 145358 292046 145426 292102
rect 145482 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 178518 292102
rect 178574 292046 178642 292102
rect 178698 292046 209238 292102
rect 209294 292046 209362 292102
rect 209418 292046 239958 292102
rect 240014 292046 240082 292102
rect 240138 292046 270678 292102
rect 270734 292046 270802 292102
rect 270858 292046 281994 292102
rect 282050 292046 282118 292102
rect 282174 292046 282242 292102
rect 282298 292046 282366 292102
rect 282422 292046 312714 292102
rect 312770 292046 312838 292102
rect 312894 292046 312962 292102
rect 313018 292046 313086 292102
rect 313142 292046 324518 292102
rect 324574 292046 324642 292102
rect 324698 292046 355238 292102
rect 355294 292046 355362 292102
rect 355418 292046 385958 292102
rect 386014 292046 386082 292102
rect 386138 292046 416678 292102
rect 416734 292046 416802 292102
rect 416858 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 448518 292102
rect 448574 292046 448642 292102
rect 448698 292046 479238 292102
rect 479294 292046 479362 292102
rect 479418 292046 509958 292102
rect 510014 292046 510082 292102
rect 510138 292046 540678 292102
rect 540734 292046 540802 292102
rect 540858 292046 571398 292102
rect 571454 292046 571522 292102
rect 571578 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 22422 291978
rect 22478 291922 22546 291978
rect 22602 291922 53142 291978
rect 53198 291922 53266 291978
rect 53322 291922 83862 291978
rect 83918 291922 83986 291978
rect 84042 291922 114582 291978
rect 114638 291922 114706 291978
rect 114762 291922 145302 291978
rect 145358 291922 145426 291978
rect 145482 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 178518 291978
rect 178574 291922 178642 291978
rect 178698 291922 209238 291978
rect 209294 291922 209362 291978
rect 209418 291922 239958 291978
rect 240014 291922 240082 291978
rect 240138 291922 270678 291978
rect 270734 291922 270802 291978
rect 270858 291922 281994 291978
rect 282050 291922 282118 291978
rect 282174 291922 282242 291978
rect 282298 291922 282366 291978
rect 282422 291922 312714 291978
rect 312770 291922 312838 291978
rect 312894 291922 312962 291978
rect 313018 291922 313086 291978
rect 313142 291922 324518 291978
rect 324574 291922 324642 291978
rect 324698 291922 355238 291978
rect 355294 291922 355362 291978
rect 355418 291922 385958 291978
rect 386014 291922 386082 291978
rect 386138 291922 416678 291978
rect 416734 291922 416802 291978
rect 416858 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 448518 291978
rect 448574 291922 448642 291978
rect 448698 291922 479238 291978
rect 479294 291922 479362 291978
rect 479418 291922 509958 291978
rect 510014 291922 510082 291978
rect 510138 291922 540678 291978
rect 540734 291922 540802 291978
rect 540858 291922 571398 291978
rect 571454 291922 571522 291978
rect 571578 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 37782 280350
rect 37838 280294 37906 280350
rect 37962 280294 68502 280350
rect 68558 280294 68626 280350
rect 68682 280294 99222 280350
rect 99278 280294 99346 280350
rect 99402 280294 129942 280350
rect 129998 280294 130066 280350
rect 130122 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 193878 280350
rect 193934 280294 194002 280350
rect 194058 280294 224598 280350
rect 224654 280294 224722 280350
rect 224778 280294 255318 280350
rect 255374 280294 255442 280350
rect 255498 280294 285714 280350
rect 285770 280294 285838 280350
rect 285894 280294 285962 280350
rect 286018 280294 286086 280350
rect 286142 280294 316434 280350
rect 316490 280294 316558 280350
rect 316614 280294 316682 280350
rect 316738 280294 316806 280350
rect 316862 280294 339878 280350
rect 339934 280294 340002 280350
rect 340058 280294 370598 280350
rect 370654 280294 370722 280350
rect 370778 280294 401318 280350
rect 401374 280294 401442 280350
rect 401498 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 463878 280350
rect 463934 280294 464002 280350
rect 464058 280294 494598 280350
rect 494654 280294 494722 280350
rect 494778 280294 525318 280350
rect 525374 280294 525442 280350
rect 525498 280294 556038 280350
rect 556094 280294 556162 280350
rect 556218 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 37782 280226
rect 37838 280170 37906 280226
rect 37962 280170 68502 280226
rect 68558 280170 68626 280226
rect 68682 280170 99222 280226
rect 99278 280170 99346 280226
rect 99402 280170 129942 280226
rect 129998 280170 130066 280226
rect 130122 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 193878 280226
rect 193934 280170 194002 280226
rect 194058 280170 224598 280226
rect 224654 280170 224722 280226
rect 224778 280170 255318 280226
rect 255374 280170 255442 280226
rect 255498 280170 285714 280226
rect 285770 280170 285838 280226
rect 285894 280170 285962 280226
rect 286018 280170 286086 280226
rect 286142 280170 316434 280226
rect 316490 280170 316558 280226
rect 316614 280170 316682 280226
rect 316738 280170 316806 280226
rect 316862 280170 339878 280226
rect 339934 280170 340002 280226
rect 340058 280170 370598 280226
rect 370654 280170 370722 280226
rect 370778 280170 401318 280226
rect 401374 280170 401442 280226
rect 401498 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 463878 280226
rect 463934 280170 464002 280226
rect 464058 280170 494598 280226
rect 494654 280170 494722 280226
rect 494778 280170 525318 280226
rect 525374 280170 525442 280226
rect 525498 280170 556038 280226
rect 556094 280170 556162 280226
rect 556218 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 37782 280102
rect 37838 280046 37906 280102
rect 37962 280046 68502 280102
rect 68558 280046 68626 280102
rect 68682 280046 99222 280102
rect 99278 280046 99346 280102
rect 99402 280046 129942 280102
rect 129998 280046 130066 280102
rect 130122 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 193878 280102
rect 193934 280046 194002 280102
rect 194058 280046 224598 280102
rect 224654 280046 224722 280102
rect 224778 280046 255318 280102
rect 255374 280046 255442 280102
rect 255498 280046 285714 280102
rect 285770 280046 285838 280102
rect 285894 280046 285962 280102
rect 286018 280046 286086 280102
rect 286142 280046 316434 280102
rect 316490 280046 316558 280102
rect 316614 280046 316682 280102
rect 316738 280046 316806 280102
rect 316862 280046 339878 280102
rect 339934 280046 340002 280102
rect 340058 280046 370598 280102
rect 370654 280046 370722 280102
rect 370778 280046 401318 280102
rect 401374 280046 401442 280102
rect 401498 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 463878 280102
rect 463934 280046 464002 280102
rect 464058 280046 494598 280102
rect 494654 280046 494722 280102
rect 494778 280046 525318 280102
rect 525374 280046 525442 280102
rect 525498 280046 556038 280102
rect 556094 280046 556162 280102
rect 556218 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 37782 279978
rect 37838 279922 37906 279978
rect 37962 279922 68502 279978
rect 68558 279922 68626 279978
rect 68682 279922 99222 279978
rect 99278 279922 99346 279978
rect 99402 279922 129942 279978
rect 129998 279922 130066 279978
rect 130122 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 193878 279978
rect 193934 279922 194002 279978
rect 194058 279922 224598 279978
rect 224654 279922 224722 279978
rect 224778 279922 255318 279978
rect 255374 279922 255442 279978
rect 255498 279922 285714 279978
rect 285770 279922 285838 279978
rect 285894 279922 285962 279978
rect 286018 279922 286086 279978
rect 286142 279922 316434 279978
rect 316490 279922 316558 279978
rect 316614 279922 316682 279978
rect 316738 279922 316806 279978
rect 316862 279922 339878 279978
rect 339934 279922 340002 279978
rect 340058 279922 370598 279978
rect 370654 279922 370722 279978
rect 370778 279922 401318 279978
rect 401374 279922 401442 279978
rect 401498 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 463878 279978
rect 463934 279922 464002 279978
rect 464058 279922 494598 279978
rect 494654 279922 494722 279978
rect 494778 279922 525318 279978
rect 525374 279922 525442 279978
rect 525498 279922 556038 279978
rect 556094 279922 556162 279978
rect 556218 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 22422 274350
rect 22478 274294 22546 274350
rect 22602 274294 53142 274350
rect 53198 274294 53266 274350
rect 53322 274294 83862 274350
rect 83918 274294 83986 274350
rect 84042 274294 114582 274350
rect 114638 274294 114706 274350
rect 114762 274294 145302 274350
rect 145358 274294 145426 274350
rect 145482 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 178518 274350
rect 178574 274294 178642 274350
rect 178698 274294 209238 274350
rect 209294 274294 209362 274350
rect 209418 274294 239958 274350
rect 240014 274294 240082 274350
rect 240138 274294 270678 274350
rect 270734 274294 270802 274350
rect 270858 274294 281994 274350
rect 282050 274294 282118 274350
rect 282174 274294 282242 274350
rect 282298 274294 282366 274350
rect 282422 274294 312714 274350
rect 312770 274294 312838 274350
rect 312894 274294 312962 274350
rect 313018 274294 313086 274350
rect 313142 274294 324518 274350
rect 324574 274294 324642 274350
rect 324698 274294 355238 274350
rect 355294 274294 355362 274350
rect 355418 274294 385958 274350
rect 386014 274294 386082 274350
rect 386138 274294 416678 274350
rect 416734 274294 416802 274350
rect 416858 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 448518 274350
rect 448574 274294 448642 274350
rect 448698 274294 479238 274350
rect 479294 274294 479362 274350
rect 479418 274294 509958 274350
rect 510014 274294 510082 274350
rect 510138 274294 540678 274350
rect 540734 274294 540802 274350
rect 540858 274294 571398 274350
rect 571454 274294 571522 274350
rect 571578 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 22422 274226
rect 22478 274170 22546 274226
rect 22602 274170 53142 274226
rect 53198 274170 53266 274226
rect 53322 274170 83862 274226
rect 83918 274170 83986 274226
rect 84042 274170 114582 274226
rect 114638 274170 114706 274226
rect 114762 274170 145302 274226
rect 145358 274170 145426 274226
rect 145482 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 178518 274226
rect 178574 274170 178642 274226
rect 178698 274170 209238 274226
rect 209294 274170 209362 274226
rect 209418 274170 239958 274226
rect 240014 274170 240082 274226
rect 240138 274170 270678 274226
rect 270734 274170 270802 274226
rect 270858 274170 281994 274226
rect 282050 274170 282118 274226
rect 282174 274170 282242 274226
rect 282298 274170 282366 274226
rect 282422 274170 312714 274226
rect 312770 274170 312838 274226
rect 312894 274170 312962 274226
rect 313018 274170 313086 274226
rect 313142 274170 324518 274226
rect 324574 274170 324642 274226
rect 324698 274170 355238 274226
rect 355294 274170 355362 274226
rect 355418 274170 385958 274226
rect 386014 274170 386082 274226
rect 386138 274170 416678 274226
rect 416734 274170 416802 274226
rect 416858 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 448518 274226
rect 448574 274170 448642 274226
rect 448698 274170 479238 274226
rect 479294 274170 479362 274226
rect 479418 274170 509958 274226
rect 510014 274170 510082 274226
rect 510138 274170 540678 274226
rect 540734 274170 540802 274226
rect 540858 274170 571398 274226
rect 571454 274170 571522 274226
rect 571578 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 22422 274102
rect 22478 274046 22546 274102
rect 22602 274046 53142 274102
rect 53198 274046 53266 274102
rect 53322 274046 83862 274102
rect 83918 274046 83986 274102
rect 84042 274046 114582 274102
rect 114638 274046 114706 274102
rect 114762 274046 145302 274102
rect 145358 274046 145426 274102
rect 145482 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 178518 274102
rect 178574 274046 178642 274102
rect 178698 274046 209238 274102
rect 209294 274046 209362 274102
rect 209418 274046 239958 274102
rect 240014 274046 240082 274102
rect 240138 274046 270678 274102
rect 270734 274046 270802 274102
rect 270858 274046 281994 274102
rect 282050 274046 282118 274102
rect 282174 274046 282242 274102
rect 282298 274046 282366 274102
rect 282422 274046 312714 274102
rect 312770 274046 312838 274102
rect 312894 274046 312962 274102
rect 313018 274046 313086 274102
rect 313142 274046 324518 274102
rect 324574 274046 324642 274102
rect 324698 274046 355238 274102
rect 355294 274046 355362 274102
rect 355418 274046 385958 274102
rect 386014 274046 386082 274102
rect 386138 274046 416678 274102
rect 416734 274046 416802 274102
rect 416858 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 448518 274102
rect 448574 274046 448642 274102
rect 448698 274046 479238 274102
rect 479294 274046 479362 274102
rect 479418 274046 509958 274102
rect 510014 274046 510082 274102
rect 510138 274046 540678 274102
rect 540734 274046 540802 274102
rect 540858 274046 571398 274102
rect 571454 274046 571522 274102
rect 571578 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 22422 273978
rect 22478 273922 22546 273978
rect 22602 273922 53142 273978
rect 53198 273922 53266 273978
rect 53322 273922 83862 273978
rect 83918 273922 83986 273978
rect 84042 273922 114582 273978
rect 114638 273922 114706 273978
rect 114762 273922 145302 273978
rect 145358 273922 145426 273978
rect 145482 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 178518 273978
rect 178574 273922 178642 273978
rect 178698 273922 209238 273978
rect 209294 273922 209362 273978
rect 209418 273922 239958 273978
rect 240014 273922 240082 273978
rect 240138 273922 270678 273978
rect 270734 273922 270802 273978
rect 270858 273922 281994 273978
rect 282050 273922 282118 273978
rect 282174 273922 282242 273978
rect 282298 273922 282366 273978
rect 282422 273922 312714 273978
rect 312770 273922 312838 273978
rect 312894 273922 312962 273978
rect 313018 273922 313086 273978
rect 313142 273922 324518 273978
rect 324574 273922 324642 273978
rect 324698 273922 355238 273978
rect 355294 273922 355362 273978
rect 355418 273922 385958 273978
rect 386014 273922 386082 273978
rect 386138 273922 416678 273978
rect 416734 273922 416802 273978
rect 416858 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 448518 273978
rect 448574 273922 448642 273978
rect 448698 273922 479238 273978
rect 479294 273922 479362 273978
rect 479418 273922 509958 273978
rect 510014 273922 510082 273978
rect 510138 273922 540678 273978
rect 540734 273922 540802 273978
rect 540858 273922 571398 273978
rect 571454 273922 571522 273978
rect 571578 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 37782 262350
rect 37838 262294 37906 262350
rect 37962 262294 68502 262350
rect 68558 262294 68626 262350
rect 68682 262294 99222 262350
rect 99278 262294 99346 262350
rect 99402 262294 129942 262350
rect 129998 262294 130066 262350
rect 130122 262294 162834 262350
rect 162890 262294 162958 262350
rect 163014 262294 163082 262350
rect 163138 262294 163206 262350
rect 163262 262294 193878 262350
rect 193934 262294 194002 262350
rect 194058 262294 224598 262350
rect 224654 262294 224722 262350
rect 224778 262294 255318 262350
rect 255374 262294 255442 262350
rect 255498 262294 285714 262350
rect 285770 262294 285838 262350
rect 285894 262294 285962 262350
rect 286018 262294 286086 262350
rect 286142 262294 316434 262350
rect 316490 262294 316558 262350
rect 316614 262294 316682 262350
rect 316738 262294 316806 262350
rect 316862 262294 339878 262350
rect 339934 262294 340002 262350
rect 340058 262294 370598 262350
rect 370654 262294 370722 262350
rect 370778 262294 401318 262350
rect 401374 262294 401442 262350
rect 401498 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 463878 262350
rect 463934 262294 464002 262350
rect 464058 262294 494598 262350
rect 494654 262294 494722 262350
rect 494778 262294 525318 262350
rect 525374 262294 525442 262350
rect 525498 262294 556038 262350
rect 556094 262294 556162 262350
rect 556218 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 37782 262226
rect 37838 262170 37906 262226
rect 37962 262170 68502 262226
rect 68558 262170 68626 262226
rect 68682 262170 99222 262226
rect 99278 262170 99346 262226
rect 99402 262170 129942 262226
rect 129998 262170 130066 262226
rect 130122 262170 162834 262226
rect 162890 262170 162958 262226
rect 163014 262170 163082 262226
rect 163138 262170 163206 262226
rect 163262 262170 193878 262226
rect 193934 262170 194002 262226
rect 194058 262170 224598 262226
rect 224654 262170 224722 262226
rect 224778 262170 255318 262226
rect 255374 262170 255442 262226
rect 255498 262170 285714 262226
rect 285770 262170 285838 262226
rect 285894 262170 285962 262226
rect 286018 262170 286086 262226
rect 286142 262170 316434 262226
rect 316490 262170 316558 262226
rect 316614 262170 316682 262226
rect 316738 262170 316806 262226
rect 316862 262170 339878 262226
rect 339934 262170 340002 262226
rect 340058 262170 370598 262226
rect 370654 262170 370722 262226
rect 370778 262170 401318 262226
rect 401374 262170 401442 262226
rect 401498 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 463878 262226
rect 463934 262170 464002 262226
rect 464058 262170 494598 262226
rect 494654 262170 494722 262226
rect 494778 262170 525318 262226
rect 525374 262170 525442 262226
rect 525498 262170 556038 262226
rect 556094 262170 556162 262226
rect 556218 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 37782 262102
rect 37838 262046 37906 262102
rect 37962 262046 68502 262102
rect 68558 262046 68626 262102
rect 68682 262046 99222 262102
rect 99278 262046 99346 262102
rect 99402 262046 129942 262102
rect 129998 262046 130066 262102
rect 130122 262046 162834 262102
rect 162890 262046 162958 262102
rect 163014 262046 163082 262102
rect 163138 262046 163206 262102
rect 163262 262046 193878 262102
rect 193934 262046 194002 262102
rect 194058 262046 224598 262102
rect 224654 262046 224722 262102
rect 224778 262046 255318 262102
rect 255374 262046 255442 262102
rect 255498 262046 285714 262102
rect 285770 262046 285838 262102
rect 285894 262046 285962 262102
rect 286018 262046 286086 262102
rect 286142 262046 316434 262102
rect 316490 262046 316558 262102
rect 316614 262046 316682 262102
rect 316738 262046 316806 262102
rect 316862 262046 339878 262102
rect 339934 262046 340002 262102
rect 340058 262046 370598 262102
rect 370654 262046 370722 262102
rect 370778 262046 401318 262102
rect 401374 262046 401442 262102
rect 401498 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 463878 262102
rect 463934 262046 464002 262102
rect 464058 262046 494598 262102
rect 494654 262046 494722 262102
rect 494778 262046 525318 262102
rect 525374 262046 525442 262102
rect 525498 262046 556038 262102
rect 556094 262046 556162 262102
rect 556218 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 37782 261978
rect 37838 261922 37906 261978
rect 37962 261922 68502 261978
rect 68558 261922 68626 261978
rect 68682 261922 99222 261978
rect 99278 261922 99346 261978
rect 99402 261922 129942 261978
rect 129998 261922 130066 261978
rect 130122 261922 162834 261978
rect 162890 261922 162958 261978
rect 163014 261922 163082 261978
rect 163138 261922 163206 261978
rect 163262 261922 193878 261978
rect 193934 261922 194002 261978
rect 194058 261922 224598 261978
rect 224654 261922 224722 261978
rect 224778 261922 255318 261978
rect 255374 261922 255442 261978
rect 255498 261922 285714 261978
rect 285770 261922 285838 261978
rect 285894 261922 285962 261978
rect 286018 261922 286086 261978
rect 286142 261922 316434 261978
rect 316490 261922 316558 261978
rect 316614 261922 316682 261978
rect 316738 261922 316806 261978
rect 316862 261922 339878 261978
rect 339934 261922 340002 261978
rect 340058 261922 370598 261978
rect 370654 261922 370722 261978
rect 370778 261922 401318 261978
rect 401374 261922 401442 261978
rect 401498 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 463878 261978
rect 463934 261922 464002 261978
rect 464058 261922 494598 261978
rect 494654 261922 494722 261978
rect 494778 261922 525318 261978
rect 525374 261922 525442 261978
rect 525498 261922 556038 261978
rect 556094 261922 556162 261978
rect 556218 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 22422 256350
rect 22478 256294 22546 256350
rect 22602 256294 53142 256350
rect 53198 256294 53266 256350
rect 53322 256294 83862 256350
rect 83918 256294 83986 256350
rect 84042 256294 114582 256350
rect 114638 256294 114706 256350
rect 114762 256294 145302 256350
rect 145358 256294 145426 256350
rect 145482 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 178518 256350
rect 178574 256294 178642 256350
rect 178698 256294 209238 256350
rect 209294 256294 209362 256350
rect 209418 256294 239958 256350
rect 240014 256294 240082 256350
rect 240138 256294 270678 256350
rect 270734 256294 270802 256350
rect 270858 256294 281994 256350
rect 282050 256294 282118 256350
rect 282174 256294 282242 256350
rect 282298 256294 282366 256350
rect 282422 256294 312714 256350
rect 312770 256294 312838 256350
rect 312894 256294 312962 256350
rect 313018 256294 313086 256350
rect 313142 256294 324518 256350
rect 324574 256294 324642 256350
rect 324698 256294 355238 256350
rect 355294 256294 355362 256350
rect 355418 256294 385958 256350
rect 386014 256294 386082 256350
rect 386138 256294 416678 256350
rect 416734 256294 416802 256350
rect 416858 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 448518 256350
rect 448574 256294 448642 256350
rect 448698 256294 479238 256350
rect 479294 256294 479362 256350
rect 479418 256294 509958 256350
rect 510014 256294 510082 256350
rect 510138 256294 540678 256350
rect 540734 256294 540802 256350
rect 540858 256294 571398 256350
rect 571454 256294 571522 256350
rect 571578 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 22422 256226
rect 22478 256170 22546 256226
rect 22602 256170 53142 256226
rect 53198 256170 53266 256226
rect 53322 256170 83862 256226
rect 83918 256170 83986 256226
rect 84042 256170 114582 256226
rect 114638 256170 114706 256226
rect 114762 256170 145302 256226
rect 145358 256170 145426 256226
rect 145482 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 178518 256226
rect 178574 256170 178642 256226
rect 178698 256170 209238 256226
rect 209294 256170 209362 256226
rect 209418 256170 239958 256226
rect 240014 256170 240082 256226
rect 240138 256170 270678 256226
rect 270734 256170 270802 256226
rect 270858 256170 281994 256226
rect 282050 256170 282118 256226
rect 282174 256170 282242 256226
rect 282298 256170 282366 256226
rect 282422 256170 312714 256226
rect 312770 256170 312838 256226
rect 312894 256170 312962 256226
rect 313018 256170 313086 256226
rect 313142 256170 324518 256226
rect 324574 256170 324642 256226
rect 324698 256170 355238 256226
rect 355294 256170 355362 256226
rect 355418 256170 385958 256226
rect 386014 256170 386082 256226
rect 386138 256170 416678 256226
rect 416734 256170 416802 256226
rect 416858 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 448518 256226
rect 448574 256170 448642 256226
rect 448698 256170 479238 256226
rect 479294 256170 479362 256226
rect 479418 256170 509958 256226
rect 510014 256170 510082 256226
rect 510138 256170 540678 256226
rect 540734 256170 540802 256226
rect 540858 256170 571398 256226
rect 571454 256170 571522 256226
rect 571578 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 22422 256102
rect 22478 256046 22546 256102
rect 22602 256046 53142 256102
rect 53198 256046 53266 256102
rect 53322 256046 83862 256102
rect 83918 256046 83986 256102
rect 84042 256046 114582 256102
rect 114638 256046 114706 256102
rect 114762 256046 145302 256102
rect 145358 256046 145426 256102
rect 145482 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 178518 256102
rect 178574 256046 178642 256102
rect 178698 256046 209238 256102
rect 209294 256046 209362 256102
rect 209418 256046 239958 256102
rect 240014 256046 240082 256102
rect 240138 256046 270678 256102
rect 270734 256046 270802 256102
rect 270858 256046 281994 256102
rect 282050 256046 282118 256102
rect 282174 256046 282242 256102
rect 282298 256046 282366 256102
rect 282422 256046 312714 256102
rect 312770 256046 312838 256102
rect 312894 256046 312962 256102
rect 313018 256046 313086 256102
rect 313142 256046 324518 256102
rect 324574 256046 324642 256102
rect 324698 256046 355238 256102
rect 355294 256046 355362 256102
rect 355418 256046 385958 256102
rect 386014 256046 386082 256102
rect 386138 256046 416678 256102
rect 416734 256046 416802 256102
rect 416858 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 448518 256102
rect 448574 256046 448642 256102
rect 448698 256046 479238 256102
rect 479294 256046 479362 256102
rect 479418 256046 509958 256102
rect 510014 256046 510082 256102
rect 510138 256046 540678 256102
rect 540734 256046 540802 256102
rect 540858 256046 571398 256102
rect 571454 256046 571522 256102
rect 571578 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 22422 255978
rect 22478 255922 22546 255978
rect 22602 255922 53142 255978
rect 53198 255922 53266 255978
rect 53322 255922 83862 255978
rect 83918 255922 83986 255978
rect 84042 255922 114582 255978
rect 114638 255922 114706 255978
rect 114762 255922 145302 255978
rect 145358 255922 145426 255978
rect 145482 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 178518 255978
rect 178574 255922 178642 255978
rect 178698 255922 209238 255978
rect 209294 255922 209362 255978
rect 209418 255922 239958 255978
rect 240014 255922 240082 255978
rect 240138 255922 270678 255978
rect 270734 255922 270802 255978
rect 270858 255922 281994 255978
rect 282050 255922 282118 255978
rect 282174 255922 282242 255978
rect 282298 255922 282366 255978
rect 282422 255922 312714 255978
rect 312770 255922 312838 255978
rect 312894 255922 312962 255978
rect 313018 255922 313086 255978
rect 313142 255922 324518 255978
rect 324574 255922 324642 255978
rect 324698 255922 355238 255978
rect 355294 255922 355362 255978
rect 355418 255922 385958 255978
rect 386014 255922 386082 255978
rect 386138 255922 416678 255978
rect 416734 255922 416802 255978
rect 416858 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 448518 255978
rect 448574 255922 448642 255978
rect 448698 255922 479238 255978
rect 479294 255922 479362 255978
rect 479418 255922 509958 255978
rect 510014 255922 510082 255978
rect 510138 255922 540678 255978
rect 540734 255922 540802 255978
rect 540858 255922 571398 255978
rect 571454 255922 571522 255978
rect 571578 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 37782 244350
rect 37838 244294 37906 244350
rect 37962 244294 68502 244350
rect 68558 244294 68626 244350
rect 68682 244294 99222 244350
rect 99278 244294 99346 244350
rect 99402 244294 129942 244350
rect 129998 244294 130066 244350
rect 130122 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193878 244350
rect 193934 244294 194002 244350
rect 194058 244294 224598 244350
rect 224654 244294 224722 244350
rect 224778 244294 255318 244350
rect 255374 244294 255442 244350
rect 255498 244294 285714 244350
rect 285770 244294 285838 244350
rect 285894 244294 285962 244350
rect 286018 244294 286086 244350
rect 286142 244294 316434 244350
rect 316490 244294 316558 244350
rect 316614 244294 316682 244350
rect 316738 244294 316806 244350
rect 316862 244294 339878 244350
rect 339934 244294 340002 244350
rect 340058 244294 370598 244350
rect 370654 244294 370722 244350
rect 370778 244294 401318 244350
rect 401374 244294 401442 244350
rect 401498 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 463878 244350
rect 463934 244294 464002 244350
rect 464058 244294 494598 244350
rect 494654 244294 494722 244350
rect 494778 244294 525318 244350
rect 525374 244294 525442 244350
rect 525498 244294 556038 244350
rect 556094 244294 556162 244350
rect 556218 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 37782 244226
rect 37838 244170 37906 244226
rect 37962 244170 68502 244226
rect 68558 244170 68626 244226
rect 68682 244170 99222 244226
rect 99278 244170 99346 244226
rect 99402 244170 129942 244226
rect 129998 244170 130066 244226
rect 130122 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193878 244226
rect 193934 244170 194002 244226
rect 194058 244170 224598 244226
rect 224654 244170 224722 244226
rect 224778 244170 255318 244226
rect 255374 244170 255442 244226
rect 255498 244170 285714 244226
rect 285770 244170 285838 244226
rect 285894 244170 285962 244226
rect 286018 244170 286086 244226
rect 286142 244170 316434 244226
rect 316490 244170 316558 244226
rect 316614 244170 316682 244226
rect 316738 244170 316806 244226
rect 316862 244170 339878 244226
rect 339934 244170 340002 244226
rect 340058 244170 370598 244226
rect 370654 244170 370722 244226
rect 370778 244170 401318 244226
rect 401374 244170 401442 244226
rect 401498 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 463878 244226
rect 463934 244170 464002 244226
rect 464058 244170 494598 244226
rect 494654 244170 494722 244226
rect 494778 244170 525318 244226
rect 525374 244170 525442 244226
rect 525498 244170 556038 244226
rect 556094 244170 556162 244226
rect 556218 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 37782 244102
rect 37838 244046 37906 244102
rect 37962 244046 68502 244102
rect 68558 244046 68626 244102
rect 68682 244046 99222 244102
rect 99278 244046 99346 244102
rect 99402 244046 129942 244102
rect 129998 244046 130066 244102
rect 130122 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193878 244102
rect 193934 244046 194002 244102
rect 194058 244046 224598 244102
rect 224654 244046 224722 244102
rect 224778 244046 255318 244102
rect 255374 244046 255442 244102
rect 255498 244046 285714 244102
rect 285770 244046 285838 244102
rect 285894 244046 285962 244102
rect 286018 244046 286086 244102
rect 286142 244046 316434 244102
rect 316490 244046 316558 244102
rect 316614 244046 316682 244102
rect 316738 244046 316806 244102
rect 316862 244046 339878 244102
rect 339934 244046 340002 244102
rect 340058 244046 370598 244102
rect 370654 244046 370722 244102
rect 370778 244046 401318 244102
rect 401374 244046 401442 244102
rect 401498 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 463878 244102
rect 463934 244046 464002 244102
rect 464058 244046 494598 244102
rect 494654 244046 494722 244102
rect 494778 244046 525318 244102
rect 525374 244046 525442 244102
rect 525498 244046 556038 244102
rect 556094 244046 556162 244102
rect 556218 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 37782 243978
rect 37838 243922 37906 243978
rect 37962 243922 68502 243978
rect 68558 243922 68626 243978
rect 68682 243922 99222 243978
rect 99278 243922 99346 243978
rect 99402 243922 129942 243978
rect 129998 243922 130066 243978
rect 130122 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193878 243978
rect 193934 243922 194002 243978
rect 194058 243922 224598 243978
rect 224654 243922 224722 243978
rect 224778 243922 255318 243978
rect 255374 243922 255442 243978
rect 255498 243922 285714 243978
rect 285770 243922 285838 243978
rect 285894 243922 285962 243978
rect 286018 243922 286086 243978
rect 286142 243922 316434 243978
rect 316490 243922 316558 243978
rect 316614 243922 316682 243978
rect 316738 243922 316806 243978
rect 316862 243922 339878 243978
rect 339934 243922 340002 243978
rect 340058 243922 370598 243978
rect 370654 243922 370722 243978
rect 370778 243922 401318 243978
rect 401374 243922 401442 243978
rect 401498 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 463878 243978
rect 463934 243922 464002 243978
rect 464058 243922 494598 243978
rect 494654 243922 494722 243978
rect 494778 243922 525318 243978
rect 525374 243922 525442 243978
rect 525498 243922 556038 243978
rect 556094 243922 556162 243978
rect 556218 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 22422 238350
rect 22478 238294 22546 238350
rect 22602 238294 53142 238350
rect 53198 238294 53266 238350
rect 53322 238294 83862 238350
rect 83918 238294 83986 238350
rect 84042 238294 114582 238350
rect 114638 238294 114706 238350
rect 114762 238294 145302 238350
rect 145358 238294 145426 238350
rect 145482 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 178518 238350
rect 178574 238294 178642 238350
rect 178698 238294 209238 238350
rect 209294 238294 209362 238350
rect 209418 238294 239958 238350
rect 240014 238294 240082 238350
rect 240138 238294 270678 238350
rect 270734 238294 270802 238350
rect 270858 238294 281994 238350
rect 282050 238294 282118 238350
rect 282174 238294 282242 238350
rect 282298 238294 282366 238350
rect 282422 238294 312714 238350
rect 312770 238294 312838 238350
rect 312894 238294 312962 238350
rect 313018 238294 313086 238350
rect 313142 238294 324518 238350
rect 324574 238294 324642 238350
rect 324698 238294 355238 238350
rect 355294 238294 355362 238350
rect 355418 238294 385958 238350
rect 386014 238294 386082 238350
rect 386138 238294 416678 238350
rect 416734 238294 416802 238350
rect 416858 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 448518 238350
rect 448574 238294 448642 238350
rect 448698 238294 479238 238350
rect 479294 238294 479362 238350
rect 479418 238294 509958 238350
rect 510014 238294 510082 238350
rect 510138 238294 540678 238350
rect 540734 238294 540802 238350
rect 540858 238294 571398 238350
rect 571454 238294 571522 238350
rect 571578 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 22422 238226
rect 22478 238170 22546 238226
rect 22602 238170 53142 238226
rect 53198 238170 53266 238226
rect 53322 238170 83862 238226
rect 83918 238170 83986 238226
rect 84042 238170 114582 238226
rect 114638 238170 114706 238226
rect 114762 238170 145302 238226
rect 145358 238170 145426 238226
rect 145482 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 178518 238226
rect 178574 238170 178642 238226
rect 178698 238170 209238 238226
rect 209294 238170 209362 238226
rect 209418 238170 239958 238226
rect 240014 238170 240082 238226
rect 240138 238170 270678 238226
rect 270734 238170 270802 238226
rect 270858 238170 281994 238226
rect 282050 238170 282118 238226
rect 282174 238170 282242 238226
rect 282298 238170 282366 238226
rect 282422 238170 312714 238226
rect 312770 238170 312838 238226
rect 312894 238170 312962 238226
rect 313018 238170 313086 238226
rect 313142 238170 324518 238226
rect 324574 238170 324642 238226
rect 324698 238170 355238 238226
rect 355294 238170 355362 238226
rect 355418 238170 385958 238226
rect 386014 238170 386082 238226
rect 386138 238170 416678 238226
rect 416734 238170 416802 238226
rect 416858 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 448518 238226
rect 448574 238170 448642 238226
rect 448698 238170 479238 238226
rect 479294 238170 479362 238226
rect 479418 238170 509958 238226
rect 510014 238170 510082 238226
rect 510138 238170 540678 238226
rect 540734 238170 540802 238226
rect 540858 238170 571398 238226
rect 571454 238170 571522 238226
rect 571578 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 22422 238102
rect 22478 238046 22546 238102
rect 22602 238046 53142 238102
rect 53198 238046 53266 238102
rect 53322 238046 83862 238102
rect 83918 238046 83986 238102
rect 84042 238046 114582 238102
rect 114638 238046 114706 238102
rect 114762 238046 145302 238102
rect 145358 238046 145426 238102
rect 145482 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 178518 238102
rect 178574 238046 178642 238102
rect 178698 238046 209238 238102
rect 209294 238046 209362 238102
rect 209418 238046 239958 238102
rect 240014 238046 240082 238102
rect 240138 238046 270678 238102
rect 270734 238046 270802 238102
rect 270858 238046 281994 238102
rect 282050 238046 282118 238102
rect 282174 238046 282242 238102
rect 282298 238046 282366 238102
rect 282422 238046 312714 238102
rect 312770 238046 312838 238102
rect 312894 238046 312962 238102
rect 313018 238046 313086 238102
rect 313142 238046 324518 238102
rect 324574 238046 324642 238102
rect 324698 238046 355238 238102
rect 355294 238046 355362 238102
rect 355418 238046 385958 238102
rect 386014 238046 386082 238102
rect 386138 238046 416678 238102
rect 416734 238046 416802 238102
rect 416858 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 448518 238102
rect 448574 238046 448642 238102
rect 448698 238046 479238 238102
rect 479294 238046 479362 238102
rect 479418 238046 509958 238102
rect 510014 238046 510082 238102
rect 510138 238046 540678 238102
rect 540734 238046 540802 238102
rect 540858 238046 571398 238102
rect 571454 238046 571522 238102
rect 571578 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 22422 237978
rect 22478 237922 22546 237978
rect 22602 237922 53142 237978
rect 53198 237922 53266 237978
rect 53322 237922 83862 237978
rect 83918 237922 83986 237978
rect 84042 237922 114582 237978
rect 114638 237922 114706 237978
rect 114762 237922 145302 237978
rect 145358 237922 145426 237978
rect 145482 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 178518 237978
rect 178574 237922 178642 237978
rect 178698 237922 209238 237978
rect 209294 237922 209362 237978
rect 209418 237922 239958 237978
rect 240014 237922 240082 237978
rect 240138 237922 270678 237978
rect 270734 237922 270802 237978
rect 270858 237922 281994 237978
rect 282050 237922 282118 237978
rect 282174 237922 282242 237978
rect 282298 237922 282366 237978
rect 282422 237922 312714 237978
rect 312770 237922 312838 237978
rect 312894 237922 312962 237978
rect 313018 237922 313086 237978
rect 313142 237922 324518 237978
rect 324574 237922 324642 237978
rect 324698 237922 355238 237978
rect 355294 237922 355362 237978
rect 355418 237922 385958 237978
rect 386014 237922 386082 237978
rect 386138 237922 416678 237978
rect 416734 237922 416802 237978
rect 416858 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 448518 237978
rect 448574 237922 448642 237978
rect 448698 237922 479238 237978
rect 479294 237922 479362 237978
rect 479418 237922 509958 237978
rect 510014 237922 510082 237978
rect 510138 237922 540678 237978
rect 540734 237922 540802 237978
rect 540858 237922 571398 237978
rect 571454 237922 571522 237978
rect 571578 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 37782 226350
rect 37838 226294 37906 226350
rect 37962 226294 68502 226350
rect 68558 226294 68626 226350
rect 68682 226294 99222 226350
rect 99278 226294 99346 226350
rect 99402 226294 129942 226350
rect 129998 226294 130066 226350
rect 130122 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193878 226350
rect 193934 226294 194002 226350
rect 194058 226294 224598 226350
rect 224654 226294 224722 226350
rect 224778 226294 255318 226350
rect 255374 226294 255442 226350
rect 255498 226294 285714 226350
rect 285770 226294 285838 226350
rect 285894 226294 285962 226350
rect 286018 226294 286086 226350
rect 286142 226294 316434 226350
rect 316490 226294 316558 226350
rect 316614 226294 316682 226350
rect 316738 226294 316806 226350
rect 316862 226294 339878 226350
rect 339934 226294 340002 226350
rect 340058 226294 370598 226350
rect 370654 226294 370722 226350
rect 370778 226294 401318 226350
rect 401374 226294 401442 226350
rect 401498 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 463878 226350
rect 463934 226294 464002 226350
rect 464058 226294 494598 226350
rect 494654 226294 494722 226350
rect 494778 226294 525318 226350
rect 525374 226294 525442 226350
rect 525498 226294 556038 226350
rect 556094 226294 556162 226350
rect 556218 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 37782 226226
rect 37838 226170 37906 226226
rect 37962 226170 68502 226226
rect 68558 226170 68626 226226
rect 68682 226170 99222 226226
rect 99278 226170 99346 226226
rect 99402 226170 129942 226226
rect 129998 226170 130066 226226
rect 130122 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193878 226226
rect 193934 226170 194002 226226
rect 194058 226170 224598 226226
rect 224654 226170 224722 226226
rect 224778 226170 255318 226226
rect 255374 226170 255442 226226
rect 255498 226170 285714 226226
rect 285770 226170 285838 226226
rect 285894 226170 285962 226226
rect 286018 226170 286086 226226
rect 286142 226170 316434 226226
rect 316490 226170 316558 226226
rect 316614 226170 316682 226226
rect 316738 226170 316806 226226
rect 316862 226170 339878 226226
rect 339934 226170 340002 226226
rect 340058 226170 370598 226226
rect 370654 226170 370722 226226
rect 370778 226170 401318 226226
rect 401374 226170 401442 226226
rect 401498 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 463878 226226
rect 463934 226170 464002 226226
rect 464058 226170 494598 226226
rect 494654 226170 494722 226226
rect 494778 226170 525318 226226
rect 525374 226170 525442 226226
rect 525498 226170 556038 226226
rect 556094 226170 556162 226226
rect 556218 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 37782 226102
rect 37838 226046 37906 226102
rect 37962 226046 68502 226102
rect 68558 226046 68626 226102
rect 68682 226046 99222 226102
rect 99278 226046 99346 226102
rect 99402 226046 129942 226102
rect 129998 226046 130066 226102
rect 130122 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193878 226102
rect 193934 226046 194002 226102
rect 194058 226046 224598 226102
rect 224654 226046 224722 226102
rect 224778 226046 255318 226102
rect 255374 226046 255442 226102
rect 255498 226046 285714 226102
rect 285770 226046 285838 226102
rect 285894 226046 285962 226102
rect 286018 226046 286086 226102
rect 286142 226046 316434 226102
rect 316490 226046 316558 226102
rect 316614 226046 316682 226102
rect 316738 226046 316806 226102
rect 316862 226046 339878 226102
rect 339934 226046 340002 226102
rect 340058 226046 370598 226102
rect 370654 226046 370722 226102
rect 370778 226046 401318 226102
rect 401374 226046 401442 226102
rect 401498 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 463878 226102
rect 463934 226046 464002 226102
rect 464058 226046 494598 226102
rect 494654 226046 494722 226102
rect 494778 226046 525318 226102
rect 525374 226046 525442 226102
rect 525498 226046 556038 226102
rect 556094 226046 556162 226102
rect 556218 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 37782 225978
rect 37838 225922 37906 225978
rect 37962 225922 68502 225978
rect 68558 225922 68626 225978
rect 68682 225922 99222 225978
rect 99278 225922 99346 225978
rect 99402 225922 129942 225978
rect 129998 225922 130066 225978
rect 130122 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193878 225978
rect 193934 225922 194002 225978
rect 194058 225922 224598 225978
rect 224654 225922 224722 225978
rect 224778 225922 255318 225978
rect 255374 225922 255442 225978
rect 255498 225922 285714 225978
rect 285770 225922 285838 225978
rect 285894 225922 285962 225978
rect 286018 225922 286086 225978
rect 286142 225922 316434 225978
rect 316490 225922 316558 225978
rect 316614 225922 316682 225978
rect 316738 225922 316806 225978
rect 316862 225922 339878 225978
rect 339934 225922 340002 225978
rect 340058 225922 370598 225978
rect 370654 225922 370722 225978
rect 370778 225922 401318 225978
rect 401374 225922 401442 225978
rect 401498 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 463878 225978
rect 463934 225922 464002 225978
rect 464058 225922 494598 225978
rect 494654 225922 494722 225978
rect 494778 225922 525318 225978
rect 525374 225922 525442 225978
rect 525498 225922 556038 225978
rect 556094 225922 556162 225978
rect 556218 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 22422 220350
rect 22478 220294 22546 220350
rect 22602 220294 53142 220350
rect 53198 220294 53266 220350
rect 53322 220294 83862 220350
rect 83918 220294 83986 220350
rect 84042 220294 114582 220350
rect 114638 220294 114706 220350
rect 114762 220294 145302 220350
rect 145358 220294 145426 220350
rect 145482 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 178518 220350
rect 178574 220294 178642 220350
rect 178698 220294 209238 220350
rect 209294 220294 209362 220350
rect 209418 220294 239958 220350
rect 240014 220294 240082 220350
rect 240138 220294 270678 220350
rect 270734 220294 270802 220350
rect 270858 220294 281994 220350
rect 282050 220294 282118 220350
rect 282174 220294 282242 220350
rect 282298 220294 282366 220350
rect 282422 220294 312714 220350
rect 312770 220294 312838 220350
rect 312894 220294 312962 220350
rect 313018 220294 313086 220350
rect 313142 220294 324518 220350
rect 324574 220294 324642 220350
rect 324698 220294 355238 220350
rect 355294 220294 355362 220350
rect 355418 220294 385958 220350
rect 386014 220294 386082 220350
rect 386138 220294 416678 220350
rect 416734 220294 416802 220350
rect 416858 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 448518 220350
rect 448574 220294 448642 220350
rect 448698 220294 479238 220350
rect 479294 220294 479362 220350
rect 479418 220294 509958 220350
rect 510014 220294 510082 220350
rect 510138 220294 540678 220350
rect 540734 220294 540802 220350
rect 540858 220294 571398 220350
rect 571454 220294 571522 220350
rect 571578 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 22422 220226
rect 22478 220170 22546 220226
rect 22602 220170 53142 220226
rect 53198 220170 53266 220226
rect 53322 220170 83862 220226
rect 83918 220170 83986 220226
rect 84042 220170 114582 220226
rect 114638 220170 114706 220226
rect 114762 220170 145302 220226
rect 145358 220170 145426 220226
rect 145482 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 178518 220226
rect 178574 220170 178642 220226
rect 178698 220170 209238 220226
rect 209294 220170 209362 220226
rect 209418 220170 239958 220226
rect 240014 220170 240082 220226
rect 240138 220170 270678 220226
rect 270734 220170 270802 220226
rect 270858 220170 281994 220226
rect 282050 220170 282118 220226
rect 282174 220170 282242 220226
rect 282298 220170 282366 220226
rect 282422 220170 312714 220226
rect 312770 220170 312838 220226
rect 312894 220170 312962 220226
rect 313018 220170 313086 220226
rect 313142 220170 324518 220226
rect 324574 220170 324642 220226
rect 324698 220170 355238 220226
rect 355294 220170 355362 220226
rect 355418 220170 385958 220226
rect 386014 220170 386082 220226
rect 386138 220170 416678 220226
rect 416734 220170 416802 220226
rect 416858 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 448518 220226
rect 448574 220170 448642 220226
rect 448698 220170 479238 220226
rect 479294 220170 479362 220226
rect 479418 220170 509958 220226
rect 510014 220170 510082 220226
rect 510138 220170 540678 220226
rect 540734 220170 540802 220226
rect 540858 220170 571398 220226
rect 571454 220170 571522 220226
rect 571578 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 22422 220102
rect 22478 220046 22546 220102
rect 22602 220046 53142 220102
rect 53198 220046 53266 220102
rect 53322 220046 83862 220102
rect 83918 220046 83986 220102
rect 84042 220046 114582 220102
rect 114638 220046 114706 220102
rect 114762 220046 145302 220102
rect 145358 220046 145426 220102
rect 145482 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 178518 220102
rect 178574 220046 178642 220102
rect 178698 220046 209238 220102
rect 209294 220046 209362 220102
rect 209418 220046 239958 220102
rect 240014 220046 240082 220102
rect 240138 220046 270678 220102
rect 270734 220046 270802 220102
rect 270858 220046 281994 220102
rect 282050 220046 282118 220102
rect 282174 220046 282242 220102
rect 282298 220046 282366 220102
rect 282422 220046 312714 220102
rect 312770 220046 312838 220102
rect 312894 220046 312962 220102
rect 313018 220046 313086 220102
rect 313142 220046 324518 220102
rect 324574 220046 324642 220102
rect 324698 220046 355238 220102
rect 355294 220046 355362 220102
rect 355418 220046 385958 220102
rect 386014 220046 386082 220102
rect 386138 220046 416678 220102
rect 416734 220046 416802 220102
rect 416858 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 448518 220102
rect 448574 220046 448642 220102
rect 448698 220046 479238 220102
rect 479294 220046 479362 220102
rect 479418 220046 509958 220102
rect 510014 220046 510082 220102
rect 510138 220046 540678 220102
rect 540734 220046 540802 220102
rect 540858 220046 571398 220102
rect 571454 220046 571522 220102
rect 571578 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 22422 219978
rect 22478 219922 22546 219978
rect 22602 219922 53142 219978
rect 53198 219922 53266 219978
rect 53322 219922 83862 219978
rect 83918 219922 83986 219978
rect 84042 219922 114582 219978
rect 114638 219922 114706 219978
rect 114762 219922 145302 219978
rect 145358 219922 145426 219978
rect 145482 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 178518 219978
rect 178574 219922 178642 219978
rect 178698 219922 209238 219978
rect 209294 219922 209362 219978
rect 209418 219922 239958 219978
rect 240014 219922 240082 219978
rect 240138 219922 270678 219978
rect 270734 219922 270802 219978
rect 270858 219922 281994 219978
rect 282050 219922 282118 219978
rect 282174 219922 282242 219978
rect 282298 219922 282366 219978
rect 282422 219922 312714 219978
rect 312770 219922 312838 219978
rect 312894 219922 312962 219978
rect 313018 219922 313086 219978
rect 313142 219922 324518 219978
rect 324574 219922 324642 219978
rect 324698 219922 355238 219978
rect 355294 219922 355362 219978
rect 355418 219922 385958 219978
rect 386014 219922 386082 219978
rect 386138 219922 416678 219978
rect 416734 219922 416802 219978
rect 416858 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 448518 219978
rect 448574 219922 448642 219978
rect 448698 219922 479238 219978
rect 479294 219922 479362 219978
rect 479418 219922 509958 219978
rect 510014 219922 510082 219978
rect 510138 219922 540678 219978
rect 540734 219922 540802 219978
rect 540858 219922 571398 219978
rect 571454 219922 571522 219978
rect 571578 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 37782 208350
rect 37838 208294 37906 208350
rect 37962 208294 68502 208350
rect 68558 208294 68626 208350
rect 68682 208294 99222 208350
rect 99278 208294 99346 208350
rect 99402 208294 129942 208350
rect 129998 208294 130066 208350
rect 130122 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 193878 208350
rect 193934 208294 194002 208350
rect 194058 208294 224598 208350
rect 224654 208294 224722 208350
rect 224778 208294 255318 208350
rect 255374 208294 255442 208350
rect 255498 208294 285714 208350
rect 285770 208294 285838 208350
rect 285894 208294 285962 208350
rect 286018 208294 286086 208350
rect 286142 208294 316434 208350
rect 316490 208294 316558 208350
rect 316614 208294 316682 208350
rect 316738 208294 316806 208350
rect 316862 208294 339878 208350
rect 339934 208294 340002 208350
rect 340058 208294 370598 208350
rect 370654 208294 370722 208350
rect 370778 208294 401318 208350
rect 401374 208294 401442 208350
rect 401498 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 463878 208350
rect 463934 208294 464002 208350
rect 464058 208294 494598 208350
rect 494654 208294 494722 208350
rect 494778 208294 525318 208350
rect 525374 208294 525442 208350
rect 525498 208294 556038 208350
rect 556094 208294 556162 208350
rect 556218 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 37782 208226
rect 37838 208170 37906 208226
rect 37962 208170 68502 208226
rect 68558 208170 68626 208226
rect 68682 208170 99222 208226
rect 99278 208170 99346 208226
rect 99402 208170 129942 208226
rect 129998 208170 130066 208226
rect 130122 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 193878 208226
rect 193934 208170 194002 208226
rect 194058 208170 224598 208226
rect 224654 208170 224722 208226
rect 224778 208170 255318 208226
rect 255374 208170 255442 208226
rect 255498 208170 285714 208226
rect 285770 208170 285838 208226
rect 285894 208170 285962 208226
rect 286018 208170 286086 208226
rect 286142 208170 316434 208226
rect 316490 208170 316558 208226
rect 316614 208170 316682 208226
rect 316738 208170 316806 208226
rect 316862 208170 339878 208226
rect 339934 208170 340002 208226
rect 340058 208170 370598 208226
rect 370654 208170 370722 208226
rect 370778 208170 401318 208226
rect 401374 208170 401442 208226
rect 401498 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 463878 208226
rect 463934 208170 464002 208226
rect 464058 208170 494598 208226
rect 494654 208170 494722 208226
rect 494778 208170 525318 208226
rect 525374 208170 525442 208226
rect 525498 208170 556038 208226
rect 556094 208170 556162 208226
rect 556218 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 37782 208102
rect 37838 208046 37906 208102
rect 37962 208046 68502 208102
rect 68558 208046 68626 208102
rect 68682 208046 99222 208102
rect 99278 208046 99346 208102
rect 99402 208046 129942 208102
rect 129998 208046 130066 208102
rect 130122 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 193878 208102
rect 193934 208046 194002 208102
rect 194058 208046 224598 208102
rect 224654 208046 224722 208102
rect 224778 208046 255318 208102
rect 255374 208046 255442 208102
rect 255498 208046 285714 208102
rect 285770 208046 285838 208102
rect 285894 208046 285962 208102
rect 286018 208046 286086 208102
rect 286142 208046 316434 208102
rect 316490 208046 316558 208102
rect 316614 208046 316682 208102
rect 316738 208046 316806 208102
rect 316862 208046 339878 208102
rect 339934 208046 340002 208102
rect 340058 208046 370598 208102
rect 370654 208046 370722 208102
rect 370778 208046 401318 208102
rect 401374 208046 401442 208102
rect 401498 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 463878 208102
rect 463934 208046 464002 208102
rect 464058 208046 494598 208102
rect 494654 208046 494722 208102
rect 494778 208046 525318 208102
rect 525374 208046 525442 208102
rect 525498 208046 556038 208102
rect 556094 208046 556162 208102
rect 556218 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 37782 207978
rect 37838 207922 37906 207978
rect 37962 207922 68502 207978
rect 68558 207922 68626 207978
rect 68682 207922 99222 207978
rect 99278 207922 99346 207978
rect 99402 207922 129942 207978
rect 129998 207922 130066 207978
rect 130122 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 193878 207978
rect 193934 207922 194002 207978
rect 194058 207922 224598 207978
rect 224654 207922 224722 207978
rect 224778 207922 255318 207978
rect 255374 207922 255442 207978
rect 255498 207922 285714 207978
rect 285770 207922 285838 207978
rect 285894 207922 285962 207978
rect 286018 207922 286086 207978
rect 286142 207922 316434 207978
rect 316490 207922 316558 207978
rect 316614 207922 316682 207978
rect 316738 207922 316806 207978
rect 316862 207922 339878 207978
rect 339934 207922 340002 207978
rect 340058 207922 370598 207978
rect 370654 207922 370722 207978
rect 370778 207922 401318 207978
rect 401374 207922 401442 207978
rect 401498 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 463878 207978
rect 463934 207922 464002 207978
rect 464058 207922 494598 207978
rect 494654 207922 494722 207978
rect 494778 207922 525318 207978
rect 525374 207922 525442 207978
rect 525498 207922 556038 207978
rect 556094 207922 556162 207978
rect 556218 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 22422 202350
rect 22478 202294 22546 202350
rect 22602 202294 53142 202350
rect 53198 202294 53266 202350
rect 53322 202294 83862 202350
rect 83918 202294 83986 202350
rect 84042 202294 114582 202350
rect 114638 202294 114706 202350
rect 114762 202294 145302 202350
rect 145358 202294 145426 202350
rect 145482 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 178518 202350
rect 178574 202294 178642 202350
rect 178698 202294 209238 202350
rect 209294 202294 209362 202350
rect 209418 202294 239958 202350
rect 240014 202294 240082 202350
rect 240138 202294 270678 202350
rect 270734 202294 270802 202350
rect 270858 202294 281994 202350
rect 282050 202294 282118 202350
rect 282174 202294 282242 202350
rect 282298 202294 282366 202350
rect 282422 202294 312714 202350
rect 312770 202294 312838 202350
rect 312894 202294 312962 202350
rect 313018 202294 313086 202350
rect 313142 202294 324518 202350
rect 324574 202294 324642 202350
rect 324698 202294 355238 202350
rect 355294 202294 355362 202350
rect 355418 202294 385958 202350
rect 386014 202294 386082 202350
rect 386138 202294 416678 202350
rect 416734 202294 416802 202350
rect 416858 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 448518 202350
rect 448574 202294 448642 202350
rect 448698 202294 479238 202350
rect 479294 202294 479362 202350
rect 479418 202294 509958 202350
rect 510014 202294 510082 202350
rect 510138 202294 540678 202350
rect 540734 202294 540802 202350
rect 540858 202294 571398 202350
rect 571454 202294 571522 202350
rect 571578 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 22422 202226
rect 22478 202170 22546 202226
rect 22602 202170 53142 202226
rect 53198 202170 53266 202226
rect 53322 202170 83862 202226
rect 83918 202170 83986 202226
rect 84042 202170 114582 202226
rect 114638 202170 114706 202226
rect 114762 202170 145302 202226
rect 145358 202170 145426 202226
rect 145482 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 178518 202226
rect 178574 202170 178642 202226
rect 178698 202170 209238 202226
rect 209294 202170 209362 202226
rect 209418 202170 239958 202226
rect 240014 202170 240082 202226
rect 240138 202170 270678 202226
rect 270734 202170 270802 202226
rect 270858 202170 281994 202226
rect 282050 202170 282118 202226
rect 282174 202170 282242 202226
rect 282298 202170 282366 202226
rect 282422 202170 312714 202226
rect 312770 202170 312838 202226
rect 312894 202170 312962 202226
rect 313018 202170 313086 202226
rect 313142 202170 324518 202226
rect 324574 202170 324642 202226
rect 324698 202170 355238 202226
rect 355294 202170 355362 202226
rect 355418 202170 385958 202226
rect 386014 202170 386082 202226
rect 386138 202170 416678 202226
rect 416734 202170 416802 202226
rect 416858 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 448518 202226
rect 448574 202170 448642 202226
rect 448698 202170 479238 202226
rect 479294 202170 479362 202226
rect 479418 202170 509958 202226
rect 510014 202170 510082 202226
rect 510138 202170 540678 202226
rect 540734 202170 540802 202226
rect 540858 202170 571398 202226
rect 571454 202170 571522 202226
rect 571578 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 22422 202102
rect 22478 202046 22546 202102
rect 22602 202046 53142 202102
rect 53198 202046 53266 202102
rect 53322 202046 83862 202102
rect 83918 202046 83986 202102
rect 84042 202046 114582 202102
rect 114638 202046 114706 202102
rect 114762 202046 145302 202102
rect 145358 202046 145426 202102
rect 145482 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 178518 202102
rect 178574 202046 178642 202102
rect 178698 202046 209238 202102
rect 209294 202046 209362 202102
rect 209418 202046 239958 202102
rect 240014 202046 240082 202102
rect 240138 202046 270678 202102
rect 270734 202046 270802 202102
rect 270858 202046 281994 202102
rect 282050 202046 282118 202102
rect 282174 202046 282242 202102
rect 282298 202046 282366 202102
rect 282422 202046 312714 202102
rect 312770 202046 312838 202102
rect 312894 202046 312962 202102
rect 313018 202046 313086 202102
rect 313142 202046 324518 202102
rect 324574 202046 324642 202102
rect 324698 202046 355238 202102
rect 355294 202046 355362 202102
rect 355418 202046 385958 202102
rect 386014 202046 386082 202102
rect 386138 202046 416678 202102
rect 416734 202046 416802 202102
rect 416858 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 448518 202102
rect 448574 202046 448642 202102
rect 448698 202046 479238 202102
rect 479294 202046 479362 202102
rect 479418 202046 509958 202102
rect 510014 202046 510082 202102
rect 510138 202046 540678 202102
rect 540734 202046 540802 202102
rect 540858 202046 571398 202102
rect 571454 202046 571522 202102
rect 571578 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 22422 201978
rect 22478 201922 22546 201978
rect 22602 201922 53142 201978
rect 53198 201922 53266 201978
rect 53322 201922 83862 201978
rect 83918 201922 83986 201978
rect 84042 201922 114582 201978
rect 114638 201922 114706 201978
rect 114762 201922 145302 201978
rect 145358 201922 145426 201978
rect 145482 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 178518 201978
rect 178574 201922 178642 201978
rect 178698 201922 209238 201978
rect 209294 201922 209362 201978
rect 209418 201922 239958 201978
rect 240014 201922 240082 201978
rect 240138 201922 270678 201978
rect 270734 201922 270802 201978
rect 270858 201922 281994 201978
rect 282050 201922 282118 201978
rect 282174 201922 282242 201978
rect 282298 201922 282366 201978
rect 282422 201922 312714 201978
rect 312770 201922 312838 201978
rect 312894 201922 312962 201978
rect 313018 201922 313086 201978
rect 313142 201922 324518 201978
rect 324574 201922 324642 201978
rect 324698 201922 355238 201978
rect 355294 201922 355362 201978
rect 355418 201922 385958 201978
rect 386014 201922 386082 201978
rect 386138 201922 416678 201978
rect 416734 201922 416802 201978
rect 416858 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 448518 201978
rect 448574 201922 448642 201978
rect 448698 201922 479238 201978
rect 479294 201922 479362 201978
rect 479418 201922 509958 201978
rect 510014 201922 510082 201978
rect 510138 201922 540678 201978
rect 540734 201922 540802 201978
rect 540858 201922 571398 201978
rect 571454 201922 571522 201978
rect 571578 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 37782 190350
rect 37838 190294 37906 190350
rect 37962 190294 68502 190350
rect 68558 190294 68626 190350
rect 68682 190294 99222 190350
rect 99278 190294 99346 190350
rect 99402 190294 129942 190350
rect 129998 190294 130066 190350
rect 130122 190294 162834 190350
rect 162890 190294 162958 190350
rect 163014 190294 163082 190350
rect 163138 190294 163206 190350
rect 163262 190294 193878 190350
rect 193934 190294 194002 190350
rect 194058 190294 224598 190350
rect 224654 190294 224722 190350
rect 224778 190294 255318 190350
rect 255374 190294 255442 190350
rect 255498 190294 285714 190350
rect 285770 190294 285838 190350
rect 285894 190294 285962 190350
rect 286018 190294 286086 190350
rect 286142 190294 316434 190350
rect 316490 190294 316558 190350
rect 316614 190294 316682 190350
rect 316738 190294 316806 190350
rect 316862 190294 339878 190350
rect 339934 190294 340002 190350
rect 340058 190294 370598 190350
rect 370654 190294 370722 190350
rect 370778 190294 401318 190350
rect 401374 190294 401442 190350
rect 401498 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 463878 190350
rect 463934 190294 464002 190350
rect 464058 190294 494598 190350
rect 494654 190294 494722 190350
rect 494778 190294 525318 190350
rect 525374 190294 525442 190350
rect 525498 190294 556038 190350
rect 556094 190294 556162 190350
rect 556218 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 37782 190226
rect 37838 190170 37906 190226
rect 37962 190170 68502 190226
rect 68558 190170 68626 190226
rect 68682 190170 99222 190226
rect 99278 190170 99346 190226
rect 99402 190170 129942 190226
rect 129998 190170 130066 190226
rect 130122 190170 162834 190226
rect 162890 190170 162958 190226
rect 163014 190170 163082 190226
rect 163138 190170 163206 190226
rect 163262 190170 193878 190226
rect 193934 190170 194002 190226
rect 194058 190170 224598 190226
rect 224654 190170 224722 190226
rect 224778 190170 255318 190226
rect 255374 190170 255442 190226
rect 255498 190170 285714 190226
rect 285770 190170 285838 190226
rect 285894 190170 285962 190226
rect 286018 190170 286086 190226
rect 286142 190170 316434 190226
rect 316490 190170 316558 190226
rect 316614 190170 316682 190226
rect 316738 190170 316806 190226
rect 316862 190170 339878 190226
rect 339934 190170 340002 190226
rect 340058 190170 370598 190226
rect 370654 190170 370722 190226
rect 370778 190170 401318 190226
rect 401374 190170 401442 190226
rect 401498 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 463878 190226
rect 463934 190170 464002 190226
rect 464058 190170 494598 190226
rect 494654 190170 494722 190226
rect 494778 190170 525318 190226
rect 525374 190170 525442 190226
rect 525498 190170 556038 190226
rect 556094 190170 556162 190226
rect 556218 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 37782 190102
rect 37838 190046 37906 190102
rect 37962 190046 68502 190102
rect 68558 190046 68626 190102
rect 68682 190046 99222 190102
rect 99278 190046 99346 190102
rect 99402 190046 129942 190102
rect 129998 190046 130066 190102
rect 130122 190046 162834 190102
rect 162890 190046 162958 190102
rect 163014 190046 163082 190102
rect 163138 190046 163206 190102
rect 163262 190046 193878 190102
rect 193934 190046 194002 190102
rect 194058 190046 224598 190102
rect 224654 190046 224722 190102
rect 224778 190046 255318 190102
rect 255374 190046 255442 190102
rect 255498 190046 285714 190102
rect 285770 190046 285838 190102
rect 285894 190046 285962 190102
rect 286018 190046 286086 190102
rect 286142 190046 316434 190102
rect 316490 190046 316558 190102
rect 316614 190046 316682 190102
rect 316738 190046 316806 190102
rect 316862 190046 339878 190102
rect 339934 190046 340002 190102
rect 340058 190046 370598 190102
rect 370654 190046 370722 190102
rect 370778 190046 401318 190102
rect 401374 190046 401442 190102
rect 401498 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 463878 190102
rect 463934 190046 464002 190102
rect 464058 190046 494598 190102
rect 494654 190046 494722 190102
rect 494778 190046 525318 190102
rect 525374 190046 525442 190102
rect 525498 190046 556038 190102
rect 556094 190046 556162 190102
rect 556218 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 37782 189978
rect 37838 189922 37906 189978
rect 37962 189922 68502 189978
rect 68558 189922 68626 189978
rect 68682 189922 99222 189978
rect 99278 189922 99346 189978
rect 99402 189922 129942 189978
rect 129998 189922 130066 189978
rect 130122 189922 162834 189978
rect 162890 189922 162958 189978
rect 163014 189922 163082 189978
rect 163138 189922 163206 189978
rect 163262 189922 193878 189978
rect 193934 189922 194002 189978
rect 194058 189922 224598 189978
rect 224654 189922 224722 189978
rect 224778 189922 255318 189978
rect 255374 189922 255442 189978
rect 255498 189922 285714 189978
rect 285770 189922 285838 189978
rect 285894 189922 285962 189978
rect 286018 189922 286086 189978
rect 286142 189922 316434 189978
rect 316490 189922 316558 189978
rect 316614 189922 316682 189978
rect 316738 189922 316806 189978
rect 316862 189922 339878 189978
rect 339934 189922 340002 189978
rect 340058 189922 370598 189978
rect 370654 189922 370722 189978
rect 370778 189922 401318 189978
rect 401374 189922 401442 189978
rect 401498 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 463878 189978
rect 463934 189922 464002 189978
rect 464058 189922 494598 189978
rect 494654 189922 494722 189978
rect 494778 189922 525318 189978
rect 525374 189922 525442 189978
rect 525498 189922 556038 189978
rect 556094 189922 556162 189978
rect 556218 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 22422 184350
rect 22478 184294 22546 184350
rect 22602 184294 53142 184350
rect 53198 184294 53266 184350
rect 53322 184294 83862 184350
rect 83918 184294 83986 184350
rect 84042 184294 114582 184350
rect 114638 184294 114706 184350
rect 114762 184294 145302 184350
rect 145358 184294 145426 184350
rect 145482 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 178518 184350
rect 178574 184294 178642 184350
rect 178698 184294 209238 184350
rect 209294 184294 209362 184350
rect 209418 184294 239958 184350
rect 240014 184294 240082 184350
rect 240138 184294 270678 184350
rect 270734 184294 270802 184350
rect 270858 184294 281994 184350
rect 282050 184294 282118 184350
rect 282174 184294 282242 184350
rect 282298 184294 282366 184350
rect 282422 184294 312714 184350
rect 312770 184294 312838 184350
rect 312894 184294 312962 184350
rect 313018 184294 313086 184350
rect 313142 184294 324518 184350
rect 324574 184294 324642 184350
rect 324698 184294 355238 184350
rect 355294 184294 355362 184350
rect 355418 184294 385958 184350
rect 386014 184294 386082 184350
rect 386138 184294 416678 184350
rect 416734 184294 416802 184350
rect 416858 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 448518 184350
rect 448574 184294 448642 184350
rect 448698 184294 479238 184350
rect 479294 184294 479362 184350
rect 479418 184294 509958 184350
rect 510014 184294 510082 184350
rect 510138 184294 540678 184350
rect 540734 184294 540802 184350
rect 540858 184294 571398 184350
rect 571454 184294 571522 184350
rect 571578 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 22422 184226
rect 22478 184170 22546 184226
rect 22602 184170 53142 184226
rect 53198 184170 53266 184226
rect 53322 184170 83862 184226
rect 83918 184170 83986 184226
rect 84042 184170 114582 184226
rect 114638 184170 114706 184226
rect 114762 184170 145302 184226
rect 145358 184170 145426 184226
rect 145482 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 178518 184226
rect 178574 184170 178642 184226
rect 178698 184170 209238 184226
rect 209294 184170 209362 184226
rect 209418 184170 239958 184226
rect 240014 184170 240082 184226
rect 240138 184170 270678 184226
rect 270734 184170 270802 184226
rect 270858 184170 281994 184226
rect 282050 184170 282118 184226
rect 282174 184170 282242 184226
rect 282298 184170 282366 184226
rect 282422 184170 312714 184226
rect 312770 184170 312838 184226
rect 312894 184170 312962 184226
rect 313018 184170 313086 184226
rect 313142 184170 324518 184226
rect 324574 184170 324642 184226
rect 324698 184170 355238 184226
rect 355294 184170 355362 184226
rect 355418 184170 385958 184226
rect 386014 184170 386082 184226
rect 386138 184170 416678 184226
rect 416734 184170 416802 184226
rect 416858 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 448518 184226
rect 448574 184170 448642 184226
rect 448698 184170 479238 184226
rect 479294 184170 479362 184226
rect 479418 184170 509958 184226
rect 510014 184170 510082 184226
rect 510138 184170 540678 184226
rect 540734 184170 540802 184226
rect 540858 184170 571398 184226
rect 571454 184170 571522 184226
rect 571578 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 22422 184102
rect 22478 184046 22546 184102
rect 22602 184046 53142 184102
rect 53198 184046 53266 184102
rect 53322 184046 83862 184102
rect 83918 184046 83986 184102
rect 84042 184046 114582 184102
rect 114638 184046 114706 184102
rect 114762 184046 145302 184102
rect 145358 184046 145426 184102
rect 145482 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 178518 184102
rect 178574 184046 178642 184102
rect 178698 184046 209238 184102
rect 209294 184046 209362 184102
rect 209418 184046 239958 184102
rect 240014 184046 240082 184102
rect 240138 184046 270678 184102
rect 270734 184046 270802 184102
rect 270858 184046 281994 184102
rect 282050 184046 282118 184102
rect 282174 184046 282242 184102
rect 282298 184046 282366 184102
rect 282422 184046 312714 184102
rect 312770 184046 312838 184102
rect 312894 184046 312962 184102
rect 313018 184046 313086 184102
rect 313142 184046 324518 184102
rect 324574 184046 324642 184102
rect 324698 184046 355238 184102
rect 355294 184046 355362 184102
rect 355418 184046 385958 184102
rect 386014 184046 386082 184102
rect 386138 184046 416678 184102
rect 416734 184046 416802 184102
rect 416858 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 448518 184102
rect 448574 184046 448642 184102
rect 448698 184046 479238 184102
rect 479294 184046 479362 184102
rect 479418 184046 509958 184102
rect 510014 184046 510082 184102
rect 510138 184046 540678 184102
rect 540734 184046 540802 184102
rect 540858 184046 571398 184102
rect 571454 184046 571522 184102
rect 571578 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 22422 183978
rect 22478 183922 22546 183978
rect 22602 183922 53142 183978
rect 53198 183922 53266 183978
rect 53322 183922 83862 183978
rect 83918 183922 83986 183978
rect 84042 183922 114582 183978
rect 114638 183922 114706 183978
rect 114762 183922 145302 183978
rect 145358 183922 145426 183978
rect 145482 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 178518 183978
rect 178574 183922 178642 183978
rect 178698 183922 209238 183978
rect 209294 183922 209362 183978
rect 209418 183922 239958 183978
rect 240014 183922 240082 183978
rect 240138 183922 270678 183978
rect 270734 183922 270802 183978
rect 270858 183922 281994 183978
rect 282050 183922 282118 183978
rect 282174 183922 282242 183978
rect 282298 183922 282366 183978
rect 282422 183922 312714 183978
rect 312770 183922 312838 183978
rect 312894 183922 312962 183978
rect 313018 183922 313086 183978
rect 313142 183922 324518 183978
rect 324574 183922 324642 183978
rect 324698 183922 355238 183978
rect 355294 183922 355362 183978
rect 355418 183922 385958 183978
rect 386014 183922 386082 183978
rect 386138 183922 416678 183978
rect 416734 183922 416802 183978
rect 416858 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 448518 183978
rect 448574 183922 448642 183978
rect 448698 183922 479238 183978
rect 479294 183922 479362 183978
rect 479418 183922 509958 183978
rect 510014 183922 510082 183978
rect 510138 183922 540678 183978
rect 540734 183922 540802 183978
rect 540858 183922 571398 183978
rect 571454 183922 571522 183978
rect 571578 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 37782 172350
rect 37838 172294 37906 172350
rect 37962 172294 68502 172350
rect 68558 172294 68626 172350
rect 68682 172294 99222 172350
rect 99278 172294 99346 172350
rect 99402 172294 129942 172350
rect 129998 172294 130066 172350
rect 130122 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 193878 172350
rect 193934 172294 194002 172350
rect 194058 172294 224598 172350
rect 224654 172294 224722 172350
rect 224778 172294 255318 172350
rect 255374 172294 255442 172350
rect 255498 172294 285714 172350
rect 285770 172294 285838 172350
rect 285894 172294 285962 172350
rect 286018 172294 286086 172350
rect 286142 172294 316434 172350
rect 316490 172294 316558 172350
rect 316614 172294 316682 172350
rect 316738 172294 316806 172350
rect 316862 172294 339878 172350
rect 339934 172294 340002 172350
rect 340058 172294 370598 172350
rect 370654 172294 370722 172350
rect 370778 172294 401318 172350
rect 401374 172294 401442 172350
rect 401498 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 463878 172350
rect 463934 172294 464002 172350
rect 464058 172294 494598 172350
rect 494654 172294 494722 172350
rect 494778 172294 525318 172350
rect 525374 172294 525442 172350
rect 525498 172294 556038 172350
rect 556094 172294 556162 172350
rect 556218 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 37782 172226
rect 37838 172170 37906 172226
rect 37962 172170 68502 172226
rect 68558 172170 68626 172226
rect 68682 172170 99222 172226
rect 99278 172170 99346 172226
rect 99402 172170 129942 172226
rect 129998 172170 130066 172226
rect 130122 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 193878 172226
rect 193934 172170 194002 172226
rect 194058 172170 224598 172226
rect 224654 172170 224722 172226
rect 224778 172170 255318 172226
rect 255374 172170 255442 172226
rect 255498 172170 285714 172226
rect 285770 172170 285838 172226
rect 285894 172170 285962 172226
rect 286018 172170 286086 172226
rect 286142 172170 316434 172226
rect 316490 172170 316558 172226
rect 316614 172170 316682 172226
rect 316738 172170 316806 172226
rect 316862 172170 339878 172226
rect 339934 172170 340002 172226
rect 340058 172170 370598 172226
rect 370654 172170 370722 172226
rect 370778 172170 401318 172226
rect 401374 172170 401442 172226
rect 401498 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 463878 172226
rect 463934 172170 464002 172226
rect 464058 172170 494598 172226
rect 494654 172170 494722 172226
rect 494778 172170 525318 172226
rect 525374 172170 525442 172226
rect 525498 172170 556038 172226
rect 556094 172170 556162 172226
rect 556218 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 37782 172102
rect 37838 172046 37906 172102
rect 37962 172046 68502 172102
rect 68558 172046 68626 172102
rect 68682 172046 99222 172102
rect 99278 172046 99346 172102
rect 99402 172046 129942 172102
rect 129998 172046 130066 172102
rect 130122 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 193878 172102
rect 193934 172046 194002 172102
rect 194058 172046 224598 172102
rect 224654 172046 224722 172102
rect 224778 172046 255318 172102
rect 255374 172046 255442 172102
rect 255498 172046 285714 172102
rect 285770 172046 285838 172102
rect 285894 172046 285962 172102
rect 286018 172046 286086 172102
rect 286142 172046 316434 172102
rect 316490 172046 316558 172102
rect 316614 172046 316682 172102
rect 316738 172046 316806 172102
rect 316862 172046 339878 172102
rect 339934 172046 340002 172102
rect 340058 172046 370598 172102
rect 370654 172046 370722 172102
rect 370778 172046 401318 172102
rect 401374 172046 401442 172102
rect 401498 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 463878 172102
rect 463934 172046 464002 172102
rect 464058 172046 494598 172102
rect 494654 172046 494722 172102
rect 494778 172046 525318 172102
rect 525374 172046 525442 172102
rect 525498 172046 556038 172102
rect 556094 172046 556162 172102
rect 556218 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 37782 171978
rect 37838 171922 37906 171978
rect 37962 171922 68502 171978
rect 68558 171922 68626 171978
rect 68682 171922 99222 171978
rect 99278 171922 99346 171978
rect 99402 171922 129942 171978
rect 129998 171922 130066 171978
rect 130122 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 193878 171978
rect 193934 171922 194002 171978
rect 194058 171922 224598 171978
rect 224654 171922 224722 171978
rect 224778 171922 255318 171978
rect 255374 171922 255442 171978
rect 255498 171922 285714 171978
rect 285770 171922 285838 171978
rect 285894 171922 285962 171978
rect 286018 171922 286086 171978
rect 286142 171922 316434 171978
rect 316490 171922 316558 171978
rect 316614 171922 316682 171978
rect 316738 171922 316806 171978
rect 316862 171922 339878 171978
rect 339934 171922 340002 171978
rect 340058 171922 370598 171978
rect 370654 171922 370722 171978
rect 370778 171922 401318 171978
rect 401374 171922 401442 171978
rect 401498 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 463878 171978
rect 463934 171922 464002 171978
rect 464058 171922 494598 171978
rect 494654 171922 494722 171978
rect 494778 171922 525318 171978
rect 525374 171922 525442 171978
rect 525498 171922 556038 171978
rect 556094 171922 556162 171978
rect 556218 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 22422 166350
rect 22478 166294 22546 166350
rect 22602 166294 53142 166350
rect 53198 166294 53266 166350
rect 53322 166294 83862 166350
rect 83918 166294 83986 166350
rect 84042 166294 114582 166350
rect 114638 166294 114706 166350
rect 114762 166294 145302 166350
rect 145358 166294 145426 166350
rect 145482 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 178518 166350
rect 178574 166294 178642 166350
rect 178698 166294 209238 166350
rect 209294 166294 209362 166350
rect 209418 166294 239958 166350
rect 240014 166294 240082 166350
rect 240138 166294 270678 166350
rect 270734 166294 270802 166350
rect 270858 166294 281994 166350
rect 282050 166294 282118 166350
rect 282174 166294 282242 166350
rect 282298 166294 282366 166350
rect 282422 166294 312714 166350
rect 312770 166294 312838 166350
rect 312894 166294 312962 166350
rect 313018 166294 313086 166350
rect 313142 166294 324518 166350
rect 324574 166294 324642 166350
rect 324698 166294 355238 166350
rect 355294 166294 355362 166350
rect 355418 166294 385958 166350
rect 386014 166294 386082 166350
rect 386138 166294 416678 166350
rect 416734 166294 416802 166350
rect 416858 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 448518 166350
rect 448574 166294 448642 166350
rect 448698 166294 479238 166350
rect 479294 166294 479362 166350
rect 479418 166294 509958 166350
rect 510014 166294 510082 166350
rect 510138 166294 540678 166350
rect 540734 166294 540802 166350
rect 540858 166294 571398 166350
rect 571454 166294 571522 166350
rect 571578 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 22422 166226
rect 22478 166170 22546 166226
rect 22602 166170 53142 166226
rect 53198 166170 53266 166226
rect 53322 166170 83862 166226
rect 83918 166170 83986 166226
rect 84042 166170 114582 166226
rect 114638 166170 114706 166226
rect 114762 166170 145302 166226
rect 145358 166170 145426 166226
rect 145482 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 178518 166226
rect 178574 166170 178642 166226
rect 178698 166170 209238 166226
rect 209294 166170 209362 166226
rect 209418 166170 239958 166226
rect 240014 166170 240082 166226
rect 240138 166170 270678 166226
rect 270734 166170 270802 166226
rect 270858 166170 281994 166226
rect 282050 166170 282118 166226
rect 282174 166170 282242 166226
rect 282298 166170 282366 166226
rect 282422 166170 312714 166226
rect 312770 166170 312838 166226
rect 312894 166170 312962 166226
rect 313018 166170 313086 166226
rect 313142 166170 324518 166226
rect 324574 166170 324642 166226
rect 324698 166170 355238 166226
rect 355294 166170 355362 166226
rect 355418 166170 385958 166226
rect 386014 166170 386082 166226
rect 386138 166170 416678 166226
rect 416734 166170 416802 166226
rect 416858 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 448518 166226
rect 448574 166170 448642 166226
rect 448698 166170 479238 166226
rect 479294 166170 479362 166226
rect 479418 166170 509958 166226
rect 510014 166170 510082 166226
rect 510138 166170 540678 166226
rect 540734 166170 540802 166226
rect 540858 166170 571398 166226
rect 571454 166170 571522 166226
rect 571578 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 22422 166102
rect 22478 166046 22546 166102
rect 22602 166046 53142 166102
rect 53198 166046 53266 166102
rect 53322 166046 83862 166102
rect 83918 166046 83986 166102
rect 84042 166046 114582 166102
rect 114638 166046 114706 166102
rect 114762 166046 145302 166102
rect 145358 166046 145426 166102
rect 145482 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 178518 166102
rect 178574 166046 178642 166102
rect 178698 166046 209238 166102
rect 209294 166046 209362 166102
rect 209418 166046 239958 166102
rect 240014 166046 240082 166102
rect 240138 166046 270678 166102
rect 270734 166046 270802 166102
rect 270858 166046 281994 166102
rect 282050 166046 282118 166102
rect 282174 166046 282242 166102
rect 282298 166046 282366 166102
rect 282422 166046 312714 166102
rect 312770 166046 312838 166102
rect 312894 166046 312962 166102
rect 313018 166046 313086 166102
rect 313142 166046 324518 166102
rect 324574 166046 324642 166102
rect 324698 166046 355238 166102
rect 355294 166046 355362 166102
rect 355418 166046 385958 166102
rect 386014 166046 386082 166102
rect 386138 166046 416678 166102
rect 416734 166046 416802 166102
rect 416858 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 448518 166102
rect 448574 166046 448642 166102
rect 448698 166046 479238 166102
rect 479294 166046 479362 166102
rect 479418 166046 509958 166102
rect 510014 166046 510082 166102
rect 510138 166046 540678 166102
rect 540734 166046 540802 166102
rect 540858 166046 571398 166102
rect 571454 166046 571522 166102
rect 571578 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 22422 165978
rect 22478 165922 22546 165978
rect 22602 165922 53142 165978
rect 53198 165922 53266 165978
rect 53322 165922 83862 165978
rect 83918 165922 83986 165978
rect 84042 165922 114582 165978
rect 114638 165922 114706 165978
rect 114762 165922 145302 165978
rect 145358 165922 145426 165978
rect 145482 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 178518 165978
rect 178574 165922 178642 165978
rect 178698 165922 209238 165978
rect 209294 165922 209362 165978
rect 209418 165922 239958 165978
rect 240014 165922 240082 165978
rect 240138 165922 270678 165978
rect 270734 165922 270802 165978
rect 270858 165922 281994 165978
rect 282050 165922 282118 165978
rect 282174 165922 282242 165978
rect 282298 165922 282366 165978
rect 282422 165922 312714 165978
rect 312770 165922 312838 165978
rect 312894 165922 312962 165978
rect 313018 165922 313086 165978
rect 313142 165922 324518 165978
rect 324574 165922 324642 165978
rect 324698 165922 355238 165978
rect 355294 165922 355362 165978
rect 355418 165922 385958 165978
rect 386014 165922 386082 165978
rect 386138 165922 416678 165978
rect 416734 165922 416802 165978
rect 416858 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 448518 165978
rect 448574 165922 448642 165978
rect 448698 165922 479238 165978
rect 479294 165922 479362 165978
rect 479418 165922 509958 165978
rect 510014 165922 510082 165978
rect 510138 165922 540678 165978
rect 540734 165922 540802 165978
rect 540858 165922 571398 165978
rect 571454 165922 571522 165978
rect 571578 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 37782 154350
rect 37838 154294 37906 154350
rect 37962 154294 68502 154350
rect 68558 154294 68626 154350
rect 68682 154294 99222 154350
rect 99278 154294 99346 154350
rect 99402 154294 129942 154350
rect 129998 154294 130066 154350
rect 130122 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 193878 154350
rect 193934 154294 194002 154350
rect 194058 154294 224598 154350
rect 224654 154294 224722 154350
rect 224778 154294 255318 154350
rect 255374 154294 255442 154350
rect 255498 154294 285714 154350
rect 285770 154294 285838 154350
rect 285894 154294 285962 154350
rect 286018 154294 286086 154350
rect 286142 154294 316434 154350
rect 316490 154294 316558 154350
rect 316614 154294 316682 154350
rect 316738 154294 316806 154350
rect 316862 154294 339878 154350
rect 339934 154294 340002 154350
rect 340058 154294 370598 154350
rect 370654 154294 370722 154350
rect 370778 154294 401318 154350
rect 401374 154294 401442 154350
rect 401498 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 463878 154350
rect 463934 154294 464002 154350
rect 464058 154294 494598 154350
rect 494654 154294 494722 154350
rect 494778 154294 525318 154350
rect 525374 154294 525442 154350
rect 525498 154294 556038 154350
rect 556094 154294 556162 154350
rect 556218 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 37782 154226
rect 37838 154170 37906 154226
rect 37962 154170 68502 154226
rect 68558 154170 68626 154226
rect 68682 154170 99222 154226
rect 99278 154170 99346 154226
rect 99402 154170 129942 154226
rect 129998 154170 130066 154226
rect 130122 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 193878 154226
rect 193934 154170 194002 154226
rect 194058 154170 224598 154226
rect 224654 154170 224722 154226
rect 224778 154170 255318 154226
rect 255374 154170 255442 154226
rect 255498 154170 285714 154226
rect 285770 154170 285838 154226
rect 285894 154170 285962 154226
rect 286018 154170 286086 154226
rect 286142 154170 316434 154226
rect 316490 154170 316558 154226
rect 316614 154170 316682 154226
rect 316738 154170 316806 154226
rect 316862 154170 339878 154226
rect 339934 154170 340002 154226
rect 340058 154170 370598 154226
rect 370654 154170 370722 154226
rect 370778 154170 401318 154226
rect 401374 154170 401442 154226
rect 401498 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 463878 154226
rect 463934 154170 464002 154226
rect 464058 154170 494598 154226
rect 494654 154170 494722 154226
rect 494778 154170 525318 154226
rect 525374 154170 525442 154226
rect 525498 154170 556038 154226
rect 556094 154170 556162 154226
rect 556218 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 37782 154102
rect 37838 154046 37906 154102
rect 37962 154046 68502 154102
rect 68558 154046 68626 154102
rect 68682 154046 99222 154102
rect 99278 154046 99346 154102
rect 99402 154046 129942 154102
rect 129998 154046 130066 154102
rect 130122 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 193878 154102
rect 193934 154046 194002 154102
rect 194058 154046 224598 154102
rect 224654 154046 224722 154102
rect 224778 154046 255318 154102
rect 255374 154046 255442 154102
rect 255498 154046 285714 154102
rect 285770 154046 285838 154102
rect 285894 154046 285962 154102
rect 286018 154046 286086 154102
rect 286142 154046 316434 154102
rect 316490 154046 316558 154102
rect 316614 154046 316682 154102
rect 316738 154046 316806 154102
rect 316862 154046 339878 154102
rect 339934 154046 340002 154102
rect 340058 154046 370598 154102
rect 370654 154046 370722 154102
rect 370778 154046 401318 154102
rect 401374 154046 401442 154102
rect 401498 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 463878 154102
rect 463934 154046 464002 154102
rect 464058 154046 494598 154102
rect 494654 154046 494722 154102
rect 494778 154046 525318 154102
rect 525374 154046 525442 154102
rect 525498 154046 556038 154102
rect 556094 154046 556162 154102
rect 556218 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 37782 153978
rect 37838 153922 37906 153978
rect 37962 153922 68502 153978
rect 68558 153922 68626 153978
rect 68682 153922 99222 153978
rect 99278 153922 99346 153978
rect 99402 153922 129942 153978
rect 129998 153922 130066 153978
rect 130122 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 193878 153978
rect 193934 153922 194002 153978
rect 194058 153922 224598 153978
rect 224654 153922 224722 153978
rect 224778 153922 255318 153978
rect 255374 153922 255442 153978
rect 255498 153922 285714 153978
rect 285770 153922 285838 153978
rect 285894 153922 285962 153978
rect 286018 153922 286086 153978
rect 286142 153922 316434 153978
rect 316490 153922 316558 153978
rect 316614 153922 316682 153978
rect 316738 153922 316806 153978
rect 316862 153922 339878 153978
rect 339934 153922 340002 153978
rect 340058 153922 370598 153978
rect 370654 153922 370722 153978
rect 370778 153922 401318 153978
rect 401374 153922 401442 153978
rect 401498 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 463878 153978
rect 463934 153922 464002 153978
rect 464058 153922 494598 153978
rect 494654 153922 494722 153978
rect 494778 153922 525318 153978
rect 525374 153922 525442 153978
rect 525498 153922 556038 153978
rect 556094 153922 556162 153978
rect 556218 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 22422 148350
rect 22478 148294 22546 148350
rect 22602 148294 53142 148350
rect 53198 148294 53266 148350
rect 53322 148294 83862 148350
rect 83918 148294 83986 148350
rect 84042 148294 114582 148350
rect 114638 148294 114706 148350
rect 114762 148294 145302 148350
rect 145358 148294 145426 148350
rect 145482 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 178518 148350
rect 178574 148294 178642 148350
rect 178698 148294 209238 148350
rect 209294 148294 209362 148350
rect 209418 148294 239958 148350
rect 240014 148294 240082 148350
rect 240138 148294 270678 148350
rect 270734 148294 270802 148350
rect 270858 148294 281994 148350
rect 282050 148294 282118 148350
rect 282174 148294 282242 148350
rect 282298 148294 282366 148350
rect 282422 148294 312714 148350
rect 312770 148294 312838 148350
rect 312894 148294 312962 148350
rect 313018 148294 313086 148350
rect 313142 148294 324518 148350
rect 324574 148294 324642 148350
rect 324698 148294 355238 148350
rect 355294 148294 355362 148350
rect 355418 148294 385958 148350
rect 386014 148294 386082 148350
rect 386138 148294 416678 148350
rect 416734 148294 416802 148350
rect 416858 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 448518 148350
rect 448574 148294 448642 148350
rect 448698 148294 479238 148350
rect 479294 148294 479362 148350
rect 479418 148294 509958 148350
rect 510014 148294 510082 148350
rect 510138 148294 540678 148350
rect 540734 148294 540802 148350
rect 540858 148294 571398 148350
rect 571454 148294 571522 148350
rect 571578 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 22422 148226
rect 22478 148170 22546 148226
rect 22602 148170 53142 148226
rect 53198 148170 53266 148226
rect 53322 148170 83862 148226
rect 83918 148170 83986 148226
rect 84042 148170 114582 148226
rect 114638 148170 114706 148226
rect 114762 148170 145302 148226
rect 145358 148170 145426 148226
rect 145482 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 178518 148226
rect 178574 148170 178642 148226
rect 178698 148170 209238 148226
rect 209294 148170 209362 148226
rect 209418 148170 239958 148226
rect 240014 148170 240082 148226
rect 240138 148170 270678 148226
rect 270734 148170 270802 148226
rect 270858 148170 281994 148226
rect 282050 148170 282118 148226
rect 282174 148170 282242 148226
rect 282298 148170 282366 148226
rect 282422 148170 312714 148226
rect 312770 148170 312838 148226
rect 312894 148170 312962 148226
rect 313018 148170 313086 148226
rect 313142 148170 324518 148226
rect 324574 148170 324642 148226
rect 324698 148170 355238 148226
rect 355294 148170 355362 148226
rect 355418 148170 385958 148226
rect 386014 148170 386082 148226
rect 386138 148170 416678 148226
rect 416734 148170 416802 148226
rect 416858 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 448518 148226
rect 448574 148170 448642 148226
rect 448698 148170 479238 148226
rect 479294 148170 479362 148226
rect 479418 148170 509958 148226
rect 510014 148170 510082 148226
rect 510138 148170 540678 148226
rect 540734 148170 540802 148226
rect 540858 148170 571398 148226
rect 571454 148170 571522 148226
rect 571578 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 22422 148102
rect 22478 148046 22546 148102
rect 22602 148046 53142 148102
rect 53198 148046 53266 148102
rect 53322 148046 83862 148102
rect 83918 148046 83986 148102
rect 84042 148046 114582 148102
rect 114638 148046 114706 148102
rect 114762 148046 145302 148102
rect 145358 148046 145426 148102
rect 145482 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 178518 148102
rect 178574 148046 178642 148102
rect 178698 148046 209238 148102
rect 209294 148046 209362 148102
rect 209418 148046 239958 148102
rect 240014 148046 240082 148102
rect 240138 148046 270678 148102
rect 270734 148046 270802 148102
rect 270858 148046 281994 148102
rect 282050 148046 282118 148102
rect 282174 148046 282242 148102
rect 282298 148046 282366 148102
rect 282422 148046 312714 148102
rect 312770 148046 312838 148102
rect 312894 148046 312962 148102
rect 313018 148046 313086 148102
rect 313142 148046 324518 148102
rect 324574 148046 324642 148102
rect 324698 148046 355238 148102
rect 355294 148046 355362 148102
rect 355418 148046 385958 148102
rect 386014 148046 386082 148102
rect 386138 148046 416678 148102
rect 416734 148046 416802 148102
rect 416858 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 448518 148102
rect 448574 148046 448642 148102
rect 448698 148046 479238 148102
rect 479294 148046 479362 148102
rect 479418 148046 509958 148102
rect 510014 148046 510082 148102
rect 510138 148046 540678 148102
rect 540734 148046 540802 148102
rect 540858 148046 571398 148102
rect 571454 148046 571522 148102
rect 571578 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 22422 147978
rect 22478 147922 22546 147978
rect 22602 147922 53142 147978
rect 53198 147922 53266 147978
rect 53322 147922 83862 147978
rect 83918 147922 83986 147978
rect 84042 147922 114582 147978
rect 114638 147922 114706 147978
rect 114762 147922 145302 147978
rect 145358 147922 145426 147978
rect 145482 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 178518 147978
rect 178574 147922 178642 147978
rect 178698 147922 209238 147978
rect 209294 147922 209362 147978
rect 209418 147922 239958 147978
rect 240014 147922 240082 147978
rect 240138 147922 270678 147978
rect 270734 147922 270802 147978
rect 270858 147922 281994 147978
rect 282050 147922 282118 147978
rect 282174 147922 282242 147978
rect 282298 147922 282366 147978
rect 282422 147922 312714 147978
rect 312770 147922 312838 147978
rect 312894 147922 312962 147978
rect 313018 147922 313086 147978
rect 313142 147922 324518 147978
rect 324574 147922 324642 147978
rect 324698 147922 355238 147978
rect 355294 147922 355362 147978
rect 355418 147922 385958 147978
rect 386014 147922 386082 147978
rect 386138 147922 416678 147978
rect 416734 147922 416802 147978
rect 416858 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 448518 147978
rect 448574 147922 448642 147978
rect 448698 147922 479238 147978
rect 479294 147922 479362 147978
rect 479418 147922 509958 147978
rect 510014 147922 510082 147978
rect 510138 147922 540678 147978
rect 540734 147922 540802 147978
rect 540858 147922 571398 147978
rect 571454 147922 571522 147978
rect 571578 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 37782 136350
rect 37838 136294 37906 136350
rect 37962 136294 68502 136350
rect 68558 136294 68626 136350
rect 68682 136294 99222 136350
rect 99278 136294 99346 136350
rect 99402 136294 129942 136350
rect 129998 136294 130066 136350
rect 130122 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 193878 136350
rect 193934 136294 194002 136350
rect 194058 136294 224598 136350
rect 224654 136294 224722 136350
rect 224778 136294 255318 136350
rect 255374 136294 255442 136350
rect 255498 136294 285714 136350
rect 285770 136294 285838 136350
rect 285894 136294 285962 136350
rect 286018 136294 286086 136350
rect 286142 136294 316434 136350
rect 316490 136294 316558 136350
rect 316614 136294 316682 136350
rect 316738 136294 316806 136350
rect 316862 136294 339878 136350
rect 339934 136294 340002 136350
rect 340058 136294 370598 136350
rect 370654 136294 370722 136350
rect 370778 136294 401318 136350
rect 401374 136294 401442 136350
rect 401498 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 463878 136350
rect 463934 136294 464002 136350
rect 464058 136294 494598 136350
rect 494654 136294 494722 136350
rect 494778 136294 525318 136350
rect 525374 136294 525442 136350
rect 525498 136294 556038 136350
rect 556094 136294 556162 136350
rect 556218 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 37782 136226
rect 37838 136170 37906 136226
rect 37962 136170 68502 136226
rect 68558 136170 68626 136226
rect 68682 136170 99222 136226
rect 99278 136170 99346 136226
rect 99402 136170 129942 136226
rect 129998 136170 130066 136226
rect 130122 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 193878 136226
rect 193934 136170 194002 136226
rect 194058 136170 224598 136226
rect 224654 136170 224722 136226
rect 224778 136170 255318 136226
rect 255374 136170 255442 136226
rect 255498 136170 285714 136226
rect 285770 136170 285838 136226
rect 285894 136170 285962 136226
rect 286018 136170 286086 136226
rect 286142 136170 316434 136226
rect 316490 136170 316558 136226
rect 316614 136170 316682 136226
rect 316738 136170 316806 136226
rect 316862 136170 339878 136226
rect 339934 136170 340002 136226
rect 340058 136170 370598 136226
rect 370654 136170 370722 136226
rect 370778 136170 401318 136226
rect 401374 136170 401442 136226
rect 401498 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 463878 136226
rect 463934 136170 464002 136226
rect 464058 136170 494598 136226
rect 494654 136170 494722 136226
rect 494778 136170 525318 136226
rect 525374 136170 525442 136226
rect 525498 136170 556038 136226
rect 556094 136170 556162 136226
rect 556218 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 37782 136102
rect 37838 136046 37906 136102
rect 37962 136046 68502 136102
rect 68558 136046 68626 136102
rect 68682 136046 99222 136102
rect 99278 136046 99346 136102
rect 99402 136046 129942 136102
rect 129998 136046 130066 136102
rect 130122 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 193878 136102
rect 193934 136046 194002 136102
rect 194058 136046 224598 136102
rect 224654 136046 224722 136102
rect 224778 136046 255318 136102
rect 255374 136046 255442 136102
rect 255498 136046 285714 136102
rect 285770 136046 285838 136102
rect 285894 136046 285962 136102
rect 286018 136046 286086 136102
rect 286142 136046 316434 136102
rect 316490 136046 316558 136102
rect 316614 136046 316682 136102
rect 316738 136046 316806 136102
rect 316862 136046 339878 136102
rect 339934 136046 340002 136102
rect 340058 136046 370598 136102
rect 370654 136046 370722 136102
rect 370778 136046 401318 136102
rect 401374 136046 401442 136102
rect 401498 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 463878 136102
rect 463934 136046 464002 136102
rect 464058 136046 494598 136102
rect 494654 136046 494722 136102
rect 494778 136046 525318 136102
rect 525374 136046 525442 136102
rect 525498 136046 556038 136102
rect 556094 136046 556162 136102
rect 556218 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 37782 135978
rect 37838 135922 37906 135978
rect 37962 135922 68502 135978
rect 68558 135922 68626 135978
rect 68682 135922 99222 135978
rect 99278 135922 99346 135978
rect 99402 135922 129942 135978
rect 129998 135922 130066 135978
rect 130122 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 193878 135978
rect 193934 135922 194002 135978
rect 194058 135922 224598 135978
rect 224654 135922 224722 135978
rect 224778 135922 255318 135978
rect 255374 135922 255442 135978
rect 255498 135922 285714 135978
rect 285770 135922 285838 135978
rect 285894 135922 285962 135978
rect 286018 135922 286086 135978
rect 286142 135922 316434 135978
rect 316490 135922 316558 135978
rect 316614 135922 316682 135978
rect 316738 135922 316806 135978
rect 316862 135922 339878 135978
rect 339934 135922 340002 135978
rect 340058 135922 370598 135978
rect 370654 135922 370722 135978
rect 370778 135922 401318 135978
rect 401374 135922 401442 135978
rect 401498 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 463878 135978
rect 463934 135922 464002 135978
rect 464058 135922 494598 135978
rect 494654 135922 494722 135978
rect 494778 135922 525318 135978
rect 525374 135922 525442 135978
rect 525498 135922 556038 135978
rect 556094 135922 556162 135978
rect 556218 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 22422 130350
rect 22478 130294 22546 130350
rect 22602 130294 53142 130350
rect 53198 130294 53266 130350
rect 53322 130294 83862 130350
rect 83918 130294 83986 130350
rect 84042 130294 114582 130350
rect 114638 130294 114706 130350
rect 114762 130294 145302 130350
rect 145358 130294 145426 130350
rect 145482 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 178518 130350
rect 178574 130294 178642 130350
rect 178698 130294 209238 130350
rect 209294 130294 209362 130350
rect 209418 130294 239958 130350
rect 240014 130294 240082 130350
rect 240138 130294 270678 130350
rect 270734 130294 270802 130350
rect 270858 130294 281994 130350
rect 282050 130294 282118 130350
rect 282174 130294 282242 130350
rect 282298 130294 282366 130350
rect 282422 130294 312714 130350
rect 312770 130294 312838 130350
rect 312894 130294 312962 130350
rect 313018 130294 313086 130350
rect 313142 130294 324518 130350
rect 324574 130294 324642 130350
rect 324698 130294 355238 130350
rect 355294 130294 355362 130350
rect 355418 130294 385958 130350
rect 386014 130294 386082 130350
rect 386138 130294 416678 130350
rect 416734 130294 416802 130350
rect 416858 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 448518 130350
rect 448574 130294 448642 130350
rect 448698 130294 479238 130350
rect 479294 130294 479362 130350
rect 479418 130294 509958 130350
rect 510014 130294 510082 130350
rect 510138 130294 540678 130350
rect 540734 130294 540802 130350
rect 540858 130294 571398 130350
rect 571454 130294 571522 130350
rect 571578 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 22422 130226
rect 22478 130170 22546 130226
rect 22602 130170 53142 130226
rect 53198 130170 53266 130226
rect 53322 130170 83862 130226
rect 83918 130170 83986 130226
rect 84042 130170 114582 130226
rect 114638 130170 114706 130226
rect 114762 130170 145302 130226
rect 145358 130170 145426 130226
rect 145482 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 178518 130226
rect 178574 130170 178642 130226
rect 178698 130170 209238 130226
rect 209294 130170 209362 130226
rect 209418 130170 239958 130226
rect 240014 130170 240082 130226
rect 240138 130170 270678 130226
rect 270734 130170 270802 130226
rect 270858 130170 281994 130226
rect 282050 130170 282118 130226
rect 282174 130170 282242 130226
rect 282298 130170 282366 130226
rect 282422 130170 312714 130226
rect 312770 130170 312838 130226
rect 312894 130170 312962 130226
rect 313018 130170 313086 130226
rect 313142 130170 324518 130226
rect 324574 130170 324642 130226
rect 324698 130170 355238 130226
rect 355294 130170 355362 130226
rect 355418 130170 385958 130226
rect 386014 130170 386082 130226
rect 386138 130170 416678 130226
rect 416734 130170 416802 130226
rect 416858 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 448518 130226
rect 448574 130170 448642 130226
rect 448698 130170 479238 130226
rect 479294 130170 479362 130226
rect 479418 130170 509958 130226
rect 510014 130170 510082 130226
rect 510138 130170 540678 130226
rect 540734 130170 540802 130226
rect 540858 130170 571398 130226
rect 571454 130170 571522 130226
rect 571578 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 22422 130102
rect 22478 130046 22546 130102
rect 22602 130046 53142 130102
rect 53198 130046 53266 130102
rect 53322 130046 83862 130102
rect 83918 130046 83986 130102
rect 84042 130046 114582 130102
rect 114638 130046 114706 130102
rect 114762 130046 145302 130102
rect 145358 130046 145426 130102
rect 145482 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 178518 130102
rect 178574 130046 178642 130102
rect 178698 130046 209238 130102
rect 209294 130046 209362 130102
rect 209418 130046 239958 130102
rect 240014 130046 240082 130102
rect 240138 130046 270678 130102
rect 270734 130046 270802 130102
rect 270858 130046 281994 130102
rect 282050 130046 282118 130102
rect 282174 130046 282242 130102
rect 282298 130046 282366 130102
rect 282422 130046 312714 130102
rect 312770 130046 312838 130102
rect 312894 130046 312962 130102
rect 313018 130046 313086 130102
rect 313142 130046 324518 130102
rect 324574 130046 324642 130102
rect 324698 130046 355238 130102
rect 355294 130046 355362 130102
rect 355418 130046 385958 130102
rect 386014 130046 386082 130102
rect 386138 130046 416678 130102
rect 416734 130046 416802 130102
rect 416858 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 448518 130102
rect 448574 130046 448642 130102
rect 448698 130046 479238 130102
rect 479294 130046 479362 130102
rect 479418 130046 509958 130102
rect 510014 130046 510082 130102
rect 510138 130046 540678 130102
rect 540734 130046 540802 130102
rect 540858 130046 571398 130102
rect 571454 130046 571522 130102
rect 571578 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 22422 129978
rect 22478 129922 22546 129978
rect 22602 129922 53142 129978
rect 53198 129922 53266 129978
rect 53322 129922 83862 129978
rect 83918 129922 83986 129978
rect 84042 129922 114582 129978
rect 114638 129922 114706 129978
rect 114762 129922 145302 129978
rect 145358 129922 145426 129978
rect 145482 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 178518 129978
rect 178574 129922 178642 129978
rect 178698 129922 209238 129978
rect 209294 129922 209362 129978
rect 209418 129922 239958 129978
rect 240014 129922 240082 129978
rect 240138 129922 270678 129978
rect 270734 129922 270802 129978
rect 270858 129922 281994 129978
rect 282050 129922 282118 129978
rect 282174 129922 282242 129978
rect 282298 129922 282366 129978
rect 282422 129922 312714 129978
rect 312770 129922 312838 129978
rect 312894 129922 312962 129978
rect 313018 129922 313086 129978
rect 313142 129922 324518 129978
rect 324574 129922 324642 129978
rect 324698 129922 355238 129978
rect 355294 129922 355362 129978
rect 355418 129922 385958 129978
rect 386014 129922 386082 129978
rect 386138 129922 416678 129978
rect 416734 129922 416802 129978
rect 416858 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 448518 129978
rect 448574 129922 448642 129978
rect 448698 129922 479238 129978
rect 479294 129922 479362 129978
rect 479418 129922 509958 129978
rect 510014 129922 510082 129978
rect 510138 129922 540678 129978
rect 540734 129922 540802 129978
rect 540858 129922 571398 129978
rect 571454 129922 571522 129978
rect 571578 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 37782 118350
rect 37838 118294 37906 118350
rect 37962 118294 68502 118350
rect 68558 118294 68626 118350
rect 68682 118294 99222 118350
rect 99278 118294 99346 118350
rect 99402 118294 129942 118350
rect 129998 118294 130066 118350
rect 130122 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 193878 118350
rect 193934 118294 194002 118350
rect 194058 118294 224598 118350
rect 224654 118294 224722 118350
rect 224778 118294 255318 118350
rect 255374 118294 255442 118350
rect 255498 118294 285714 118350
rect 285770 118294 285838 118350
rect 285894 118294 285962 118350
rect 286018 118294 286086 118350
rect 286142 118294 316434 118350
rect 316490 118294 316558 118350
rect 316614 118294 316682 118350
rect 316738 118294 316806 118350
rect 316862 118294 339878 118350
rect 339934 118294 340002 118350
rect 340058 118294 370598 118350
rect 370654 118294 370722 118350
rect 370778 118294 401318 118350
rect 401374 118294 401442 118350
rect 401498 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 463878 118350
rect 463934 118294 464002 118350
rect 464058 118294 494598 118350
rect 494654 118294 494722 118350
rect 494778 118294 525318 118350
rect 525374 118294 525442 118350
rect 525498 118294 556038 118350
rect 556094 118294 556162 118350
rect 556218 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 37782 118226
rect 37838 118170 37906 118226
rect 37962 118170 68502 118226
rect 68558 118170 68626 118226
rect 68682 118170 99222 118226
rect 99278 118170 99346 118226
rect 99402 118170 129942 118226
rect 129998 118170 130066 118226
rect 130122 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 193878 118226
rect 193934 118170 194002 118226
rect 194058 118170 224598 118226
rect 224654 118170 224722 118226
rect 224778 118170 255318 118226
rect 255374 118170 255442 118226
rect 255498 118170 285714 118226
rect 285770 118170 285838 118226
rect 285894 118170 285962 118226
rect 286018 118170 286086 118226
rect 286142 118170 316434 118226
rect 316490 118170 316558 118226
rect 316614 118170 316682 118226
rect 316738 118170 316806 118226
rect 316862 118170 339878 118226
rect 339934 118170 340002 118226
rect 340058 118170 370598 118226
rect 370654 118170 370722 118226
rect 370778 118170 401318 118226
rect 401374 118170 401442 118226
rect 401498 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 463878 118226
rect 463934 118170 464002 118226
rect 464058 118170 494598 118226
rect 494654 118170 494722 118226
rect 494778 118170 525318 118226
rect 525374 118170 525442 118226
rect 525498 118170 556038 118226
rect 556094 118170 556162 118226
rect 556218 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 37782 118102
rect 37838 118046 37906 118102
rect 37962 118046 68502 118102
rect 68558 118046 68626 118102
rect 68682 118046 99222 118102
rect 99278 118046 99346 118102
rect 99402 118046 129942 118102
rect 129998 118046 130066 118102
rect 130122 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 193878 118102
rect 193934 118046 194002 118102
rect 194058 118046 224598 118102
rect 224654 118046 224722 118102
rect 224778 118046 255318 118102
rect 255374 118046 255442 118102
rect 255498 118046 285714 118102
rect 285770 118046 285838 118102
rect 285894 118046 285962 118102
rect 286018 118046 286086 118102
rect 286142 118046 316434 118102
rect 316490 118046 316558 118102
rect 316614 118046 316682 118102
rect 316738 118046 316806 118102
rect 316862 118046 339878 118102
rect 339934 118046 340002 118102
rect 340058 118046 370598 118102
rect 370654 118046 370722 118102
rect 370778 118046 401318 118102
rect 401374 118046 401442 118102
rect 401498 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 463878 118102
rect 463934 118046 464002 118102
rect 464058 118046 494598 118102
rect 494654 118046 494722 118102
rect 494778 118046 525318 118102
rect 525374 118046 525442 118102
rect 525498 118046 556038 118102
rect 556094 118046 556162 118102
rect 556218 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 37782 117978
rect 37838 117922 37906 117978
rect 37962 117922 68502 117978
rect 68558 117922 68626 117978
rect 68682 117922 99222 117978
rect 99278 117922 99346 117978
rect 99402 117922 129942 117978
rect 129998 117922 130066 117978
rect 130122 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 193878 117978
rect 193934 117922 194002 117978
rect 194058 117922 224598 117978
rect 224654 117922 224722 117978
rect 224778 117922 255318 117978
rect 255374 117922 255442 117978
rect 255498 117922 285714 117978
rect 285770 117922 285838 117978
rect 285894 117922 285962 117978
rect 286018 117922 286086 117978
rect 286142 117922 316434 117978
rect 316490 117922 316558 117978
rect 316614 117922 316682 117978
rect 316738 117922 316806 117978
rect 316862 117922 339878 117978
rect 339934 117922 340002 117978
rect 340058 117922 370598 117978
rect 370654 117922 370722 117978
rect 370778 117922 401318 117978
rect 401374 117922 401442 117978
rect 401498 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 463878 117978
rect 463934 117922 464002 117978
rect 464058 117922 494598 117978
rect 494654 117922 494722 117978
rect 494778 117922 525318 117978
rect 525374 117922 525442 117978
rect 525498 117922 556038 117978
rect 556094 117922 556162 117978
rect 556218 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 22422 112350
rect 22478 112294 22546 112350
rect 22602 112294 53142 112350
rect 53198 112294 53266 112350
rect 53322 112294 83862 112350
rect 83918 112294 83986 112350
rect 84042 112294 114582 112350
rect 114638 112294 114706 112350
rect 114762 112294 145302 112350
rect 145358 112294 145426 112350
rect 145482 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 178518 112350
rect 178574 112294 178642 112350
rect 178698 112294 209238 112350
rect 209294 112294 209362 112350
rect 209418 112294 239958 112350
rect 240014 112294 240082 112350
rect 240138 112294 270678 112350
rect 270734 112294 270802 112350
rect 270858 112294 281994 112350
rect 282050 112294 282118 112350
rect 282174 112294 282242 112350
rect 282298 112294 282366 112350
rect 282422 112294 312714 112350
rect 312770 112294 312838 112350
rect 312894 112294 312962 112350
rect 313018 112294 313086 112350
rect 313142 112294 324518 112350
rect 324574 112294 324642 112350
rect 324698 112294 355238 112350
rect 355294 112294 355362 112350
rect 355418 112294 385958 112350
rect 386014 112294 386082 112350
rect 386138 112294 416678 112350
rect 416734 112294 416802 112350
rect 416858 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 448518 112350
rect 448574 112294 448642 112350
rect 448698 112294 479238 112350
rect 479294 112294 479362 112350
rect 479418 112294 509958 112350
rect 510014 112294 510082 112350
rect 510138 112294 540678 112350
rect 540734 112294 540802 112350
rect 540858 112294 571398 112350
rect 571454 112294 571522 112350
rect 571578 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 22422 112226
rect 22478 112170 22546 112226
rect 22602 112170 53142 112226
rect 53198 112170 53266 112226
rect 53322 112170 83862 112226
rect 83918 112170 83986 112226
rect 84042 112170 114582 112226
rect 114638 112170 114706 112226
rect 114762 112170 145302 112226
rect 145358 112170 145426 112226
rect 145482 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 178518 112226
rect 178574 112170 178642 112226
rect 178698 112170 209238 112226
rect 209294 112170 209362 112226
rect 209418 112170 239958 112226
rect 240014 112170 240082 112226
rect 240138 112170 270678 112226
rect 270734 112170 270802 112226
rect 270858 112170 281994 112226
rect 282050 112170 282118 112226
rect 282174 112170 282242 112226
rect 282298 112170 282366 112226
rect 282422 112170 312714 112226
rect 312770 112170 312838 112226
rect 312894 112170 312962 112226
rect 313018 112170 313086 112226
rect 313142 112170 324518 112226
rect 324574 112170 324642 112226
rect 324698 112170 355238 112226
rect 355294 112170 355362 112226
rect 355418 112170 385958 112226
rect 386014 112170 386082 112226
rect 386138 112170 416678 112226
rect 416734 112170 416802 112226
rect 416858 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 448518 112226
rect 448574 112170 448642 112226
rect 448698 112170 479238 112226
rect 479294 112170 479362 112226
rect 479418 112170 509958 112226
rect 510014 112170 510082 112226
rect 510138 112170 540678 112226
rect 540734 112170 540802 112226
rect 540858 112170 571398 112226
rect 571454 112170 571522 112226
rect 571578 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 22422 112102
rect 22478 112046 22546 112102
rect 22602 112046 53142 112102
rect 53198 112046 53266 112102
rect 53322 112046 83862 112102
rect 83918 112046 83986 112102
rect 84042 112046 114582 112102
rect 114638 112046 114706 112102
rect 114762 112046 145302 112102
rect 145358 112046 145426 112102
rect 145482 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 178518 112102
rect 178574 112046 178642 112102
rect 178698 112046 209238 112102
rect 209294 112046 209362 112102
rect 209418 112046 239958 112102
rect 240014 112046 240082 112102
rect 240138 112046 270678 112102
rect 270734 112046 270802 112102
rect 270858 112046 281994 112102
rect 282050 112046 282118 112102
rect 282174 112046 282242 112102
rect 282298 112046 282366 112102
rect 282422 112046 312714 112102
rect 312770 112046 312838 112102
rect 312894 112046 312962 112102
rect 313018 112046 313086 112102
rect 313142 112046 324518 112102
rect 324574 112046 324642 112102
rect 324698 112046 355238 112102
rect 355294 112046 355362 112102
rect 355418 112046 385958 112102
rect 386014 112046 386082 112102
rect 386138 112046 416678 112102
rect 416734 112046 416802 112102
rect 416858 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 448518 112102
rect 448574 112046 448642 112102
rect 448698 112046 479238 112102
rect 479294 112046 479362 112102
rect 479418 112046 509958 112102
rect 510014 112046 510082 112102
rect 510138 112046 540678 112102
rect 540734 112046 540802 112102
rect 540858 112046 571398 112102
rect 571454 112046 571522 112102
rect 571578 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 22422 111978
rect 22478 111922 22546 111978
rect 22602 111922 53142 111978
rect 53198 111922 53266 111978
rect 53322 111922 83862 111978
rect 83918 111922 83986 111978
rect 84042 111922 114582 111978
rect 114638 111922 114706 111978
rect 114762 111922 145302 111978
rect 145358 111922 145426 111978
rect 145482 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 178518 111978
rect 178574 111922 178642 111978
rect 178698 111922 209238 111978
rect 209294 111922 209362 111978
rect 209418 111922 239958 111978
rect 240014 111922 240082 111978
rect 240138 111922 270678 111978
rect 270734 111922 270802 111978
rect 270858 111922 281994 111978
rect 282050 111922 282118 111978
rect 282174 111922 282242 111978
rect 282298 111922 282366 111978
rect 282422 111922 312714 111978
rect 312770 111922 312838 111978
rect 312894 111922 312962 111978
rect 313018 111922 313086 111978
rect 313142 111922 324518 111978
rect 324574 111922 324642 111978
rect 324698 111922 355238 111978
rect 355294 111922 355362 111978
rect 355418 111922 385958 111978
rect 386014 111922 386082 111978
rect 386138 111922 416678 111978
rect 416734 111922 416802 111978
rect 416858 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 448518 111978
rect 448574 111922 448642 111978
rect 448698 111922 479238 111978
rect 479294 111922 479362 111978
rect 479418 111922 509958 111978
rect 510014 111922 510082 111978
rect 510138 111922 540678 111978
rect 540734 111922 540802 111978
rect 540858 111922 571398 111978
rect 571454 111922 571522 111978
rect 571578 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect 271500 108298 286372 108314
rect 271500 108242 271516 108298
rect 271572 108242 286300 108298
rect 286356 108242 286372 108298
rect 271500 108226 286372 108242
rect 267916 104158 273044 104174
rect 267916 104102 267932 104158
rect 267988 104102 272972 104158
rect 273028 104102 273044 104158
rect 267916 104086 273044 104102
rect 243500 101998 424244 102014
rect 243500 101942 243516 101998
rect 243572 101942 424172 101998
rect 424228 101942 424244 101998
rect 243500 101926 424244 101942
rect 226588 101818 443284 101834
rect 226588 101762 226604 101818
rect 226660 101762 443212 101818
rect 443268 101762 443284 101818
rect 226588 101746 443284 101762
rect 226700 101638 443508 101654
rect 226700 101582 226716 101638
rect 226772 101582 443436 101638
rect 443492 101582 443508 101638
rect 226700 101566 443508 101582
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 37782 100350
rect 37838 100294 37906 100350
rect 37962 100294 68502 100350
rect 68558 100294 68626 100350
rect 68682 100294 99222 100350
rect 99278 100294 99346 100350
rect 99402 100294 129942 100350
rect 129998 100294 130066 100350
rect 130122 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 285714 100350
rect 285770 100294 285838 100350
rect 285894 100294 285962 100350
rect 286018 100294 286086 100350
rect 286142 100294 316434 100350
rect 316490 100294 316558 100350
rect 316614 100294 316682 100350
rect 316738 100294 316806 100350
rect 316862 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 463878 100350
rect 463934 100294 464002 100350
rect 464058 100294 494598 100350
rect 494654 100294 494722 100350
rect 494778 100294 525318 100350
rect 525374 100294 525442 100350
rect 525498 100294 556038 100350
rect 556094 100294 556162 100350
rect 556218 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 37782 100226
rect 37838 100170 37906 100226
rect 37962 100170 68502 100226
rect 68558 100170 68626 100226
rect 68682 100170 99222 100226
rect 99278 100170 99346 100226
rect 99402 100170 129942 100226
rect 129998 100170 130066 100226
rect 130122 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 285714 100226
rect 285770 100170 285838 100226
rect 285894 100170 285962 100226
rect 286018 100170 286086 100226
rect 286142 100170 316434 100226
rect 316490 100170 316558 100226
rect 316614 100170 316682 100226
rect 316738 100170 316806 100226
rect 316862 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 463878 100226
rect 463934 100170 464002 100226
rect 464058 100170 494598 100226
rect 494654 100170 494722 100226
rect 494778 100170 525318 100226
rect 525374 100170 525442 100226
rect 525498 100170 556038 100226
rect 556094 100170 556162 100226
rect 556218 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 37782 100102
rect 37838 100046 37906 100102
rect 37962 100046 68502 100102
rect 68558 100046 68626 100102
rect 68682 100046 99222 100102
rect 99278 100046 99346 100102
rect 99402 100046 129942 100102
rect 129998 100046 130066 100102
rect 130122 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 285714 100102
rect 285770 100046 285838 100102
rect 285894 100046 285962 100102
rect 286018 100046 286086 100102
rect 286142 100046 316434 100102
rect 316490 100046 316558 100102
rect 316614 100046 316682 100102
rect 316738 100046 316806 100102
rect 316862 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 463878 100102
rect 463934 100046 464002 100102
rect 464058 100046 494598 100102
rect 494654 100046 494722 100102
rect 494778 100046 525318 100102
rect 525374 100046 525442 100102
rect 525498 100046 556038 100102
rect 556094 100046 556162 100102
rect 556218 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 37782 99978
rect 37838 99922 37906 99978
rect 37962 99922 68502 99978
rect 68558 99922 68626 99978
rect 68682 99922 99222 99978
rect 99278 99922 99346 99978
rect 99402 99922 129942 99978
rect 129998 99922 130066 99978
rect 130122 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99923 285714 99978
rect 163262 99922 193554 99923
rect -1916 99867 193554 99922
rect 193610 99867 193678 99923
rect 193734 99867 193802 99923
rect 193858 99867 193926 99923
rect 193982 99867 224274 99923
rect 224330 99867 224398 99923
rect 224454 99867 224522 99923
rect 224578 99867 224646 99923
rect 224702 99867 254994 99923
rect 255050 99867 255118 99923
rect 255174 99867 255242 99923
rect 255298 99867 255366 99923
rect 255422 99922 285714 99923
rect 285770 99922 285838 99978
rect 285894 99922 285962 99978
rect 286018 99922 286086 99978
rect 286142 99922 316434 99978
rect 316490 99922 316558 99978
rect 316614 99922 316682 99978
rect 316738 99922 316806 99978
rect 316862 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 463878 99978
rect 463934 99922 464002 99978
rect 464058 99922 494598 99978
rect 494654 99922 494722 99978
rect 494778 99922 525318 99978
rect 525374 99922 525442 99978
rect 525498 99922 556038 99978
rect 556094 99922 556162 99978
rect 556218 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 255422 99867 597980 99922
rect -1916 99826 597980 99867
rect 235100 98578 432756 98594
rect 235100 98522 235116 98578
rect 235172 98522 432684 98578
rect 432740 98522 432756 98578
rect 235100 98506 432756 98522
rect 233420 98398 440148 98414
rect 233420 98342 233436 98398
rect 233492 98342 440076 98398
rect 440132 98342 440148 98398
rect 233420 98326 440148 98342
rect 230060 98218 443172 98234
rect 230060 98162 230076 98218
rect 230132 98162 443100 98218
rect 443156 98162 443172 98218
rect 230060 98146 443172 98162
rect 241820 96778 437796 96794
rect 241820 96722 241836 96778
rect 241892 96722 437724 96778
rect 437780 96722 437796 96778
rect 241820 96706 437796 96722
rect 228380 96598 442948 96614
rect 228380 96542 228396 96598
rect 228452 96542 442876 96598
rect 442932 96542 442948 96598
rect 228380 96526 442948 96542
rect 236780 94978 437684 94994
rect 236780 94922 236796 94978
rect 236852 94922 437612 94978
rect 437668 94922 437684 94978
rect 236780 94906 437684 94922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 22422 94350
rect 22478 94294 22546 94350
rect 22602 94294 53142 94350
rect 53198 94294 53266 94350
rect 53322 94294 83862 94350
rect 83918 94294 83986 94350
rect 84042 94294 114582 94350
rect 114638 94294 114706 94350
rect 114762 94294 145302 94350
rect 145358 94294 145426 94350
rect 145482 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 281994 94350
rect 282050 94294 282118 94350
rect 282174 94294 282242 94350
rect 282298 94294 282366 94350
rect 282422 94294 312714 94350
rect 312770 94294 312838 94350
rect 312894 94294 312962 94350
rect 313018 94294 313086 94350
rect 313142 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 448518 94350
rect 448574 94294 448642 94350
rect 448698 94294 479238 94350
rect 479294 94294 479362 94350
rect 479418 94294 509958 94350
rect 510014 94294 510082 94350
rect 510138 94294 540678 94350
rect 540734 94294 540802 94350
rect 540858 94294 571398 94350
rect 571454 94294 571522 94350
rect 571578 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 22422 94226
rect 22478 94170 22546 94226
rect 22602 94170 53142 94226
rect 53198 94170 53266 94226
rect 53322 94170 83862 94226
rect 83918 94170 83986 94226
rect 84042 94170 114582 94226
rect 114638 94170 114706 94226
rect 114762 94170 145302 94226
rect 145358 94170 145426 94226
rect 145482 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 281994 94226
rect 282050 94170 282118 94226
rect 282174 94170 282242 94226
rect 282298 94170 282366 94226
rect 282422 94170 312714 94226
rect 312770 94170 312838 94226
rect 312894 94170 312962 94226
rect 313018 94170 313086 94226
rect 313142 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 448518 94226
rect 448574 94170 448642 94226
rect 448698 94170 479238 94226
rect 479294 94170 479362 94226
rect 479418 94170 509958 94226
rect 510014 94170 510082 94226
rect 510138 94170 540678 94226
rect 540734 94170 540802 94226
rect 540858 94170 571398 94226
rect 571454 94170 571522 94226
rect 571578 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 22422 94102
rect 22478 94046 22546 94102
rect 22602 94046 53142 94102
rect 53198 94046 53266 94102
rect 53322 94046 83862 94102
rect 83918 94046 83986 94102
rect 84042 94046 114582 94102
rect 114638 94046 114706 94102
rect 114762 94046 145302 94102
rect 145358 94046 145426 94102
rect 145482 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 281994 94102
rect 282050 94046 282118 94102
rect 282174 94046 282242 94102
rect 282298 94046 282366 94102
rect 282422 94046 312714 94102
rect 312770 94046 312838 94102
rect 312894 94046 312962 94102
rect 313018 94046 313086 94102
rect 313142 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 448518 94102
rect 448574 94046 448642 94102
rect 448698 94046 479238 94102
rect 479294 94046 479362 94102
rect 479418 94046 509958 94102
rect 510014 94046 510082 94102
rect 510138 94046 540678 94102
rect 540734 94046 540802 94102
rect 540858 94046 571398 94102
rect 571454 94046 571522 94102
rect 571578 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 22422 93978
rect 22478 93922 22546 93978
rect 22602 93922 53142 93978
rect 53198 93922 53266 93978
rect 53322 93922 83862 93978
rect 83918 93922 83986 93978
rect 84042 93922 114582 93978
rect 114638 93922 114706 93978
rect 114762 93922 145302 93978
rect 145358 93922 145426 93978
rect 145482 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 281994 93978
rect 282050 93922 282118 93978
rect 282174 93922 282242 93978
rect 282298 93922 282366 93978
rect 282422 93922 312714 93978
rect 312770 93922 312838 93978
rect 312894 93922 312962 93978
rect 313018 93922 313086 93978
rect 313142 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 448518 93978
rect 448574 93922 448642 93978
rect 448698 93922 479238 93978
rect 479294 93922 479362 93978
rect 479418 93922 509958 93978
rect 510014 93922 510082 93978
rect 510138 93922 540678 93978
rect 540734 93922 540802 93978
rect 540858 93922 571398 93978
rect 571454 93922 571522 93978
rect 571578 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect 238460 93178 436340 93194
rect 238460 93122 238476 93178
rect 238532 93122 436268 93178
rect 436324 93122 436340 93178
rect 238460 93106 436340 93122
rect 229948 92458 274052 92474
rect 229948 92402 229964 92458
rect 230020 92402 273980 92458
rect 274036 92402 274052 92458
rect 229948 92386 274052 92402
rect 245180 91558 438020 91574
rect 245180 91502 245196 91558
rect 245252 91502 437948 91558
rect 438004 91502 438020 91558
rect 245180 91486 438020 91502
rect 254700 91198 433204 91214
rect 254700 91142 254716 91198
rect 254772 91142 433132 91198
rect 433188 91142 433204 91198
rect 254700 91126 433204 91142
rect 253468 91018 432532 91034
rect 253468 90962 253484 91018
rect 253540 90962 432460 91018
rect 432516 90962 432532 91018
rect 253468 90946 432532 90962
rect 251900 90838 433428 90854
rect 251900 90782 251916 90838
rect 251972 90782 433356 90838
rect 433412 90782 433428 90838
rect 251900 90766 433428 90782
rect 232076 89938 432644 89954
rect 232076 89882 232092 89938
rect 232148 89882 432572 89938
rect 432628 89882 432644 89938
rect 232076 89866 432644 89882
rect 259628 89398 431300 89414
rect 259628 89342 259644 89398
rect 259700 89342 431228 89398
rect 431284 89342 431300 89398
rect 259628 89326 431300 89342
rect 249548 89218 433092 89234
rect 249548 89162 249564 89218
rect 249620 89162 433020 89218
rect 433076 89162 433092 89218
rect 249548 89146 433092 89162
rect 206540 88498 294100 88514
rect 206540 88442 206556 88498
rect 206612 88442 294028 88498
rect 294084 88442 294100 88498
rect 206540 88426 294100 88442
rect 202508 88318 290740 88334
rect 202508 88262 202524 88318
rect 202580 88262 290668 88318
rect 290724 88262 290740 88318
rect 202508 88246 290740 88262
rect 204860 88138 292420 88154
rect 204860 88082 204876 88138
rect 204932 88082 292348 88138
rect 292404 88082 292420 88138
rect 204860 88066 292420 88082
rect 268140 87598 436564 87614
rect 268140 87542 268156 87598
rect 268212 87542 436492 87598
rect 436548 87542 436564 87598
rect 268140 87526 436564 87542
rect 246860 87418 440148 87434
rect 246860 87362 246876 87418
rect 246932 87362 440076 87418
rect 440132 87362 440148 87418
rect 246860 87346 440148 87362
rect 269932 86698 317508 86714
rect 269932 86642 269948 86698
rect 270004 86642 317436 86698
rect 317492 86642 317508 86698
rect 269932 86626 317508 86642
rect 189516 86518 282676 86534
rect 189516 86462 189532 86518
rect 189588 86462 282604 86518
rect 282660 86462 282676 86518
rect 189516 86446 282676 86462
rect 268812 85978 432980 85994
rect 268812 85922 268828 85978
rect 268884 85922 432908 85978
rect 432964 85922 432980 85978
rect 268812 85906 432980 85922
rect 266348 85798 443172 85814
rect 266348 85742 266364 85798
rect 266420 85742 443100 85798
rect 443156 85742 443172 85798
rect 266348 85726 443172 85742
rect 268028 85258 283908 85274
rect 268028 85202 268044 85258
rect 268100 85202 283836 85258
rect 283892 85202 283908 85258
rect 268028 85186 283908 85202
rect 213932 85078 296564 85094
rect 213932 85022 213948 85078
rect 214004 85022 296492 85078
rect 296548 85022 296564 85078
rect 213932 85006 296564 85022
rect 214828 84898 299140 84914
rect 214828 84842 214844 84898
rect 214900 84842 299068 84898
rect 299124 84842 299140 84898
rect 214828 84826 299140 84842
rect 317420 84358 436676 84374
rect 317420 84302 317436 84358
rect 317492 84302 436604 84358
rect 436660 84302 436676 84358
rect 317420 84286 436676 84302
rect 268252 84178 442948 84194
rect 268252 84122 268268 84178
rect 268324 84122 442876 84178
rect 442932 84122 442948 84178
rect 268252 84106 442948 84122
rect 270716 83098 317508 83114
rect 270716 83042 270732 83098
rect 270788 83042 317436 83098
rect 317492 83042 317508 83098
rect 270716 83026 317508 83042
rect 268924 82918 436340 82934
rect 268924 82862 268940 82918
rect 268996 82862 436268 82918
rect 436324 82862 436340 82918
rect 268924 82846 436340 82862
rect 254476 82738 439140 82754
rect 254476 82682 254492 82738
rect 254548 82682 439068 82738
rect 439124 82682 439140 82738
rect 254476 82666 439140 82682
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 37782 82350
rect 37838 82294 37906 82350
rect 37962 82294 68502 82350
rect 68558 82294 68626 82350
rect 68682 82294 99222 82350
rect 99278 82294 99346 82350
rect 99402 82294 129942 82350
rect 129998 82294 130066 82350
rect 130122 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 285714 82350
rect 285770 82294 285838 82350
rect 285894 82294 285962 82350
rect 286018 82294 286086 82350
rect 286142 82294 316434 82350
rect 316490 82294 316558 82350
rect 316614 82294 316682 82350
rect 316738 82294 316806 82350
rect 316862 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 463878 82350
rect 463934 82294 464002 82350
rect 464058 82294 494598 82350
rect 494654 82294 494722 82350
rect 494778 82294 525318 82350
rect 525374 82294 525442 82350
rect 525498 82294 556038 82350
rect 556094 82294 556162 82350
rect 556218 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 37782 82226
rect 37838 82170 37906 82226
rect 37962 82170 68502 82226
rect 68558 82170 68626 82226
rect 68682 82170 99222 82226
rect 99278 82170 99346 82226
rect 99402 82170 129942 82226
rect 129998 82170 130066 82226
rect 130122 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 285714 82226
rect 285770 82170 285838 82226
rect 285894 82170 285962 82226
rect 286018 82170 286086 82226
rect 286142 82170 316434 82226
rect 316490 82170 316558 82226
rect 316614 82170 316682 82226
rect 316738 82170 316806 82226
rect 316862 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 463878 82226
rect 463934 82170 464002 82226
rect 464058 82170 494598 82226
rect 494654 82170 494722 82226
rect 494778 82170 525318 82226
rect 525374 82170 525442 82226
rect 525498 82170 556038 82226
rect 556094 82170 556162 82226
rect 556218 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 37782 82102
rect 37838 82046 37906 82102
rect 37962 82046 68502 82102
rect 68558 82046 68626 82102
rect 68682 82046 99222 82102
rect 99278 82046 99346 82102
rect 99402 82046 129942 82102
rect 129998 82046 130066 82102
rect 130122 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 285714 82102
rect 285770 82046 285838 82102
rect 285894 82046 285962 82102
rect 286018 82046 286086 82102
rect 286142 82046 316434 82102
rect 316490 82046 316558 82102
rect 316614 82046 316682 82102
rect 316738 82046 316806 82102
rect 316862 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 463878 82102
rect 463934 82046 464002 82102
rect 464058 82046 494598 82102
rect 494654 82046 494722 82102
rect 494778 82046 525318 82102
rect 525374 82046 525442 82102
rect 525498 82046 556038 82102
rect 556094 82046 556162 82102
rect 556218 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 37782 81978
rect 37838 81922 37906 81978
rect 37962 81922 68502 81978
rect 68558 81922 68626 81978
rect 68682 81922 99222 81978
rect 99278 81922 99346 81978
rect 99402 81922 129942 81978
rect 129998 81922 130066 81978
rect 130122 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 285714 81978
rect 285770 81922 285838 81978
rect 285894 81922 285962 81978
rect 286018 81922 286086 81978
rect 286142 81922 316434 81978
rect 316490 81922 316558 81978
rect 316614 81922 316682 81978
rect 316738 81922 316806 81978
rect 316862 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 463878 81978
rect 463934 81922 464002 81978
rect 464058 81922 494598 81978
rect 494654 81922 494722 81978
rect 494778 81922 525318 81978
rect 525374 81922 525442 81978
rect 525498 81922 556038 81978
rect 556094 81922 556162 81978
rect 556218 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect 181452 81478 273940 81494
rect 181452 81422 181468 81478
rect 181524 81422 273868 81478
rect 273924 81422 273940 81478
rect 181452 81406 273940 81422
rect 252908 80938 438916 80954
rect 252908 80882 252924 80938
rect 252980 80882 438844 80938
rect 438900 80882 438916 80938
rect 252908 80866 438916 80882
rect 256940 80758 443284 80774
rect 256940 80702 256956 80758
rect 257012 80702 443212 80758
rect 443268 80702 443284 80758
rect 256940 80686 443284 80702
rect 234764 80578 442724 80594
rect 234764 80522 234780 80578
rect 234836 80522 442652 80578
rect 442708 80522 442724 80578
rect 234764 80506 442724 80522
rect 229948 80398 434548 80414
rect 229948 80342 229964 80398
rect 230020 80342 434476 80398
rect 434532 80342 434548 80398
rect 229948 80326 434548 80342
rect 231404 80218 434324 80234
rect 231404 80162 231420 80218
rect 231476 80162 434252 80218
rect 434308 80162 434324 80218
rect 231404 80146 434324 80162
rect 232748 80038 427604 80054
rect 232748 79982 232764 80038
rect 232820 79982 427532 80038
rect 427588 79982 427604 80038
rect 232748 79966 427604 79982
rect 230732 79858 425924 79874
rect 230732 79802 230748 79858
rect 230804 79802 425852 79858
rect 425908 79802 425924 79858
rect 230732 79786 425924 79802
rect 227260 78958 315044 78974
rect 227260 78902 227276 78958
rect 227332 78902 314972 78958
rect 315028 78902 315044 78958
rect 227260 78886 315044 78902
rect 250892 78058 438692 78074
rect 250892 78002 250908 78058
rect 250964 78002 438620 78058
rect 438676 78002 438692 78058
rect 250892 77986 438692 78002
rect 268700 77698 436788 77714
rect 268700 77642 268716 77698
rect 268772 77642 436716 77698
rect 436772 77642 436788 77698
rect 268700 77626 436788 77642
rect 267916 77338 440036 77354
rect 267916 77282 267932 77338
rect 267988 77282 439964 77338
rect 440020 77282 440036 77338
rect 267916 77266 440036 77282
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 22422 76350
rect 22478 76294 22546 76350
rect 22602 76294 53142 76350
rect 53198 76294 53266 76350
rect 53322 76294 83862 76350
rect 83918 76294 83986 76350
rect 84042 76294 114582 76350
rect 114638 76294 114706 76350
rect 114762 76294 145302 76350
rect 145358 76294 145426 76350
rect 145482 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 271702 76350
rect 271758 76294 271826 76350
rect 271882 76294 302422 76350
rect 302478 76294 302546 76350
rect 302602 76294 333142 76350
rect 333198 76294 333266 76350
rect 333322 76294 363862 76350
rect 363918 76294 363986 76350
rect 364042 76294 394582 76350
rect 394638 76294 394706 76350
rect 394762 76294 425302 76350
rect 425358 76294 425426 76350
rect 425482 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 448518 76350
rect 448574 76294 448642 76350
rect 448698 76294 479238 76350
rect 479294 76294 479362 76350
rect 479418 76294 509958 76350
rect 510014 76294 510082 76350
rect 510138 76294 540678 76350
rect 540734 76294 540802 76350
rect 540858 76294 571398 76350
rect 571454 76294 571522 76350
rect 571578 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 22422 76226
rect 22478 76170 22546 76226
rect 22602 76170 53142 76226
rect 53198 76170 53266 76226
rect 53322 76170 83862 76226
rect 83918 76170 83986 76226
rect 84042 76170 114582 76226
rect 114638 76170 114706 76226
rect 114762 76170 145302 76226
rect 145358 76170 145426 76226
rect 145482 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 271702 76226
rect 271758 76170 271826 76226
rect 271882 76170 302422 76226
rect 302478 76170 302546 76226
rect 302602 76170 333142 76226
rect 333198 76170 333266 76226
rect 333322 76170 363862 76226
rect 363918 76170 363986 76226
rect 364042 76170 394582 76226
rect 394638 76170 394706 76226
rect 394762 76170 425302 76226
rect 425358 76170 425426 76226
rect 425482 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 448518 76226
rect 448574 76170 448642 76226
rect 448698 76170 479238 76226
rect 479294 76170 479362 76226
rect 479418 76170 509958 76226
rect 510014 76170 510082 76226
rect 510138 76170 540678 76226
rect 540734 76170 540802 76226
rect 540858 76170 571398 76226
rect 571454 76170 571522 76226
rect 571578 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 22422 76102
rect 22478 76046 22546 76102
rect 22602 76046 53142 76102
rect 53198 76046 53266 76102
rect 53322 76046 83862 76102
rect 83918 76046 83986 76102
rect 84042 76046 114582 76102
rect 114638 76046 114706 76102
rect 114762 76046 145302 76102
rect 145358 76046 145426 76102
rect 145482 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 271702 76102
rect 271758 76046 271826 76102
rect 271882 76046 302422 76102
rect 302478 76046 302546 76102
rect 302602 76046 333142 76102
rect 333198 76046 333266 76102
rect 333322 76046 363862 76102
rect 363918 76046 363986 76102
rect 364042 76046 394582 76102
rect 394638 76046 394706 76102
rect 394762 76046 425302 76102
rect 425358 76046 425426 76102
rect 425482 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 448518 76102
rect 448574 76046 448642 76102
rect 448698 76046 479238 76102
rect 479294 76046 479362 76102
rect 479418 76046 509958 76102
rect 510014 76046 510082 76102
rect 510138 76046 540678 76102
rect 540734 76046 540802 76102
rect 540858 76046 571398 76102
rect 571454 76046 571522 76102
rect 571578 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 22422 75978
rect 22478 75922 22546 75978
rect 22602 75922 53142 75978
rect 53198 75922 53266 75978
rect 53322 75922 83862 75978
rect 83918 75922 83986 75978
rect 84042 75922 114582 75978
rect 114638 75922 114706 75978
rect 114762 75922 145302 75978
rect 145358 75922 145426 75978
rect 145482 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 271702 75978
rect 271758 75922 271826 75978
rect 271882 75922 302422 75978
rect 302478 75922 302546 75978
rect 302602 75922 333142 75978
rect 333198 75922 333266 75978
rect 333322 75922 363862 75978
rect 363918 75922 363986 75978
rect 364042 75922 394582 75978
rect 394638 75922 394706 75978
rect 394762 75922 425302 75978
rect 425358 75922 425426 75978
rect 425482 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 448518 75978
rect 448574 75922 448642 75978
rect 448698 75922 479238 75978
rect 479294 75922 479362 75978
rect 479418 75922 509958 75978
rect 510014 75922 510082 75978
rect 510138 75922 540678 75978
rect 540734 75922 540802 75978
rect 540858 75922 571398 75978
rect 571454 75922 571522 75978
rect 571578 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect 428076 75538 428724 75554
rect 428076 75482 428092 75538
rect 428148 75482 428652 75538
rect 428708 75482 428724 75538
rect 428076 75466 428724 75482
rect 268588 74098 274164 74114
rect 268588 74042 268604 74098
rect 268660 74042 274092 74098
rect 274148 74042 274164 74098
rect 268588 74026 274164 74042
rect 268476 73198 273380 73214
rect 268476 73142 268492 73198
rect 268548 73142 273308 73198
rect 273364 73142 273380 73198
rect 268476 73126 273380 73142
rect 266908 73018 273604 73034
rect 266908 72962 266924 73018
rect 266980 72962 273532 73018
rect 273588 72962 273604 73018
rect 266908 72946 273604 72962
rect 266796 69778 273716 69794
rect 266796 69722 266812 69778
rect 266868 69722 273644 69778
rect 273700 69722 273716 69778
rect 266796 69706 273716 69722
rect 420796 67978 442724 67994
rect 420796 67922 420812 67978
rect 420868 67922 442652 67978
rect 442708 67922 442724 67978
rect 420796 67906 442724 67922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 37782 64350
rect 37838 64294 37906 64350
rect 37962 64294 68502 64350
rect 68558 64294 68626 64350
rect 68682 64294 99222 64350
rect 99278 64294 99346 64350
rect 99402 64294 129942 64350
rect 129998 64294 130066 64350
rect 130122 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 185878 64350
rect 185934 64294 186002 64350
rect 186058 64294 216598 64350
rect 216654 64294 216722 64350
rect 216778 64294 247318 64350
rect 247374 64294 247442 64350
rect 247498 64294 287062 64350
rect 287118 64294 287186 64350
rect 287242 64294 317782 64350
rect 317838 64294 317906 64350
rect 317962 64294 348502 64350
rect 348558 64294 348626 64350
rect 348682 64294 379222 64350
rect 379278 64294 379346 64350
rect 379402 64294 409942 64350
rect 409998 64294 410066 64350
rect 410122 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 463878 64350
rect 463934 64294 464002 64350
rect 464058 64294 494598 64350
rect 494654 64294 494722 64350
rect 494778 64294 525318 64350
rect 525374 64294 525442 64350
rect 525498 64294 556038 64350
rect 556094 64294 556162 64350
rect 556218 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 37782 64226
rect 37838 64170 37906 64226
rect 37962 64170 68502 64226
rect 68558 64170 68626 64226
rect 68682 64170 99222 64226
rect 99278 64170 99346 64226
rect 99402 64170 129942 64226
rect 129998 64170 130066 64226
rect 130122 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 185878 64226
rect 185934 64170 186002 64226
rect 186058 64170 216598 64226
rect 216654 64170 216722 64226
rect 216778 64170 247318 64226
rect 247374 64170 247442 64226
rect 247498 64170 287062 64226
rect 287118 64170 287186 64226
rect 287242 64170 317782 64226
rect 317838 64170 317906 64226
rect 317962 64170 348502 64226
rect 348558 64170 348626 64226
rect 348682 64170 379222 64226
rect 379278 64170 379346 64226
rect 379402 64170 409942 64226
rect 409998 64170 410066 64226
rect 410122 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 463878 64226
rect 463934 64170 464002 64226
rect 464058 64170 494598 64226
rect 494654 64170 494722 64226
rect 494778 64170 525318 64226
rect 525374 64170 525442 64226
rect 525498 64170 556038 64226
rect 556094 64170 556162 64226
rect 556218 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 37782 64102
rect 37838 64046 37906 64102
rect 37962 64046 68502 64102
rect 68558 64046 68626 64102
rect 68682 64046 99222 64102
rect 99278 64046 99346 64102
rect 99402 64046 129942 64102
rect 129998 64046 130066 64102
rect 130122 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 185878 64102
rect 185934 64046 186002 64102
rect 186058 64046 216598 64102
rect 216654 64046 216722 64102
rect 216778 64046 247318 64102
rect 247374 64046 247442 64102
rect 247498 64046 287062 64102
rect 287118 64046 287186 64102
rect 287242 64046 317782 64102
rect 317838 64046 317906 64102
rect 317962 64046 348502 64102
rect 348558 64046 348626 64102
rect 348682 64046 379222 64102
rect 379278 64046 379346 64102
rect 379402 64046 409942 64102
rect 409998 64046 410066 64102
rect 410122 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 463878 64102
rect 463934 64046 464002 64102
rect 464058 64046 494598 64102
rect 494654 64046 494722 64102
rect 494778 64046 525318 64102
rect 525374 64046 525442 64102
rect 525498 64046 556038 64102
rect 556094 64046 556162 64102
rect 556218 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 37782 63978
rect 37838 63922 37906 63978
rect 37962 63922 68502 63978
rect 68558 63922 68626 63978
rect 68682 63922 99222 63978
rect 99278 63922 99346 63978
rect 99402 63922 129942 63978
rect 129998 63922 130066 63978
rect 130122 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 185878 63978
rect 185934 63922 186002 63978
rect 186058 63922 216598 63978
rect 216654 63922 216722 63978
rect 216778 63922 247318 63978
rect 247374 63922 247442 63978
rect 247498 63922 287062 63978
rect 287118 63922 287186 63978
rect 287242 63922 317782 63978
rect 317838 63922 317906 63978
rect 317962 63922 348502 63978
rect 348558 63922 348626 63978
rect 348682 63922 379222 63978
rect 379278 63922 379346 63978
rect 379402 63922 409942 63978
rect 409998 63922 410066 63978
rect 410122 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 463878 63978
rect 463934 63922 464002 63978
rect 464058 63922 494598 63978
rect 494654 63922 494722 63978
rect 494778 63922 525318 63978
rect 525374 63922 525442 63978
rect 525498 63922 556038 63978
rect 556094 63922 556162 63978
rect 556218 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 22422 58350
rect 22478 58294 22546 58350
rect 22602 58294 53142 58350
rect 53198 58294 53266 58350
rect 53322 58294 83862 58350
rect 83918 58294 83986 58350
rect 84042 58294 114582 58350
rect 114638 58294 114706 58350
rect 114762 58294 145302 58350
rect 145358 58294 145426 58350
rect 145482 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 170518 58350
rect 170574 58294 170642 58350
rect 170698 58294 201238 58350
rect 201294 58294 201362 58350
rect 201418 58294 231958 58350
rect 232014 58294 232082 58350
rect 232138 58294 262678 58350
rect 262734 58294 262802 58350
rect 262858 58294 271702 58350
rect 271758 58294 271826 58350
rect 271882 58294 302422 58350
rect 302478 58294 302546 58350
rect 302602 58294 333142 58350
rect 333198 58294 333266 58350
rect 333322 58294 363862 58350
rect 363918 58294 363986 58350
rect 364042 58294 394582 58350
rect 394638 58294 394706 58350
rect 394762 58294 425302 58350
rect 425358 58294 425426 58350
rect 425482 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 448518 58350
rect 448574 58294 448642 58350
rect 448698 58294 479238 58350
rect 479294 58294 479362 58350
rect 479418 58294 509958 58350
rect 510014 58294 510082 58350
rect 510138 58294 540678 58350
rect 540734 58294 540802 58350
rect 540858 58294 571398 58350
rect 571454 58294 571522 58350
rect 571578 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 22422 58226
rect 22478 58170 22546 58226
rect 22602 58170 53142 58226
rect 53198 58170 53266 58226
rect 53322 58170 83862 58226
rect 83918 58170 83986 58226
rect 84042 58170 114582 58226
rect 114638 58170 114706 58226
rect 114762 58170 145302 58226
rect 145358 58170 145426 58226
rect 145482 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 170518 58226
rect 170574 58170 170642 58226
rect 170698 58170 201238 58226
rect 201294 58170 201362 58226
rect 201418 58170 231958 58226
rect 232014 58170 232082 58226
rect 232138 58170 262678 58226
rect 262734 58170 262802 58226
rect 262858 58170 271702 58226
rect 271758 58170 271826 58226
rect 271882 58170 302422 58226
rect 302478 58170 302546 58226
rect 302602 58170 333142 58226
rect 333198 58170 333266 58226
rect 333322 58170 363862 58226
rect 363918 58170 363986 58226
rect 364042 58170 394582 58226
rect 394638 58170 394706 58226
rect 394762 58170 425302 58226
rect 425358 58170 425426 58226
rect 425482 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 448518 58226
rect 448574 58170 448642 58226
rect 448698 58170 479238 58226
rect 479294 58170 479362 58226
rect 479418 58170 509958 58226
rect 510014 58170 510082 58226
rect 510138 58170 540678 58226
rect 540734 58170 540802 58226
rect 540858 58170 571398 58226
rect 571454 58170 571522 58226
rect 571578 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 22422 58102
rect 22478 58046 22546 58102
rect 22602 58046 53142 58102
rect 53198 58046 53266 58102
rect 53322 58046 83862 58102
rect 83918 58046 83986 58102
rect 84042 58046 114582 58102
rect 114638 58046 114706 58102
rect 114762 58046 145302 58102
rect 145358 58046 145426 58102
rect 145482 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 170518 58102
rect 170574 58046 170642 58102
rect 170698 58046 201238 58102
rect 201294 58046 201362 58102
rect 201418 58046 231958 58102
rect 232014 58046 232082 58102
rect 232138 58046 262678 58102
rect 262734 58046 262802 58102
rect 262858 58046 271702 58102
rect 271758 58046 271826 58102
rect 271882 58046 302422 58102
rect 302478 58046 302546 58102
rect 302602 58046 333142 58102
rect 333198 58046 333266 58102
rect 333322 58046 363862 58102
rect 363918 58046 363986 58102
rect 364042 58046 394582 58102
rect 394638 58046 394706 58102
rect 394762 58046 425302 58102
rect 425358 58046 425426 58102
rect 425482 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 448518 58102
rect 448574 58046 448642 58102
rect 448698 58046 479238 58102
rect 479294 58046 479362 58102
rect 479418 58046 509958 58102
rect 510014 58046 510082 58102
rect 510138 58046 540678 58102
rect 540734 58046 540802 58102
rect 540858 58046 571398 58102
rect 571454 58046 571522 58102
rect 571578 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 22422 57978
rect 22478 57922 22546 57978
rect 22602 57922 53142 57978
rect 53198 57922 53266 57978
rect 53322 57922 83862 57978
rect 83918 57922 83986 57978
rect 84042 57922 114582 57978
rect 114638 57922 114706 57978
rect 114762 57922 145302 57978
rect 145358 57922 145426 57978
rect 145482 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 170518 57978
rect 170574 57922 170642 57978
rect 170698 57922 201238 57978
rect 201294 57922 201362 57978
rect 201418 57922 231958 57978
rect 232014 57922 232082 57978
rect 232138 57922 262678 57978
rect 262734 57922 262802 57978
rect 262858 57922 271702 57978
rect 271758 57922 271826 57978
rect 271882 57922 302422 57978
rect 302478 57922 302546 57978
rect 302602 57922 333142 57978
rect 333198 57922 333266 57978
rect 333322 57922 363862 57978
rect 363918 57922 363986 57978
rect 364042 57922 394582 57978
rect 394638 57922 394706 57978
rect 394762 57922 425302 57978
rect 425358 57922 425426 57978
rect 425482 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 448518 57978
rect 448574 57922 448642 57978
rect 448698 57922 479238 57978
rect 479294 57922 479362 57978
rect 479418 57922 509958 57978
rect 510014 57922 510082 57978
rect 510138 57922 540678 57978
rect 540734 57922 540802 57978
rect 540858 57922 571398 57978
rect 571454 57922 571522 57978
rect 571578 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 264556 54658 273156 54674
rect 264556 54602 264572 54658
rect 264628 54602 273084 54658
rect 273140 54602 273156 54658
rect 264556 54586 273156 54602
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 37782 46350
rect 37838 46294 37906 46350
rect 37962 46294 68502 46350
rect 68558 46294 68626 46350
rect 68682 46294 99222 46350
rect 99278 46294 99346 46350
rect 99402 46294 129942 46350
rect 129998 46294 130066 46350
rect 130122 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 185878 46350
rect 185934 46294 186002 46350
rect 186058 46294 216598 46350
rect 216654 46294 216722 46350
rect 216778 46294 247318 46350
rect 247374 46294 247442 46350
rect 247498 46294 287062 46350
rect 287118 46294 287186 46350
rect 287242 46294 317782 46350
rect 317838 46294 317906 46350
rect 317962 46294 348502 46350
rect 348558 46294 348626 46350
rect 348682 46294 379222 46350
rect 379278 46294 379346 46350
rect 379402 46294 409942 46350
rect 409998 46294 410066 46350
rect 410122 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 463878 46350
rect 463934 46294 464002 46350
rect 464058 46294 494598 46350
rect 494654 46294 494722 46350
rect 494778 46294 525318 46350
rect 525374 46294 525442 46350
rect 525498 46294 556038 46350
rect 556094 46294 556162 46350
rect 556218 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 37782 46226
rect 37838 46170 37906 46226
rect 37962 46170 68502 46226
rect 68558 46170 68626 46226
rect 68682 46170 99222 46226
rect 99278 46170 99346 46226
rect 99402 46170 129942 46226
rect 129998 46170 130066 46226
rect 130122 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 185878 46226
rect 185934 46170 186002 46226
rect 186058 46170 216598 46226
rect 216654 46170 216722 46226
rect 216778 46170 247318 46226
rect 247374 46170 247442 46226
rect 247498 46170 287062 46226
rect 287118 46170 287186 46226
rect 287242 46170 317782 46226
rect 317838 46170 317906 46226
rect 317962 46170 348502 46226
rect 348558 46170 348626 46226
rect 348682 46170 379222 46226
rect 379278 46170 379346 46226
rect 379402 46170 409942 46226
rect 409998 46170 410066 46226
rect 410122 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 463878 46226
rect 463934 46170 464002 46226
rect 464058 46170 494598 46226
rect 494654 46170 494722 46226
rect 494778 46170 525318 46226
rect 525374 46170 525442 46226
rect 525498 46170 556038 46226
rect 556094 46170 556162 46226
rect 556218 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 37782 46102
rect 37838 46046 37906 46102
rect 37962 46046 68502 46102
rect 68558 46046 68626 46102
rect 68682 46046 99222 46102
rect 99278 46046 99346 46102
rect 99402 46046 129942 46102
rect 129998 46046 130066 46102
rect 130122 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 185878 46102
rect 185934 46046 186002 46102
rect 186058 46046 216598 46102
rect 216654 46046 216722 46102
rect 216778 46046 247318 46102
rect 247374 46046 247442 46102
rect 247498 46046 287062 46102
rect 287118 46046 287186 46102
rect 287242 46046 317782 46102
rect 317838 46046 317906 46102
rect 317962 46046 348502 46102
rect 348558 46046 348626 46102
rect 348682 46046 379222 46102
rect 379278 46046 379346 46102
rect 379402 46046 409942 46102
rect 409998 46046 410066 46102
rect 410122 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 463878 46102
rect 463934 46046 464002 46102
rect 464058 46046 494598 46102
rect 494654 46046 494722 46102
rect 494778 46046 525318 46102
rect 525374 46046 525442 46102
rect 525498 46046 556038 46102
rect 556094 46046 556162 46102
rect 556218 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 37782 45978
rect 37838 45922 37906 45978
rect 37962 45922 68502 45978
rect 68558 45922 68626 45978
rect 68682 45922 99222 45978
rect 99278 45922 99346 45978
rect 99402 45922 129942 45978
rect 129998 45922 130066 45978
rect 130122 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 185878 45978
rect 185934 45922 186002 45978
rect 186058 45922 216598 45978
rect 216654 45922 216722 45978
rect 216778 45922 247318 45978
rect 247374 45922 247442 45978
rect 247498 45922 287062 45978
rect 287118 45922 287186 45978
rect 287242 45922 317782 45978
rect 317838 45922 317906 45978
rect 317962 45922 348502 45978
rect 348558 45922 348626 45978
rect 348682 45922 379222 45978
rect 379278 45922 379346 45978
rect 379402 45922 409942 45978
rect 409998 45922 410066 45978
rect 410122 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 463878 45978
rect 463934 45922 464002 45978
rect 464058 45922 494598 45978
rect 494654 45922 494722 45978
rect 494778 45922 525318 45978
rect 525374 45922 525442 45978
rect 525498 45922 556038 45978
rect 556094 45922 556162 45978
rect 556218 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 22422 40350
rect 22478 40294 22546 40350
rect 22602 40294 53142 40350
rect 53198 40294 53266 40350
rect 53322 40294 83862 40350
rect 83918 40294 83986 40350
rect 84042 40294 114582 40350
rect 114638 40294 114706 40350
rect 114762 40294 145302 40350
rect 145358 40294 145426 40350
rect 145482 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 170518 40350
rect 170574 40294 170642 40350
rect 170698 40294 201238 40350
rect 201294 40294 201362 40350
rect 201418 40294 231958 40350
rect 232014 40294 232082 40350
rect 232138 40294 262678 40350
rect 262734 40294 262802 40350
rect 262858 40294 271702 40350
rect 271758 40294 271826 40350
rect 271882 40294 302422 40350
rect 302478 40294 302546 40350
rect 302602 40294 333142 40350
rect 333198 40294 333266 40350
rect 333322 40294 363862 40350
rect 363918 40294 363986 40350
rect 364042 40294 394582 40350
rect 394638 40294 394706 40350
rect 394762 40294 425302 40350
rect 425358 40294 425426 40350
rect 425482 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 448518 40350
rect 448574 40294 448642 40350
rect 448698 40294 479238 40350
rect 479294 40294 479362 40350
rect 479418 40294 509958 40350
rect 510014 40294 510082 40350
rect 510138 40294 540678 40350
rect 540734 40294 540802 40350
rect 540858 40294 571398 40350
rect 571454 40294 571522 40350
rect 571578 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 22422 40226
rect 22478 40170 22546 40226
rect 22602 40170 53142 40226
rect 53198 40170 53266 40226
rect 53322 40170 83862 40226
rect 83918 40170 83986 40226
rect 84042 40170 114582 40226
rect 114638 40170 114706 40226
rect 114762 40170 145302 40226
rect 145358 40170 145426 40226
rect 145482 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 170518 40226
rect 170574 40170 170642 40226
rect 170698 40170 201238 40226
rect 201294 40170 201362 40226
rect 201418 40170 231958 40226
rect 232014 40170 232082 40226
rect 232138 40170 262678 40226
rect 262734 40170 262802 40226
rect 262858 40170 271702 40226
rect 271758 40170 271826 40226
rect 271882 40170 302422 40226
rect 302478 40170 302546 40226
rect 302602 40170 333142 40226
rect 333198 40170 333266 40226
rect 333322 40170 363862 40226
rect 363918 40170 363986 40226
rect 364042 40170 394582 40226
rect 394638 40170 394706 40226
rect 394762 40170 425302 40226
rect 425358 40170 425426 40226
rect 425482 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 448518 40226
rect 448574 40170 448642 40226
rect 448698 40170 479238 40226
rect 479294 40170 479362 40226
rect 479418 40170 509958 40226
rect 510014 40170 510082 40226
rect 510138 40170 540678 40226
rect 540734 40170 540802 40226
rect 540858 40170 571398 40226
rect 571454 40170 571522 40226
rect 571578 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 22422 40102
rect 22478 40046 22546 40102
rect 22602 40046 53142 40102
rect 53198 40046 53266 40102
rect 53322 40046 83862 40102
rect 83918 40046 83986 40102
rect 84042 40046 114582 40102
rect 114638 40046 114706 40102
rect 114762 40046 145302 40102
rect 145358 40046 145426 40102
rect 145482 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 170518 40102
rect 170574 40046 170642 40102
rect 170698 40046 201238 40102
rect 201294 40046 201362 40102
rect 201418 40046 231958 40102
rect 232014 40046 232082 40102
rect 232138 40046 262678 40102
rect 262734 40046 262802 40102
rect 262858 40046 271702 40102
rect 271758 40046 271826 40102
rect 271882 40046 302422 40102
rect 302478 40046 302546 40102
rect 302602 40046 333142 40102
rect 333198 40046 333266 40102
rect 333322 40046 363862 40102
rect 363918 40046 363986 40102
rect 364042 40046 394582 40102
rect 394638 40046 394706 40102
rect 394762 40046 425302 40102
rect 425358 40046 425426 40102
rect 425482 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 448518 40102
rect 448574 40046 448642 40102
rect 448698 40046 479238 40102
rect 479294 40046 479362 40102
rect 479418 40046 509958 40102
rect 510014 40046 510082 40102
rect 510138 40046 540678 40102
rect 540734 40046 540802 40102
rect 540858 40046 571398 40102
rect 571454 40046 571522 40102
rect 571578 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 22422 39978
rect 22478 39922 22546 39978
rect 22602 39922 53142 39978
rect 53198 39922 53266 39978
rect 53322 39922 83862 39978
rect 83918 39922 83986 39978
rect 84042 39922 114582 39978
rect 114638 39922 114706 39978
rect 114762 39922 145302 39978
rect 145358 39922 145426 39978
rect 145482 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 170518 39978
rect 170574 39922 170642 39978
rect 170698 39922 201238 39978
rect 201294 39922 201362 39978
rect 201418 39922 231958 39978
rect 232014 39922 232082 39978
rect 232138 39922 262678 39978
rect 262734 39922 262802 39978
rect 262858 39922 271702 39978
rect 271758 39922 271826 39978
rect 271882 39922 302422 39978
rect 302478 39922 302546 39978
rect 302602 39922 333142 39978
rect 333198 39922 333266 39978
rect 333322 39922 363862 39978
rect 363918 39922 363986 39978
rect 364042 39922 394582 39978
rect 394638 39922 394706 39978
rect 394762 39922 425302 39978
rect 425358 39922 425426 39978
rect 425482 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 448518 39978
rect 448574 39922 448642 39978
rect 448698 39922 479238 39978
rect 479294 39922 479362 39978
rect 479418 39922 509958 39978
rect 510014 39922 510082 39978
rect 510138 39922 540678 39978
rect 540734 39922 540802 39978
rect 540858 39922 571398 39978
rect 571454 39922 571522 39978
rect 571578 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 37782 28350
rect 37838 28294 37906 28350
rect 37962 28294 68502 28350
rect 68558 28294 68626 28350
rect 68682 28294 99222 28350
rect 99278 28294 99346 28350
rect 99402 28294 129942 28350
rect 129998 28294 130066 28350
rect 130122 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 185878 28350
rect 185934 28294 186002 28350
rect 186058 28294 216598 28350
rect 216654 28294 216722 28350
rect 216778 28294 247318 28350
rect 247374 28294 247442 28350
rect 247498 28294 287062 28350
rect 287118 28294 287186 28350
rect 287242 28294 317782 28350
rect 317838 28294 317906 28350
rect 317962 28294 348502 28350
rect 348558 28294 348626 28350
rect 348682 28294 379222 28350
rect 379278 28294 379346 28350
rect 379402 28294 409942 28350
rect 409998 28294 410066 28350
rect 410122 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 463878 28350
rect 463934 28294 464002 28350
rect 464058 28294 494598 28350
rect 494654 28294 494722 28350
rect 494778 28294 525318 28350
rect 525374 28294 525442 28350
rect 525498 28294 556038 28350
rect 556094 28294 556162 28350
rect 556218 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 37782 28226
rect 37838 28170 37906 28226
rect 37962 28170 68502 28226
rect 68558 28170 68626 28226
rect 68682 28170 99222 28226
rect 99278 28170 99346 28226
rect 99402 28170 129942 28226
rect 129998 28170 130066 28226
rect 130122 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 185878 28226
rect 185934 28170 186002 28226
rect 186058 28170 216598 28226
rect 216654 28170 216722 28226
rect 216778 28170 247318 28226
rect 247374 28170 247442 28226
rect 247498 28170 287062 28226
rect 287118 28170 287186 28226
rect 287242 28170 317782 28226
rect 317838 28170 317906 28226
rect 317962 28170 348502 28226
rect 348558 28170 348626 28226
rect 348682 28170 379222 28226
rect 379278 28170 379346 28226
rect 379402 28170 409942 28226
rect 409998 28170 410066 28226
rect 410122 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 463878 28226
rect 463934 28170 464002 28226
rect 464058 28170 494598 28226
rect 494654 28170 494722 28226
rect 494778 28170 525318 28226
rect 525374 28170 525442 28226
rect 525498 28170 556038 28226
rect 556094 28170 556162 28226
rect 556218 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 37782 28102
rect 37838 28046 37906 28102
rect 37962 28046 68502 28102
rect 68558 28046 68626 28102
rect 68682 28046 99222 28102
rect 99278 28046 99346 28102
rect 99402 28046 129942 28102
rect 129998 28046 130066 28102
rect 130122 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 185878 28102
rect 185934 28046 186002 28102
rect 186058 28046 216598 28102
rect 216654 28046 216722 28102
rect 216778 28046 247318 28102
rect 247374 28046 247442 28102
rect 247498 28046 287062 28102
rect 287118 28046 287186 28102
rect 287242 28046 317782 28102
rect 317838 28046 317906 28102
rect 317962 28046 348502 28102
rect 348558 28046 348626 28102
rect 348682 28046 379222 28102
rect 379278 28046 379346 28102
rect 379402 28046 409942 28102
rect 409998 28046 410066 28102
rect 410122 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 463878 28102
rect 463934 28046 464002 28102
rect 464058 28046 494598 28102
rect 494654 28046 494722 28102
rect 494778 28046 525318 28102
rect 525374 28046 525442 28102
rect 525498 28046 556038 28102
rect 556094 28046 556162 28102
rect 556218 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 37782 27978
rect 37838 27922 37906 27978
rect 37962 27922 68502 27978
rect 68558 27922 68626 27978
rect 68682 27922 99222 27978
rect 99278 27922 99346 27978
rect 99402 27922 129942 27978
rect 129998 27922 130066 27978
rect 130122 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 185878 27978
rect 185934 27922 186002 27978
rect 186058 27922 216598 27978
rect 216654 27922 216722 27978
rect 216778 27922 247318 27978
rect 247374 27922 247442 27978
rect 247498 27922 287062 27978
rect 287118 27922 287186 27978
rect 287242 27922 317782 27978
rect 317838 27922 317906 27978
rect 317962 27922 348502 27978
rect 348558 27922 348626 27978
rect 348682 27922 379222 27978
rect 379278 27922 379346 27978
rect 379402 27922 409942 27978
rect 409998 27922 410066 27978
rect 410122 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 463878 27978
rect 463934 27922 464002 27978
rect 464058 27922 494598 27978
rect 494654 27922 494722 27978
rect 494778 27922 525318 27978
rect 525374 27922 525442 27978
rect 525498 27922 556038 27978
rect 556094 27922 556162 27978
rect 556218 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 170518 22350
rect 170574 22294 170642 22350
rect 170698 22294 201238 22350
rect 201294 22294 201362 22350
rect 201418 22294 231958 22350
rect 232014 22294 232082 22350
rect 232138 22294 262678 22350
rect 262734 22294 262802 22350
rect 262858 22294 271702 22350
rect 271758 22294 271826 22350
rect 271882 22294 302422 22350
rect 302478 22294 302546 22350
rect 302602 22294 333142 22350
rect 333198 22294 333266 22350
rect 333322 22294 363862 22350
rect 363918 22294 363986 22350
rect 364042 22294 394582 22350
rect 394638 22294 394706 22350
rect 394762 22294 425302 22350
rect 425358 22294 425426 22350
rect 425482 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 170518 22226
rect 170574 22170 170642 22226
rect 170698 22170 201238 22226
rect 201294 22170 201362 22226
rect 201418 22170 231958 22226
rect 232014 22170 232082 22226
rect 232138 22170 262678 22226
rect 262734 22170 262802 22226
rect 262858 22170 271702 22226
rect 271758 22170 271826 22226
rect 271882 22170 302422 22226
rect 302478 22170 302546 22226
rect 302602 22170 333142 22226
rect 333198 22170 333266 22226
rect 333322 22170 363862 22226
rect 363918 22170 363986 22226
rect 364042 22170 394582 22226
rect 394638 22170 394706 22226
rect 394762 22170 425302 22226
rect 425358 22170 425426 22226
rect 425482 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 170518 22102
rect 170574 22046 170642 22102
rect 170698 22046 201238 22102
rect 201294 22046 201362 22102
rect 201418 22046 231958 22102
rect 232014 22046 232082 22102
rect 232138 22046 262678 22102
rect 262734 22046 262802 22102
rect 262858 22046 271702 22102
rect 271758 22046 271826 22102
rect 271882 22046 302422 22102
rect 302478 22046 302546 22102
rect 302602 22046 333142 22102
rect 333198 22046 333266 22102
rect 333322 22046 363862 22102
rect 363918 22046 363986 22102
rect 364042 22046 394582 22102
rect 394638 22046 394706 22102
rect 394762 22046 425302 22102
rect 425358 22046 425426 22102
rect 425482 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 170518 21978
rect 170574 21922 170642 21978
rect 170698 21922 201238 21978
rect 201294 21922 201362 21978
rect 201418 21922 231958 21978
rect 232014 21922 232082 21978
rect 232138 21922 262678 21978
rect 262734 21922 262802 21978
rect 262858 21922 271702 21978
rect 271758 21922 271826 21978
rect 271882 21922 302422 21978
rect 302478 21922 302546 21978
rect 302602 21922 333142 21978
rect 333198 21922 333266 21978
rect 333322 21922 363862 21978
rect 363918 21922 363986 21978
rect 364042 21922 394582 21978
rect 394638 21922 394706 21978
rect 394762 21922 425302 21978
rect 425358 21922 425426 21978
rect 425482 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect 241932 21358 266660 21374
rect 241932 21302 241948 21358
rect 242004 21302 266588 21358
rect 266644 21302 266660 21358
rect 241932 21286 266660 21302
rect 240588 21178 270356 21194
rect 240588 21122 240604 21178
rect 240660 21122 270284 21178
rect 270340 21122 270356 21178
rect 240588 21106 270356 21122
rect 240364 20998 270580 21014
rect 240364 20942 240380 20998
rect 240436 20942 270508 20998
rect 270564 20942 270580 20998
rect 240364 20926 270580 20942
rect 264668 20098 273492 20114
rect 264668 20042 264684 20098
rect 264740 20042 273420 20098
rect 273476 20042 273492 20098
rect 264668 20026 273492 20042
rect 432668 20098 587204 20114
rect 432668 20042 432684 20098
rect 432740 20042 587132 20098
rect 587188 20042 587204 20098
rect 432668 20026 587204 20042
rect 231180 19918 242020 19934
rect 231180 19862 231196 19918
rect 231252 19862 241948 19918
rect 242004 19862 242020 19918
rect 231180 19846 242020 19862
rect 243724 19918 266772 19934
rect 243724 19862 243740 19918
rect 243796 19862 266700 19918
rect 266756 19862 266772 19918
rect 243724 19846 266772 19862
rect 241932 19738 273268 19754
rect 241932 19682 241948 19738
rect 242004 19682 273196 19738
rect 273252 19682 273268 19738
rect 241932 19666 273268 19682
rect 239244 19558 271364 19574
rect 239244 19502 239260 19558
rect 239316 19502 271292 19558
rect 271348 19502 271364 19558
rect 239244 19486 271364 19502
rect 236556 19378 273044 19394
rect 236556 19322 236572 19378
rect 236628 19322 272972 19378
rect 273028 19322 273044 19378
rect 236556 19306 273044 19322
rect 245068 17578 266436 17594
rect 245068 17522 245084 17578
rect 245140 17522 266364 17578
rect 266420 17522 266436 17578
rect 245068 17506 266436 17522
rect 230732 17218 257028 17234
rect 230732 17162 230748 17218
rect 230804 17162 256956 17218
rect 257012 17162 257028 17218
rect 230732 17146 257028 17162
rect 236780 17038 273380 17054
rect 236780 16982 236796 17038
rect 236852 16982 273308 17038
rect 273364 16982 273380 17038
rect 236780 16966 273380 16982
rect 226252 16858 272932 16874
rect 226252 16802 226268 16858
rect 226324 16802 272860 16858
rect 272916 16802 272932 16858
rect 226252 16786 272932 16802
rect 4156 16678 152084 16694
rect 4156 16622 4172 16678
rect 4228 16622 152012 16678
rect 152068 16622 152084 16678
rect 4156 16606 152084 16622
rect 245292 16318 268228 16334
rect 245292 16262 245308 16318
rect 245364 16262 268156 16318
rect 268212 16262 268228 16318
rect 245292 16246 268228 16262
rect 269036 16318 273268 16334
rect 269036 16262 269052 16318
rect 269108 16262 273196 16318
rect 273252 16262 273268 16318
rect 269036 16246 273268 16262
rect 217292 16138 272260 16154
rect 217292 16082 217308 16138
rect 217364 16082 272188 16138
rect 272244 16082 272260 16138
rect 217292 16066 272260 16082
rect 226028 15958 267892 15974
rect 226028 15902 226044 15958
rect 226100 15902 267820 15958
rect 267876 15902 267892 15958
rect 226028 15886 267892 15902
rect 436588 15958 581380 15974
rect 436588 15902 436604 15958
rect 436660 15902 581308 15958
rect 581364 15902 581380 15958
rect 436588 15886 581380 15902
rect 238572 15238 272148 15254
rect 238572 15182 238588 15238
rect 238644 15182 272076 15238
rect 272132 15182 272148 15238
rect 238572 15166 272148 15182
rect 243052 14338 268452 14354
rect 243052 14282 243068 14338
rect 243124 14282 268380 14338
rect 268436 14282 268452 14338
rect 243052 14266 268452 14282
rect 221324 13978 268676 13994
rect 221324 13922 221340 13978
rect 221396 13922 268604 13978
rect 268660 13922 268676 13978
rect 221324 13906 268676 13922
rect 222220 13798 273044 13814
rect 222220 13742 222236 13798
rect 222292 13742 272972 13798
rect 273028 13742 273044 13798
rect 222220 13726 273044 13742
rect 23420 13618 187140 13634
rect 23420 13562 23436 13618
rect 23492 13562 187068 13618
rect 187124 13562 187140 13618
rect 23420 13546 187140 13562
rect 218636 13618 274164 13634
rect 218636 13562 218652 13618
rect 218708 13562 274092 13618
rect 274148 13562 274164 13618
rect 218636 13546 274164 13562
rect 169580 13438 209764 13454
rect 169580 13382 169596 13438
rect 169652 13382 209692 13438
rect 209748 13382 209764 13438
rect 169580 13366 209764 13382
rect 210124 13438 268004 13454
rect 210124 13382 210140 13438
rect 210196 13382 267932 13438
rect 267988 13382 268004 13438
rect 210124 13366 268004 13382
rect 424156 13438 428276 13454
rect 424156 13382 424172 13438
rect 424228 13382 428204 13438
rect 428260 13382 428276 13438
rect 424156 13366 428276 13382
rect 209900 13258 268340 13274
rect 209900 13202 209916 13258
rect 209972 13202 268268 13258
rect 268324 13202 268340 13258
rect 209900 13186 268340 13202
rect 209452 13078 269012 13094
rect 209452 13022 209468 13078
rect 209524 13022 268940 13078
rect 268996 13022 269012 13078
rect 209452 13006 269012 13022
rect 245964 12898 270020 12914
rect 245964 12842 245980 12898
rect 246036 12842 269948 12898
rect 270004 12842 270020 12898
rect 245964 12826 270020 12842
rect 265452 12538 273156 12554
rect 265452 12482 265468 12538
rect 265524 12482 273084 12538
rect 273140 12482 273156 12538
rect 265452 12466 273156 12482
rect 134412 11998 190612 12014
rect 134412 11942 134428 11998
rect 134484 11942 190540 11998
rect 190596 11942 190612 11998
rect 134412 11926 190612 11942
rect 44476 11818 186916 11834
rect 44476 11762 44492 11818
rect 44548 11762 186844 11818
rect 186900 11762 186916 11818
rect 44476 11746 186916 11762
rect 243500 11818 273492 11834
rect 243500 11762 243516 11818
rect 243572 11762 273420 11818
rect 273476 11762 273492 11818
rect 243500 11746 273492 11762
rect 236108 11638 273940 11654
rect 236108 11582 236124 11638
rect 236180 11582 273868 11638
rect 273924 11582 273940 11638
rect 236108 11566 273940 11582
rect 241484 11458 269684 11474
rect 241484 11402 241500 11458
rect 241556 11402 269612 11458
rect 269668 11402 269684 11458
rect 241484 11386 269684 11402
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 221996 9658 289060 9674
rect 221996 9602 222012 9658
rect 222068 9602 288988 9658
rect 289044 9602 289060 9658
rect 221996 9586 289060 9602
rect 242380 9478 531204 9494
rect 242380 9422 242396 9478
rect 242452 9422 531132 9478
rect 531188 9422 531204 9478
rect 242380 9406 531204 9422
rect 17260 9298 186244 9314
rect 17260 9242 17276 9298
rect 17332 9242 186172 9298
rect 186228 9242 186244 9298
rect 17260 9226 186244 9242
rect 231404 9298 571300 9314
rect 231404 9242 231420 9298
rect 231476 9242 571228 9298
rect 571284 9242 571300 9298
rect 231404 9226 571300 9242
rect 288972 8578 523588 8594
rect 288972 8522 523516 8578
rect 523572 8522 523588 8578
rect 288972 8506 523588 8522
rect 288972 8414 289060 8506
rect 226588 8398 289060 8414
rect 226588 8342 226604 8398
rect 226660 8342 289060 8398
rect 226588 8326 289060 8342
rect 238236 8038 479796 8054
rect 238236 7982 238252 8038
rect 238308 7982 479724 8038
rect 479780 7982 479796 8038
rect 238236 7966 479796 7982
rect 241036 7858 540724 7874
rect 241036 7802 241052 7858
rect 241108 7802 540652 7858
rect 540708 7802 540724 7858
rect 241036 7786 540724 7802
rect 55340 7678 190500 7694
rect 55340 7622 55356 7678
rect 55412 7622 190428 7678
rect 190484 7622 190500 7678
rect 55340 7606 190500 7622
rect 228380 7678 546436 7694
rect 228380 7622 228396 7678
rect 228452 7622 546364 7678
rect 546420 7622 546436 7678
rect 228380 7606 546436 7622
rect 41788 7498 188260 7514
rect 41788 7442 41804 7498
rect 41860 7442 188188 7498
rect 188244 7442 188260 7498
rect 41788 7426 188260 7442
rect 230060 7498 557860 7514
rect 230060 7442 230076 7498
rect 230132 7442 557788 7498
rect 557844 7442 557860 7498
rect 230060 7426 557860 7442
rect 231740 6598 394116 6614
rect 231740 6542 231756 6598
rect 231812 6542 394044 6598
rect 394100 6542 394116 6598
rect 231740 6526 394116 6542
rect 223340 6418 506452 6434
rect 223340 6362 223356 6418
rect 223412 6362 506380 6418
rect 506436 6362 506452 6418
rect 223340 6346 506452 6362
rect 225020 6238 512164 6254
rect 225020 6182 225036 6238
rect 225092 6182 512092 6238
rect 512148 6182 512164 6238
rect 225020 6166 512164 6182
rect 26780 6058 186580 6074
rect 26780 6002 26796 6058
rect 26852 6002 186508 6058
rect 186564 6002 186580 6058
rect 26780 5986 186580 6002
rect 224908 6058 517876 6074
rect 224908 6002 224924 6058
rect 224980 6002 517804 6058
rect 517860 6002 517876 6058
rect 224908 5986 517876 6002
rect 11548 5878 185012 5894
rect 11548 5822 11564 5878
rect 11620 5822 184940 5878
rect 184996 5822 185012 5878
rect 11548 5806 185012 5822
rect 226700 5878 535012 5894
rect 226700 5822 226716 5878
rect 226772 5822 534940 5878
rect 534996 5822 535012 5878
rect 226700 5806 535012 5822
rect 246860 4978 571300 4994
rect 246860 4922 246876 4978
rect 246932 4922 571228 4978
rect 571284 4922 571300 4978
rect 246860 4906 571300 4922
rect 245068 4798 559764 4814
rect 245068 4742 245084 4798
rect 245140 4742 559692 4798
rect 559748 4742 559764 4798
rect 245068 4726 559764 4742
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect 13340 3358 185124 3374
rect 13340 3302 13356 3358
rect 13412 3302 185052 3358
rect 185108 3302 185124 3358
rect 13340 3286 185124 3302
rect 245180 3358 552708 3374
rect 245180 3302 245196 3358
rect 245252 3302 552636 3358
rect 552692 3302 552708 3358
rect 245180 3286 552708 3302
rect 241708 3178 515972 3194
rect 241708 3122 241724 3178
rect 241780 3122 515900 3178
rect 515956 3122 515972 3178
rect 241708 3106 515972 3122
rect 273404 2998 542740 3014
rect 273404 2942 273420 2998
rect 273476 2942 542668 2998
rect 542724 2942 542740 2998
rect 273404 2926 542740 2942
rect 238348 2818 265540 2834
rect 238348 2762 238364 2818
rect 238420 2762 265468 2818
rect 265524 2762 265540 2818
rect 238348 2746 265540 2762
rect 270380 2818 475988 2834
rect 270380 2762 270396 2818
rect 270452 2762 475916 2818
rect 475972 2762 475988 2818
rect 270380 2746 475988 2762
rect 267132 2638 304180 2654
rect 267132 2582 267148 2638
rect 267204 2582 304108 2638
rect 304164 2582 304180 2638
rect 267132 2566 304180 2582
rect 240028 2458 277300 2474
rect 240028 2402 240044 2458
rect 240100 2402 277228 2458
rect 277284 2402 277300 2458
rect 240028 2386 277300 2402
rect 238460 838 474084 854
rect 238460 782 238476 838
rect 238532 782 474012 838
rect 474068 782 474084 838
rect 238460 766 474084 782
rect 240140 658 485620 674
rect 240140 602 240156 658
rect 240212 602 485548 658
rect 485604 602 485620 658
rect 240140 586 485620 602
rect 271276 478 554052 494
rect 271276 422 271292 478
rect 271348 422 553980 478
rect 554036 422 554052 478
rect 271276 406 554052 422
rect 243276 298 527396 314
rect 243276 242 243292 298
rect 243348 242 527324 298
rect 527380 242 527396 298
rect 243276 226 527396 242
rect 243388 118 533108 134
rect 243388 62 243404 118
rect 243460 62 533036 118
rect 533092 62 533108 118
rect 243388 46 533108 62
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use logo  logo
timestamp 0
transform 1 0 20000 0 1 578000
box -2000 -2000 150000 18000
use core0  mprj_core0
timestamp 0
transform 1 0 174000 0 1 99000
box 802 3076 98560 200000
use core1  mprj_core1
timestamp 0
transform 1 0 320000 0 1 99000
box 914 3076 98560 200000
use dcache  mprj_dcache
timestamp 0
transform 1 0 18000 0 1 395000
box 1258 0 534662 178958
use icache  mprj_icache_0
timestamp 0
transform -1 0 150000 0 1 20000
box 0 1138 138862 350508
use icache  mprj_icache_1
timestamp 0
transform 1 0 444000 0 1 20000
box 0 1138 138862 350508
use int_ram  mprj_int_ram
timestamp 0
transform -1 0 430000 0 1 10000
box 1258 578 160000 67966
use interconnect_inner  mprj_interconnect_inner
timestamp 0
transform 1 0 174000 0 1 308000
box 0 0 240000 74000
use interconnect_outer  mprj_interconnect_outer
timestamp 0
transform 1 0 166000 0 1 16000
box 0 0 100000 60000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 393242 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 19842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 74766 190358 104970 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 575846 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 19842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 74766 221078 104970 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 575846 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 19842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 74766 251798 104970 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 575846 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 79630 282518 306466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 575846 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 79630 313238 306466 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 575846 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 575846 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 575846 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 8578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 575846 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 393242 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 575846 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 575846 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 575846 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 575846 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 19026 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 372094 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 17816 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s 170184 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 372094 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 393242 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 19842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 74766 194078 99964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 575846 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 19842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 74766 224798 99964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 575846 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 19842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 74766 255518 99964 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 575846 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 79630 286238 306466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 575846 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 79630 316958 306466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 575846 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 79630 347678 102954 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 297430 347678 306466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 575846 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 79630 378398 102954 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 297430 378398 306466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 575846 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 79630 409118 102954 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 297430 409118 306466 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 575846 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 393242 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 575846 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 575846 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 575846 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 575846 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 19026 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 372094 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 17816 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s 170184 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 262830 58322 262830 58322 0 vdd
rlabel via4 247470 64322 247470 64322 0 vss
rlabel metal2 261016 85134 261016 85134 0 io_in[0]
rlabel metal3 593026 403592 593026 403592 0 io_in[10]
rlabel metal2 238840 77854 238840 77854 0 io_in[11]
rlabel metal2 236824 78022 236824 78022 0 io_in[12]
rlabel metal3 593250 522536 593250 522536 0 io_in[13]
rlabel metal3 593138 562184 593138 562184 0 io_in[14]
rlabel metal4 425880 229335 425880 229335 0 io_in[15]
rlabel metal2 518728 593306 518728 593306 0 io_in[16]
rlabel metal2 452536 593138 452536 593138 0 io_in[17]
rlabel metal2 309176 94192 309176 94192 0 io_in[18]
rlabel metal3 27272 389816 27272 389816 0 io_in[19]
rlabel metal3 592858 46760 592858 46760 0 io_in[1]
rlabel metal3 164122 69608 164122 69608 0 io_in[20]
rlabel metal2 46984 377776 46984 377776 0 io_in[21]
rlabel metal4 29400 475944 29400 475944 0 io_in[22]
rlabel metal2 55160 593250 55160 593250 0 io_in[23]
rlabel metal3 1918 587160 1918 587160 0 io_in[24]
rlabel metal3 2310 544824 2310 544824 0 io_in[25]
rlabel metal3 2422 502488 2422 502488 0 io_in[26]
rlabel metal3 164122 50792 164122 50792 0 io_in[27]
rlabel metal3 2198 417816 2198 417816 0 io_in[28]
rlabel metal4 163688 46648 163688 46648 0 io_in[29]
rlabel metal4 256984 80209 256984 80209 0 io_in[2]
rlabel metal3 3990 333144 3990 333144 0 io_in[30]
rlabel metal2 3528 20552 3528 20552 0 io_in[31]
rlabel metal3 164472 18200 164472 18200 0 io_in[32]
rlabel metal3 4214 206136 4214 206136 0 io_in[33]
rlabel metal3 164962 31976 164962 31976 0 io_in[34]
rlabel metal3 4326 121464 4326 121464 0 io_in[35]
rlabel metal3 165186 26600 165186 26600 0 io_in[36]
rlabel metal4 4928 26010 4928 26010 0 io_in[37]
rlabel metal3 593362 126056 593362 126056 0 io_in[3]
rlabel metal3 593250 165704 593250 165704 0 io_in[4]
rlabel metal3 593138 205352 593138 205352 0 io_in[5]
rlabel metal3 593082 245000 593082 245000 0 io_in[6]
rlabel metal3 591402 284648 591402 284648 0 io_in[7]
rlabel metal3 593306 324520 593306 324520 0 io_in[8]
rlabel metal2 242872 86254 242872 86254 0 io_in[9]
rlabel metal4 259672 84977 259672 84977 0 io_oeb[0]
rlabel metal3 593306 430136 593306 430136 0 io_oeb[10]
rlabel metal3 593082 469672 593082 469672 0 io_oeb[11]
rlabel metal2 235480 87094 235480 87094 0 io_oeb[12]
rlabel metal3 593194 548968 593194 548968 0 io_oeb[13]
rlabel metal3 593082 588616 593082 588616 0 io_oeb[14]
rlabel metal2 540792 593362 540792 593362 0 io_oeb[15]
rlabel metal2 474600 593194 474600 593194 0 io_oeb[16]
rlabel metal3 282352 245224 282352 245224 0 io_oeb[17]
rlabel metal3 28224 377944 28224 377944 0 io_oeb[18]
rlabel metal3 167664 359576 167664 359576 0 io_oeb[19]
rlabel metal3 593418 73192 593418 73192 0 io_oeb[1]
rlabel metal3 164234 67816 164234 67816 0 io_oeb[20]
rlabel metal2 143416 593082 143416 593082 0 io_oeb[21]
rlabel metal2 77336 593194 77336 593194 0 io_oeb[22]
rlabel metal3 166376 60046 166376 60046 0 io_oeb[23]
rlabel metal3 4256 403256 4256 403256 0 io_oeb[24]
rlabel metal3 2366 516600 2366 516600 0 io_oeb[25]
rlabel metal3 2590 474264 2590 474264 0 io_oeb[26]
rlabel metal3 164066 49000 164066 49000 0 io_oeb[27]
rlabel metal3 165298 46312 165298 46312 0 io_oeb[28]
rlabel metal3 2310 347480 2310 347480 0 io_oeb[29]
rlabel metal2 255640 83342 255640 83342 0 io_oeb[2]
rlabel metal3 165018 40936 165018 40936 0 io_oeb[30]
rlabel metal3 2310 262584 2310 262584 0 io_oeb[31]
rlabel metal3 4102 220248 4102 220248 0 io_oeb[32]
rlabel metal3 2422 177912 2422 177912 0 io_oeb[33]
rlabel metal3 2534 135576 2534 135576 0 io_oeb[34]
rlabel metal3 165130 27496 165130 27496 0 io_oeb[35]
rlabel metal4 4816 26190 4816 26190 0 io_oeb[36]
rlabel metal3 2310 8792 2310 8792 0 io_oeb[37]
rlabel metal3 593306 152488 593306 152488 0 io_oeb[3]
rlabel metal3 593250 192136 593250 192136 0 io_oeb[4]
rlabel metal3 593194 231896 593194 231896 0 io_oeb[5]
rlabel metal3 591514 271432 591514 271432 0 io_oeb[6]
rlabel metal3 593082 311304 593082 311304 0 io_oeb[7]
rlabel metal3 593250 350952 593250 350952 0 io_oeb[8]
rlabel metal2 241710 75880 241710 75880 0 io_oeb[9]
rlabel metal3 593474 20328 593474 20328 0 io_out[0]
rlabel metal2 240184 77910 240184 77910 0 io_out[10]
rlabel metal2 238350 75880 238350 75880 0 io_out[11]
rlabel metal3 593362 496104 593362 496104 0 io_out[12]
rlabel metal3 234640 80584 234640 80584 0 io_out[13]
rlabel metal4 232120 85247 232120 85247 0 io_out[14]
rlabel metal2 562632 488138 562632 488138 0 io_out[15]
rlabel metal2 496664 593250 496664 593250 0 io_out[16]
rlabel metal2 430472 593082 430472 593082 0 io_out[17]
rlabel metal3 546112 374584 546112 374584 0 io_out[18]
rlabel metal2 48664 381752 48664 381752 0 io_out[19]
rlabel metal2 258328 85918 258328 85918 0 io_out[1]
rlabel metal2 48664 375872 48664 375872 0 io_out[20]
rlabel metal3 163800 590184 163800 590184 0 io_out[21]
rlabel metal2 99288 593138 99288 593138 0 io_out[22]
rlabel metal3 164906 60648 164906 60648 0 io_out[23]
rlabel metal3 165018 57960 165018 57960 0 io_out[24]
rlabel metal3 164962 55272 164962 55272 0 io_out[25]
rlabel metal3 165914 52584 165914 52584 0 io_out[26]
rlabel metal3 164906 49896 164906 49896 0 io_out[27]
rlabel metal3 2702 403704 2702 403704 0 io_out[28]
rlabel metal3 2310 361592 2310 361592 0 io_out[29]
rlabel metal3 591570 99624 591570 99624 0 io_out[2]
rlabel metal4 4200 16697 4200 16697 0 io_out[30]
rlabel metal3 1470 276696 1470 276696 0 io_out[31]
rlabel metal3 2366 234360 2366 234360 0 io_out[32]
rlabel metal3 3318 192024 3318 192024 0 io_out[33]
rlabel metal3 4368 26600 4368 26600 0 io_out[34]
rlabel metal3 165018 28392 165018 28392 0 io_out[35]
rlabel metal3 4648 26376 4648 26376 0 io_out[36]
rlabel metal3 2702 22680 2702 22680 0 io_out[37]
rlabel metal3 591738 139272 591738 139272 0 io_out[3]
rlabel metal3 591458 178920 591458 178920 0 io_out[4]
rlabel metal3 591626 218568 591626 218568 0 io_out[5]
rlabel metal3 591402 258216 591402 258216 0 io_out[6]
rlabel metal3 593194 298088 593194 298088 0 io_out[7]
rlabel metal3 593138 337624 593138 337624 0 io_out[8]
rlabel metal3 242872 80584 242872 80584 0 io_out[9]
rlabel metal3 211792 4200 211792 4200 0 la_data_in[0]
rlabel metal2 217112 14658 217112 14658 0 la_data_in[10]
rlabel metal2 217784 13706 217784 13706 0 la_data_in[11]
rlabel metal2 281736 3654 281736 3654 0 la_data_in[12]
rlabel metal2 280504 2632 280504 2632 0 la_data_in[13]
rlabel metal3 281232 8120 281232 8120 0 la_data_in[14]
rlabel metal2 265496 1736 265496 1736 0 la_data_in[15]
rlabel metal2 280840 6664 280840 6664 0 la_data_in[16]
rlabel metal2 280392 1904 280392 1904 0 la_data_in[17]
rlabel metal2 265720 13104 265720 13104 0 la_data_in[18]
rlabel metal2 305704 1736 305704 1736 0 la_data_in[19]
rlabel metal3 214984 11592 214984 11592 0 la_data_in[1]
rlabel metal2 327432 2366 327432 2366 0 la_data_in[20]
rlabel metal2 333144 2478 333144 2478 0 la_data_in[21]
rlabel metal2 282184 2688 282184 2688 0 la_data_in[22]
rlabel metal2 344568 2534 344568 2534 0 la_data_in[23]
rlabel metal2 350280 3374 350280 3374 0 la_data_in[24]
rlabel metal2 355992 1750 355992 1750 0 la_data_in[25]
rlabel metal2 289016 8512 289016 8512 0 la_data_in[26]
rlabel metal2 307384 4144 307384 4144 0 la_data_in[27]
rlabel metal2 265720 3416 265720 3416 0 la_data_in[28]
rlabel metal2 265608 2912 265608 2912 0 la_data_in[29]
rlabel metal2 211736 11074 211736 11074 0 la_data_in[2]
rlabel metal2 384440 448 384440 448 0 la_data_in[30]
rlabel metal4 241976 20610 241976 20610 0 la_data_in[31]
rlabel metal3 234360 616 234360 616 0 la_data_in[32]
rlabel metal2 401912 3374 401912 3374 0 la_data_in[33]
rlabel metal2 407624 2422 407624 2422 0 la_data_in[34]
rlabel metal2 233240 9058 233240 9058 0 la_data_in[35]
rlabel metal2 233688 8778 233688 8778 0 la_data_in[36]
rlabel metal3 424200 4200 424200 4200 0 la_data_in[37]
rlabel metal2 234584 8722 234584 8722 0 la_data_in[38]
rlabel metal2 235032 9674 235032 9674 0 la_data_in[39]
rlabel metal2 212408 13762 212408 13762 0 la_data_in[3]
rlabel metal2 235480 8610 235480 8610 0 la_data_in[40]
rlabel metal2 235928 9394 235928 9394 0 la_data_in[41]
rlabel metal3 236376 336 236376 336 0 la_data_in[42]
rlabel metal2 240520 12712 240520 12712 0 la_data_in[43]
rlabel metal3 237832 11816 237832 11816 0 la_data_in[44]
rlabel metal2 470232 518 470232 518 0 la_data_in[45]
rlabel metal4 475944 2263 475944 2263 0 la_data_in[46]
rlabel metal3 240296 16632 240296 16632 0 la_data_in[47]
rlabel metal2 239064 14378 239064 14378 0 la_data_in[48]
rlabel metal2 239512 10514 239512 10514 0 la_data_in[49]
rlabel metal2 236040 2310 236040 2310 0 la_data_in[4]
rlabel metal3 240072 16744 240072 16744 0 la_data_in[50]
rlabel metal4 240408 18857 240408 18857 0 la_data_in[51]
rlabel metal2 240856 14490 240856 14490 0 la_data_in[52]
rlabel metal4 515928 2443 515928 2443 0 la_data_in[53]
rlabel metal3 517944 6776 517944 6776 0 la_data_in[54]
rlabel metal3 242760 12376 242760 12376 0 la_data_in[55]
rlabel metal3 243040 11816 243040 11816 0 la_data_in[56]
rlabel metal4 243096 14631 243096 14631 0 la_data_in[57]
rlabel metal2 243432 12152 243432 12152 0 la_data_in[58]
rlabel metal2 265496 4928 265496 4928 0 la_data_in[59]
rlabel metal2 235144 6216 235144 6216 0 la_data_in[5]
rlabel metal4 552664 3373 552664 3373 0 la_data_in[60]
rlabel metal4 429240 54320 429240 54320 0 la_data_in[61]
rlabel metal2 567336 8246 567336 8246 0 la_data_in[62]
rlabel metal3 354872 97720 354872 97720 0 la_data_in[63]
rlabel metal2 214424 11186 214424 11186 0 la_data_in[6]
rlabel metal2 215096 14042 215096 14042 0 la_data_in[7]
rlabel metal2 215768 15162 215768 15162 0 la_data_in[8]
rlabel metal3 218232 13440 218232 13440 0 la_data_in[9]
rlabel metal3 212856 6776 212856 6776 0 la_data_out[0]
rlabel via4 217336 16091 217336 16091 0 la_data_out[10]
rlabel metal2 218008 11130 218008 11130 0 la_data_out[11]
rlabel metal2 283640 4326 283640 4326 0 la_data_out[12]
rlabel metal2 219352 9338 219352 9338 0 la_data_out[13]
rlabel metal2 220024 15498 220024 15498 0 la_data_out[14]
rlabel metal2 300776 3094 300776 3094 0 la_data_out[15]
rlabel metal2 306712 462 306712 462 0 la_data_out[16]
rlabel metal3 420336 285656 420336 285656 0 la_data_out[17]
rlabel metal4 426776 153944 426776 153944 0 la_data_out[18]
rlabel metal4 422184 43232 422184 43232 0 la_data_out[19]
rlabel metal2 211288 12698 211288 12698 0 la_data_out[1]
rlabel metal2 329560 2366 329560 2366 0 la_data_out[20]
rlabel metal2 335272 2478 335272 2478 0 la_data_out[21]
rlabel metal2 218456 299838 218456 299838 0 la_data_out[22]
rlabel metal4 420728 50512 420728 50512 0 la_data_out[23]
rlabel metal2 352408 2254 352408 2254 0 la_data_out[24]
rlabel metal2 233688 301518 233688 301518 0 la_data_out[25]
rlabel metal2 238168 300846 238168 300846 0 la_data_out[26]
rlabel metal4 421848 45024 421848 45024 0 la_data_out[27]
rlabel metal2 375256 2030 375256 2030 0 la_data_out[28]
rlabel metal2 380968 4158 380968 4158 0 la_data_out[29]
rlabel metal2 211960 14434 211960 14434 0 la_data_out[2]
rlabel metal2 256214 298872 256214 298872 0 la_data_out[30]
rlabel metal2 260568 299838 260568 299838 0 la_data_out[31]
rlabel metal2 397992 4214 397992 4214 0 la_data_out[32]
rlabel metal2 403816 4270 403816 4270 0 la_data_out[33]
rlabel metal3 421736 4256 421736 4256 0 la_data_out[34]
rlabel metal4 428456 151872 428456 151872 0 la_data_out[35]
rlabel metal2 420952 2254 420952 2254 0 la_data_out[36]
rlabel metal2 426664 2310 426664 2310 0 la_data_out[37]
rlabel metal2 218008 299166 218008 299166 0 la_data_out[38]
rlabel metal3 437360 4200 437360 4200 0 la_data_out[39]
rlabel metal2 212632 12642 212632 12642 0 la_data_out[3]
rlabel metal2 443576 45262 443576 45262 0 la_data_out[40]
rlabel metal2 449288 4270 449288 4270 0 la_data_out[41]
rlabel metal2 455000 2646 455000 2646 0 la_data_out[42]
rlabel metal4 437864 159199 437864 159199 0 la_data_out[43]
rlabel metal2 466424 2590 466424 2590 0 la_data_out[44]
rlabel metal4 310856 301171 310856 301171 0 la_data_out[45]
rlabel metal2 477848 2478 477848 2478 0 la_data_out[46]
rlabel metal4 260120 297584 260120 297584 0 la_data_out[47]
rlabel metal2 320936 3808 320936 3808 0 la_data_out[48]
rlabel metal2 308280 2520 308280 2520 0 la_data_out[49]
rlabel metal2 237944 4270 237944 4270 0 la_data_out[4]
rlabel metal2 500696 4158 500696 4158 0 la_data_out[50]
rlabel metal4 506408 4903 506408 4903 0 la_data_out[51]
rlabel metal4 512120 4813 512120 4813 0 la_data_out[52]
rlabel metal4 517832 4723 517832 4723 0 la_data_out[53]
rlabel metal2 523544 2366 523544 2366 0 la_data_out[54]
rlabel metal2 282184 81032 282184 81032 0 la_data_out[55]
rlabel metal4 534968 4633 534968 4633 0 la_data_out[56]
rlabel metal4 540680 5903 540680 5903 0 la_data_out[57]
rlabel metal4 546392 5757 546392 5757 0 la_data_out[58]
rlabel metal2 444136 52696 444136 52696 0 la_data_out[59]
rlabel metal2 236824 6216 236824 6216 0 la_data_out[5]
rlabel metal4 557816 5611 557816 5611 0 la_data_out[60]
rlabel metal2 431256 48496 431256 48496 0 la_data_out[61]
rlabel metal4 256984 17807 256984 17807 0 la_data_out[62]
rlabel metal4 571256 8023 571256 8023 0 la_data_out[63]
rlabel metal2 214648 15778 214648 15778 0 la_data_out[6]
rlabel metal2 215320 15834 215320 15834 0 la_data_out[7]
rlabel metal2 215992 15946 215992 15946 0 la_data_out[8]
rlabel metal3 231840 16128 231840 16128 0 la_data_out[9]
rlabel metal3 213920 4312 213920 4312 0 la_oenb[0]
rlabel metal3 217560 16856 217560 16856 0 la_oenb[10]
rlabel metal2 279832 2646 279832 2646 0 la_oenb[11]
rlabel metal2 285488 504 285488 504 0 la_oenb[12]
rlabel metal2 219576 11018 219576 11018 0 la_oenb[13]
rlabel metal3 286160 4424 286160 4424 0 la_oenb[14]
rlabel metal2 285656 6664 285656 6664 0 la_oenb[15]
rlabel metal2 308392 3486 308392 3486 0 la_oenb[16]
rlabel metal4 222264 14361 222264 14361 0 la_oenb[17]
rlabel metal2 319816 4214 319816 4214 0 la_oenb[18]
rlabel metal3 288148 3752 288148 3752 0 la_oenb[19]
rlabel metal2 211512 11242 211512 11242 0 la_oenb[1]
rlabel metal2 331240 4998 331240 4998 0 la_oenb[20]
rlabel metal2 336952 4942 336952 4942 0 la_oenb[21]
rlabel metal2 225624 12698 225624 12698 0 la_oenb[22]
rlabel metal2 289128 7616 289128 7616 0 la_oenb[23]
rlabel metal2 265832 5544 265832 5544 0 la_oenb[24]
rlabel metal2 359800 3262 359800 3262 0 la_oenb[25]
rlabel metal4 238616 13681 238616 13681 0 la_oenb[26]
rlabel metal3 275464 5320 275464 5320 0 la_oenb[27]
rlabel metal2 376936 4158 376936 4158 0 la_oenb[28]
rlabel metal2 382648 4102 382648 4102 0 la_oenb[29]
rlabel metal2 212184 14378 212184 14378 0 la_oenb[2]
rlabel metal2 388360 3150 388360 3150 0 la_oenb[30]
rlabel metal4 394072 4993 394072 4993 0 la_oenb[31]
rlabel metal2 234920 10976 234920 10976 0 la_oenb[32]
rlabel metal2 405496 1694 405496 1694 0 la_oenb[33]
rlabel metal3 235424 12264 235424 12264 0 la_oenb[34]
rlabel metal2 425096 5768 425096 5768 0 la_oenb[35]
rlabel metal3 422296 4200 422296 4200 0 la_oenb[36]
rlabel metal2 428456 4046 428456 4046 0 la_oenb[37]
rlabel metal3 241976 12320 241976 12320 0 la_oenb[38]
rlabel metal2 235256 14658 235256 14658 0 la_oenb[39]
rlabel metal2 234136 2366 234136 2366 0 la_oenb[3]
rlabel metal2 445480 3990 445480 3990 0 la_oenb[40]
rlabel metal2 451192 3206 451192 3206 0 la_oenb[41]
rlabel metal4 236600 18047 236600 18047 0 la_oenb[42]
rlabel metal2 237048 13818 237048 13818 0 la_oenb[43]
rlabel metal2 237496 11242 237496 11242 0 la_oenb[44]
rlabel metal4 474040 713 474040 713 0 la_oenb[45]
rlabel metal4 238336 12150 238336 12150 0 la_oenb[46]
rlabel metal3 239512 11816 239512 11816 0 la_oenb[47]
rlabel metal4 239288 18137 239288 18137 0 la_oenb[48]
rlabel metal2 496888 2422 496888 2422 0 la_oenb[49]
rlabel metal2 239848 2534 239848 2534 0 la_oenb[4]
rlabel metal4 240128 12150 240128 12150 0 la_oenb[50]
rlabel metal4 240632 18947 240632 18947 0 la_oenb[51]
rlabel metal2 241080 12138 241080 12138 0 la_oenb[52]
rlabel metal4 241528 12407 241528 12407 0 la_oenb[53]
rlabel metal2 241976 10458 241976 10458 0 la_oenb[54]
rlabel metal4 242424 11137 242424 11137 0 la_oenb[55]
rlabel metal2 352744 3472 352744 3472 0 la_oenb[56]
rlabel metal4 542696 2353 542696 2353 0 la_oenb[57]
rlabel metal2 548296 2366 548296 2366 0 la_oenb[58]
rlabel metal4 554008 533 554008 533 0 la_oenb[59]
rlabel metal2 214200 11914 214200 11914 0 la_oenb[5]
rlabel metal4 559720 4093 559720 4093 0 la_oenb[60]
rlabel metal2 565432 8302 565432 8302 0 la_oenb[61]
rlabel metal4 571256 4183 571256 4183 0 la_oenb[62]
rlabel metal4 429688 51128 429688 51128 0 la_oenb[63]
rlabel metal2 214872 10962 214872 10962 0 la_oenb[6]
rlabel metal2 233464 6048 233464 6048 0 la_oenb[7]
rlabel metal2 262696 2366 262696 2366 0 la_oenb[8]
rlabel metal3 216888 16912 216888 16912 0 la_oenb[9]
rlabel metal2 171640 188286 171640 188286 0 mprj/c0_clk
rlabel metal2 191128 306530 191128 306530 0 mprj/c0_disable
rlabel metal2 185752 302246 185752 302246 0 mprj/c0_i_core_int_sreg\[0\]
rlabel metal2 238616 300622 238616 300622 0 mprj/c0_i_core_int_sreg\[10\]
rlabel metal2 243096 301014 243096 301014 0 mprj/c0_i_core_int_sreg\[11\]
rlabel metal2 247576 301014 247576 301014 0 mprj/c0_i_core_int_sreg\[12\]
rlabel metal2 252224 305480 252224 305480 0 mprj/c0_i_core_int_sreg\[13\]
rlabel metal2 256802 308056 256802 308056 0 mprj/c0_i_core_int_sreg\[14\]
rlabel metal2 260694 308056 260694 308056 0 mprj/c0_i_core_int_sreg\[15\]
rlabel metal2 191702 298872 191702 298872 0 mprj/c0_i_core_int_sreg\[1\]
rlabel metal2 208600 305018 208600 305018 0 mprj/c0_i_core_int_sreg\[2\]
rlabel metal2 213080 306026 213080 306026 0 mprj/c0_i_core_int_sreg\[3\]
rlabel metal2 217560 304850 217560 304850 0 mprj/c0_i_core_int_sreg\[4\]
rlabel metal2 213528 300678 213528 300678 0 mprj/c0_i_core_int_sreg\[5\]
rlabel metal2 218904 300566 218904 300566 0 mprj/c0_i_core_int_sreg\[6\]
rlabel metal3 227752 305256 227752 305256 0 mprj/c0_i_core_int_sreg\[7\]
rlabel metal2 235480 305858 235480 305858 0 mprj/c0_i_core_int_sreg\[8\]
rlabel metal2 234262 298872 234262 298872 0 mprj/c0_i_core_int_sreg\[9\]
rlabel metal2 191576 304794 191576 304794 0 mprj/c0_i_irq
rlabel metal2 192024 305802 192024 305802 0 mprj/c0_i_mc_core_int
rlabel metal2 192472 305746 192472 305746 0 mprj/c0_i_mem_ack
rlabel metal2 186200 300566 186200 300566 0 mprj/c0_i_mem_data\[0\]
rlabel metal2 239064 300566 239064 300566 0 mprj/c0_i_mem_data\[10\]
rlabel metal2 243544 301070 243544 301070 0 mprj/c0_i_mem_data\[11\]
rlabel metal2 248024 301070 248024 301070 0 mprj/c0_i_mem_data\[12\]
rlabel metal3 253176 304024 253176 304024 0 mprj/c0_i_mem_data\[13\]
rlabel metal2 257250 308056 257250 308056 0 mprj/c0_i_mem_data\[14\]
rlabel metal2 261142 308056 261142 308056 0 mprj/c0_i_mem_data\[15\]
rlabel metal2 192024 300958 192024 300958 0 mprj/c0_i_mem_data\[1\]
rlabel metal2 209048 305858 209048 305858 0 mprj/c0_i_mem_data\[2\]
rlabel metal2 213528 306754 213528 306754 0 mprj/c0_i_mem_data\[3\]
rlabel metal2 208600 299838 208600 299838 0 mprj/c0_i_mem_data\[4\]
rlabel metal2 214102 298872 214102 298872 0 mprj/c0_i_mem_data\[5\]
rlabel metal2 219352 301462 219352 301462 0 mprj/c0_i_mem_data\[6\]
rlabel metal3 228088 303912 228088 303912 0 mprj/c0_i_mem_data\[7\]
rlabel metal2 235592 305816 235592 305816 0 mprj/c0_i_mem_data\[8\]
rlabel metal2 234710 298872 234710 298872 0 mprj/c0_i_mem_data\[9\]
rlabel metal2 192920 306474 192920 306474 0 mprj/c0_i_mem_exception
rlabel metal2 186648 301462 186648 301462 0 mprj/c0_i_req_data\[0\]
rlabel metal2 239512 300510 239512 300510 0 mprj/c0_i_req_data\[10\]
rlabel metal2 243992 301630 243992 301630 0 mprj/c0_i_req_data\[11\]
rlabel metal2 250712 304514 250712 304514 0 mprj/c0_i_req_data\[12\]
rlabel metal3 253624 303912 253624 303912 0 mprj/c0_i_req_data\[13\]
rlabel metal2 257698 308056 257698 308056 0 mprj/c0_i_req_data\[14\]
rlabel metal2 261590 308056 261590 308056 0 mprj/c0_i_req_data\[15\]
rlabel metal2 264278 308056 264278 308056 0 mprj/c0_i_req_data\[16\]
rlabel metal2 264726 308056 264726 308056 0 mprj/c0_i_req_data\[17\]
rlabel metal2 265384 305256 265384 305256 0 mprj/c0_i_req_data\[18\]
rlabel metal2 265622 308056 265622 308056 0 mprj/c0_i_req_data\[19\]
rlabel metal2 192472 301014 192472 301014 0 mprj/c0_i_req_data\[1\]
rlabel metal2 266070 308056 266070 308056 0 mprj/c0_i_req_data\[20\]
rlabel metal2 266518 308056 266518 308056 0 mprj/c0_i_req_data\[21\]
rlabel metal2 267064 306908 267064 306908 0 mprj/c0_i_req_data\[22\]
rlabel metal2 267414 308056 267414 308056 0 mprj/c0_i_req_data\[23\]
rlabel metal2 267862 308056 267862 308056 0 mprj/c0_i_req_data\[24\]
rlabel metal2 268310 308056 268310 308056 0 mprj/c0_i_req_data\[25\]
rlabel metal2 268800 305144 268800 305144 0 mprj/c0_i_req_data\[26\]
rlabel metal2 269206 308056 269206 308056 0 mprj/c0_i_req_data\[27\]
rlabel metal2 269654 308056 269654 308056 0 mprj/c0_i_req_data\[28\]
rlabel metal2 270102 308056 270102 308056 0 mprj/c0_i_req_data\[29\]
rlabel metal2 209496 306698 209496 306698 0 mprj/c0_i_req_data\[2\]
rlabel metal2 270648 305368 270648 305368 0 mprj/c0_i_req_data\[30\]
rlabel metal2 270998 308056 270998 308056 0 mprj/c0_i_req_data\[31\]
rlabel metal2 213976 305354 213976 305354 0 mprj/c0_i_req_data\[3\]
rlabel metal3 213808 304696 213808 304696 0 mprj/c0_i_req_data\[4\]
rlabel metal2 214550 298872 214550 298872 0 mprj/c0_i_req_data\[5\]
rlabel metal2 219800 300286 219800 300286 0 mprj/c0_i_req_data\[6\]
rlabel metal2 231896 306138 231896 306138 0 mprj/c0_i_req_data\[7\]
rlabel metal2 236376 306418 236376 306418 0 mprj/c0_i_req_data\[8\]
rlabel metal2 235032 301350 235032 301350 0 mprj/c0_i_req_data\[9\]
rlabel metal2 193368 304850 193368 304850 0 mprj/c0_i_req_data_valid
rlabel metal2 193816 305970 193816 305970 0 mprj/c0_o_c_data_page
rlabel metal2 194264 305914 194264 305914 0 mprj/c0_o_c_instr_long
rlabel metal2 194712 305858 194712 305858 0 mprj/c0_o_c_instr_page
rlabel metal2 195160 304962 195160 304962 0 mprj/c0_o_icache_flush
rlabel metal3 189448 303128 189448 303128 0 mprj/c0_o_instr_long_addr\[0\]
rlabel metal2 192920 301798 192920 301798 0 mprj/c0_o_instr_long_addr\[1\]
rlabel metal2 209944 306586 209944 306586 0 mprj/c0_o_instr_long_addr\[2\]
rlabel metal2 214424 305970 214424 305970 0 mprj/c0_o_instr_long_addr\[3\]
rlabel metal3 214200 304808 214200 304808 0 mprj/c0_o_instr_long_addr\[4\]
rlabel metal2 214872 300398 214872 300398 0 mprj/c0_o_instr_long_addr\[5\]
rlabel metal2 220248 300454 220248 300454 0 mprj/c0_o_instr_long_addr\[6\]
rlabel metal2 232344 306194 232344 306194 0 mprj/c0_o_instr_long_addr\[7\]
rlabel metal2 187544 299446 187544 299446 0 mprj/c0_o_mem_addr\[0\]
rlabel metal2 240086 298872 240086 298872 0 mprj/c0_o_mem_addr\[10\]
rlabel metal2 244440 301686 244440 301686 0 mprj/c0_o_mem_addr\[11\]
rlabel metal2 251160 305914 251160 305914 0 mprj/c0_o_mem_addr\[12\]
rlabel metal3 254072 303800 254072 303800 0 mprj/c0_o_mem_addr\[13\]
rlabel metal2 258146 308056 258146 308056 0 mprj/c0_o_mem_addr\[14\]
rlabel metal2 262080 305144 262080 305144 0 mprj/c0_o_mem_addr\[15\]
rlabel metal2 193494 298872 193494 298872 0 mprj/c0_o_mem_addr\[1\]
rlabel metal2 210392 305634 210392 305634 0 mprj/c0_o_mem_addr\[2\]
rlabel metal2 214872 305466 214872 305466 0 mprj/c0_o_mem_addr\[3\]
rlabel metal3 214592 305368 214592 305368 0 mprj/c0_o_mem_addr\[4\]
rlabel metal2 215446 298872 215446 298872 0 mprj/c0_o_mem_addr\[5\]
rlabel metal2 220696 300510 220696 300510 0 mprj/c0_o_mem_addr\[6\]
rlabel metal2 232792 306250 232792 306250 0 mprj/c0_o_mem_addr\[7\]
rlabel metal2 236824 305018 236824 305018 0 mprj/c0_o_mem_addr\[8\]
rlabel metal2 235480 301182 235480 301182 0 mprj/c0_o_mem_addr\[9\]
rlabel metal2 187992 302190 187992 302190 0 mprj/c0_o_mem_addr_high\[0\]
rlabel metal2 193816 301182 193816 301182 0 mprj/c0_o_mem_addr_high\[1\]
rlabel metal2 211288 306530 211288 306530 0 mprj/c0_o_mem_addr_high\[2\]
rlabel metal2 215768 305690 215768 305690 0 mprj/c0_o_mem_addr_high\[3\]
rlabel metal2 210462 298872 210462 298872 0 mprj/c0_o_mem_addr_high\[4\]
rlabel metal2 215894 298872 215894 298872 0 mprj/c0_o_mem_addr_high\[5\]
rlabel metal2 221144 299950 221144 299950 0 mprj/c0_o_mem_addr_high\[6\]
rlabel metal2 233688 306306 233688 306306 0 mprj/c0_o_mem_addr_high\[7\]
rlabel metal2 188440 300174 188440 300174 0 mprj/c0_o_mem_data\[0\]
rlabel metal2 240408 300454 240408 300454 0 mprj/c0_o_mem_data\[10\]
rlabel metal2 244888 300622 244888 300622 0 mprj/c0_o_mem_data\[11\]
rlabel metal2 251608 306026 251608 306026 0 mprj/c0_o_mem_data\[12\]
rlabel metal2 254408 303576 254408 303576 0 mprj/c0_o_mem_data\[13\]
rlabel metal2 258776 305214 258776 305214 0 mprj/c0_o_mem_data\[14\]
rlabel metal2 262486 308056 262486 308056 0 mprj/c0_o_mem_data\[15\]
rlabel metal2 194264 300062 194264 300062 0 mprj/c0_o_mem_data\[1\]
rlabel metal2 210840 305914 210840 305914 0 mprj/c0_o_mem_data\[2\]
rlabel metal2 215320 305578 215320 305578 0 mprj/c0_o_mem_data\[3\]
rlabel metal3 215320 303240 215320 303240 0 mprj/c0_o_mem_data\[4\]
rlabel metal2 216216 301406 216216 301406 0 mprj/c0_o_mem_data\[5\]
rlabel metal3 225176 303240 225176 303240 0 mprj/c0_o_mem_data\[6\]
rlabel metal2 232904 305256 232904 305256 0 mprj/c0_o_mem_data\[7\]
rlabel metal2 237272 306698 237272 306698 0 mprj/c0_o_mem_data\[8\]
rlabel metal2 235928 301462 235928 301462 0 mprj/c0_o_mem_data\[9\]
rlabel metal2 195608 305018 195608 305018 0 mprj/c0_o_mem_long
rlabel metal2 196056 306586 196056 306586 0 mprj/c0_o_mem_req
rlabel metal2 188888 300622 188888 300622 0 mprj/c0_o_mem_sel\[0\]
rlabel metal2 194712 300230 194712 300230 0 mprj/c0_o_mem_sel\[1\]
rlabel metal2 196504 306642 196504 306642 0 mprj/c0_o_mem_we
rlabel metal2 196952 306698 196952 306698 0 mprj/c0_o_req_active
rlabel metal2 189336 302302 189336 302302 0 mprj/c0_o_req_addr\[0\]
rlabel metal2 240856 300398 240856 300398 0 mprj/c0_o_req_addr\[10\]
rlabel metal2 245336 300958 245336 300958 0 mprj/c0_o_req_addr\[11\]
rlabel metal2 252056 304402 252056 304402 0 mprj/c0_o_req_addr\[12\]
rlabel metal2 255640 305354 255640 305354 0 mprj/c0_o_req_addr\[13\]
rlabel metal2 259042 308056 259042 308056 0 mprj/c0_o_req_addr\[14\]
rlabel metal2 262934 308056 262934 308056 0 mprj/c0_o_req_addr\[15\]
rlabel metal2 195160 300118 195160 300118 0 mprj/c0_o_req_addr\[1\]
rlabel metal2 211736 304906 211736 304906 0 mprj/c0_o_req_addr\[2\]
rlabel metal2 216216 306810 216216 306810 0 mprj/c0_o_req_addr\[3\]
rlabel metal2 211288 301742 211288 301742 0 mprj/c0_o_req_addr\[4\]
rlabel metal2 216664 301350 216664 301350 0 mprj/c0_o_req_addr\[5\]
rlabel metal3 225848 305144 225848 305144 0 mprj/c0_o_req_addr\[6\]
rlabel metal2 234136 304682 234136 304682 0 mprj/c0_o_req_addr\[7\]
rlabel metal2 231896 299838 231896 299838 0 mprj/c0_o_req_addr\[8\]
rlabel metal2 236502 298872 236502 298872 0 mprj/c0_o_req_addr\[9\]
rlabel metal2 197330 308056 197330 308056 0 mprj/c0_o_req_ppl_submit
rlabel metal2 197848 305634 197848 305634 0 mprj/c0_rst
rlabel metal2 189784 301854 189784 301854 0 mprj/c0_sr_bus_addr\[0\]
rlabel metal2 241304 301798 241304 301798 0 mprj/c0_sr_bus_addr\[10\]
rlabel metal2 245784 300566 245784 300566 0 mprj/c0_sr_bus_addr\[11\]
rlabel metal2 252434 308056 252434 308056 0 mprj/c0_sr_bus_addr\[12\]
rlabel metal2 256088 305410 256088 305410 0 mprj/c0_sr_bus_addr\[13\]
rlabel metal2 259490 308056 259490 308056 0 mprj/c0_sr_bus_addr\[14\]
rlabel metal2 263382 308056 263382 308056 0 mprj/c0_sr_bus_addr\[15\]
rlabel metal2 195608 300286 195608 300286 0 mprj/c0_sr_bus_addr\[1\]
rlabel metal2 212184 304962 212184 304962 0 mprj/c0_sr_bus_addr\[2\]
rlabel metal2 216664 306866 216664 306866 0 mprj/c0_sr_bus_addr\[3\]
rlabel metal2 211862 298872 211862 298872 0 mprj/c0_sr_bus_addr\[4\]
rlabel metal2 217112 300342 217112 300342 0 mprj/c0_sr_bus_addr\[5\]
rlabel metal3 226296 303464 226296 303464 0 mprj/c0_sr_bus_addr\[6\]
rlabel metal2 234584 304906 234584 304906 0 mprj/c0_sr_bus_addr\[7\]
rlabel metal3 235256 303352 235256 303352 0 mprj/c0_sr_bus_addr\[8\]
rlabel metal2 236754 298872 236754 298872 0 mprj/c0_sr_bus_addr\[9\]
rlabel metal2 190232 300510 190232 300510 0 mprj/c0_sr_bus_data_o\[0\]
rlabel metal2 241822 298872 241822 298872 0 mprj/c0_sr_bus_data_o\[10\]
rlabel metal2 246232 300510 246232 300510 0 mprj/c0_sr_bus_data_o\[11\]
rlabel metal3 251776 303912 251776 303912 0 mprj/c0_sr_bus_data_o\[12\]
rlabel metal2 256536 305466 256536 305466 0 mprj/c0_sr_bus_data_o\[13\]
rlabel metal2 259938 308056 259938 308056 0 mprj/c0_sr_bus_data_o\[14\]
rlabel metal2 263760 305256 263760 305256 0 mprj/c0_sr_bus_data_o\[15\]
rlabel metal2 196056 301742 196056 301742 0 mprj/c0_sr_bus_data_o\[1\]
rlabel metal2 212632 306642 212632 306642 0 mprj/c0_sr_bus_data_o\[2\]
rlabel metal2 217112 305074 217112 305074 0 mprj/c0_sr_bus_data_o\[3\]
rlabel metal2 212310 298872 212310 298872 0 mprj/c0_sr_bus_data_o\[4\]
rlabel metal2 217686 298872 217686 298872 0 mprj/c0_sr_bus_data_o\[5\]
rlabel metal2 222936 299894 222936 299894 0 mprj/c0_sr_bus_data_o\[6\]
rlabel metal2 234962 308056 234962 308056 0 mprj/c0_sr_bus_data_o\[7\]
rlabel metal2 232918 298872 232918 298872 0 mprj/c0_sr_bus_data_o\[8\]
rlabel metal2 237272 300062 237272 300062 0 mprj/c0_sr_bus_data_o\[9\]
rlabel metal2 198296 305690 198296 305690 0 mprj/c0_sr_bus_we
rlabel metal2 220024 85470 220024 85470 0 mprj/c1_clk
rlabel metal2 310296 303954 310296 303954 0 mprj/c1_dbg_pc\[0\]
rlabel metal2 383656 303030 383656 303030 0 mprj/c1_dbg_pc\[10\]
rlabel metal2 388136 299838 388136 299838 0 mprj/c1_dbg_pc\[11\]
rlabel metal2 372120 307258 372120 307258 0 mprj/c1_dbg_pc\[12\]
rlabel metal2 376600 307538 376600 307538 0 mprj/c1_dbg_pc\[13\]
rlabel metal4 381080 305267 381080 305267 0 mprj/c1_dbg_pc\[14\]
rlabel metal2 406056 302918 406056 302918 0 mprj/c1_dbg_pc\[15\]
rlabel metal2 336616 303142 336616 303142 0 mprj/c1_dbg_pc\[1\]
rlabel metal2 321944 307538 321944 307538 0 mprj/c1_dbg_pc\[2\]
rlabel metal4 327320 304457 327320 304457 0 mprj/c1_dbg_pc\[3\]
rlabel metal2 332696 307426 332696 307426 0 mprj/c1_dbg_pc\[4\]
rlabel metal2 338072 307706 338072 307706 0 mprj/c1_dbg_pc\[5\]
rlabel metal2 343448 307538 343448 307538 0 mprj/c1_dbg_pc\[6\]
rlabel metal2 348824 307314 348824 307314 0 mprj/c1_dbg_pc\[7\]
rlabel metal2 354200 307426 354200 307426 0 mprj/c1_dbg_pc\[8\]
rlabel metal2 379176 302918 379176 302918 0 mprj/c1_dbg_pc\[9\]
rlabel metal2 310744 307482 310744 307482 0 mprj/c1_dbg_r0\[0\]
rlabel metal2 384104 302582 384104 302582 0 mprj/c1_dbg_r0\[10\]
rlabel metal2 368088 304066 368088 304066 0 mprj/c1_dbg_r0\[11\]
rlabel metal2 372568 307314 372568 307314 0 mprj/c1_dbg_r0\[12\]
rlabel metal2 377048 303954 377048 303954 0 mprj/c1_dbg_r0\[13\]
rlabel metal2 381528 307370 381528 307370 0 mprj/c1_dbg_r0\[14\]
rlabel metal2 406504 299726 406504 299726 0 mprj/c1_dbg_r0\[15\]
rlabel metal2 337064 302694 337064 302694 0 mprj/c1_dbg_r0\[1\]
rlabel metal2 322392 307650 322392 307650 0 mprj/c1_dbg_r0\[2\]
rlabel metal2 327768 307314 327768 307314 0 mprj/c1_dbg_r0\[3\]
rlabel metal2 333144 303954 333144 303954 0 mprj/c1_dbg_r0\[4\]
rlabel metal2 338520 305858 338520 305858 0 mprj/c1_dbg_r0\[5\]
rlabel metal2 343896 307650 343896 307650 0 mprj/c1_dbg_r0\[6\]
rlabel metal2 349272 304178 349272 304178 0 mprj/c1_dbg_r0\[7\]
rlabel metal2 354648 307370 354648 307370 0 mprj/c1_dbg_r0\[8\]
rlabel metal2 379624 301238 379624 301238 0 mprj/c1_dbg_r0\[9\]
rlabel metal2 302680 306474 302680 306474 0 mprj/c1_disable
rlabel metal2 311192 307426 311192 307426 0 mprj/c1_i_core_int_sreg\[0\]
rlabel metal2 384552 301350 384552 301350 0 mprj/c1_i_core_int_sreg\[10\]
rlabel metal2 371336 303520 371336 303520 0 mprj/c1_i_core_int_sreg\[11\]
rlabel metal2 373016 306474 373016 306474 0 mprj/c1_i_core_int_sreg\[12\]
rlabel metal2 377496 305634 377496 305634 0 mprj/c1_i_core_int_sreg\[13\]
rlabel metal2 381976 305802 381976 305802 0 mprj/c1_i_core_int_sreg\[14\]
rlabel metal2 406952 301294 406952 301294 0 mprj/c1_i_core_int_sreg\[15\]
rlabel metal2 337512 299502 337512 299502 0 mprj/c1_i_core_int_sreg\[1\]
rlabel metal2 322840 304178 322840 304178 0 mprj/c1_i_core_int_sreg\[2\]
rlabel metal2 328216 305746 328216 305746 0 mprj/c1_i_core_int_sreg\[3\]
rlabel metal2 333592 305802 333592 305802 0 mprj/c1_i_core_int_sreg\[4\]
rlabel metal2 338968 305914 338968 305914 0 mprj/c1_i_core_int_sreg\[5\]
rlabel metal4 344344 301799 344344 301799 0 mprj/c1_i_core_int_sreg\[6\]
rlabel metal2 349720 305634 349720 305634 0 mprj/c1_i_core_int_sreg\[7\]
rlabel metal2 355096 305746 355096 305746 0 mprj/c1_i_core_int_sreg\[8\]
rlabel metal2 380072 301294 380072 301294 0 mprj/c1_i_core_int_sreg\[9\]
rlabel metal2 303128 304850 303128 304850 0 mprj/c1_i_irq
rlabel metal2 303576 305746 303576 305746 0 mprj/c1_i_mc_core_int
rlabel metal4 309176 303617 309176 303617 0 mprj/c1_i_mem_ack
rlabel metal2 311640 305914 311640 305914 0 mprj/c1_i_mem_data\[0\]
rlabel metal4 385000 298144 385000 298144 0 mprj/c1_i_mem_data\[10\]
rlabel metal2 368984 305970 368984 305970 0 mprj/c1_i_mem_data\[11\]
rlabel metal2 373464 305690 373464 305690 0 mprj/c1_i_mem_data\[12\]
rlabel metal4 379624 304727 379624 304727 0 mprj/c1_i_mem_data\[13\]
rlabel metal2 382424 307426 382424 307426 0 mprj/c1_i_mem_data\[14\]
rlabel metal2 407400 301462 407400 301462 0 mprj/c1_i_mem_data\[15\]
rlabel metal2 317464 303058 317464 303058 0 mprj/c1_i_mem_data\[1\]
rlabel metal2 323288 305578 323288 305578 0 mprj/c1_i_mem_data\[2\]
rlabel metal2 328664 305634 328664 305634 0 mprj/c1_i_mem_data\[3\]
rlabel metal4 336056 303741 336056 303741 0 mprj/c1_i_mem_data\[4\]
rlabel metal2 339416 307594 339416 307594 0 mprj/c1_i_mem_data\[5\]
rlabel metal2 344792 306026 344792 306026 0 mprj/c1_i_mem_data\[6\]
rlabel metal2 350168 307258 350168 307258 0 mprj/c1_i_mem_data\[7\]
rlabel metal2 376040 301014 376040 301014 0 mprj/c1_i_mem_data\[8\]
rlabel metal2 380520 303142 380520 303142 0 mprj/c1_i_mem_data\[9\]
rlabel metal2 304472 305858 304472 305858 0 mprj/c1_i_mem_exception
rlabel metal2 312088 305802 312088 305802 0 mprj/c1_i_req_data\[0\]
rlabel metal3 370440 302904 370440 302904 0 mprj/c1_i_req_data\[10\]
rlabel metal4 369432 304817 369432 304817 0 mprj/c1_i_req_data\[11\]
rlabel metal2 376264 304024 376264 304024 0 mprj/c1_i_req_data\[12\]
rlabel metal2 398888 303478 398888 303478 0 mprj/c1_i_req_data\[13\]
rlabel metal2 382872 304122 382872 304122 0 mprj/c1_i_req_data\[14\]
rlabel metal2 407848 300958 407848 300958 0 mprj/c1_i_req_data\[15\]
rlabel metal2 390040 305914 390040 305914 0 mprj/c1_i_req_data\[16\]
rlabel metal2 390488 304066 390488 304066 0 mprj/c1_i_req_data\[17\]
rlabel metal2 390936 305970 390936 305970 0 mprj/c1_i_req_data\[18\]
rlabel metal4 398104 303576 398104 303576 0 mprj/c1_i_req_data\[19\]
rlabel metal2 317912 307594 317912 307594 0 mprj/c1_i_req_data\[1\]
rlabel metal2 391832 307146 391832 307146 0 mprj/c1_i_req_data\[20\]
rlabel metal2 392280 307594 392280 307594 0 mprj/c1_i_req_data\[21\]
rlabel metal2 392728 306866 392728 306866 0 mprj/c1_i_req_data\[22\]
rlabel metal2 393176 306698 393176 306698 0 mprj/c1_i_req_data\[23\]
rlabel metal2 393624 306754 393624 306754 0 mprj/c1_i_req_data\[24\]
rlabel metal2 394072 306810 394072 306810 0 mprj/c1_i_req_data\[25\]
rlabel metal4 394520 304233 394520 304233 0 mprj/c1_i_req_data\[26\]
rlabel metal2 394968 305746 394968 305746 0 mprj/c1_i_req_data\[27\]
rlabel metal2 395416 306530 395416 306530 0 mprj/c1_i_req_data\[28\]
rlabel metal2 395864 306642 395864 306642 0 mprj/c1_i_req_data\[29\]
rlabel metal4 329224 303632 329224 303632 0 mprj/c1_i_req_data\[2\]
rlabel metal2 396312 305690 396312 305690 0 mprj/c1_i_req_data\[30\]
rlabel metal2 396760 306474 396760 306474 0 mprj/c1_i_req_data\[31\]
rlabel metal4 330904 304615 330904 304615 0 mprj/c1_i_req_data\[3\]
rlabel metal2 334488 305522 334488 305522 0 mprj/c1_i_req_data\[4\]
rlabel metal2 339864 305970 339864 305970 0 mprj/c1_i_req_data\[5\]
rlabel metal2 345240 305690 345240 305690 0 mprj/c1_i_req_data\[6\]
rlabel metal2 350616 304122 350616 304122 0 mprj/c1_i_req_data\[7\]
rlabel metal2 355992 306866 355992 306866 0 mprj/c1_i_req_data\[8\]
rlabel metal2 380968 299726 380968 299726 0 mprj/c1_i_req_data\[9\]
rlabel metal2 304920 307370 304920 307370 0 mprj/c1_i_req_data_valid
rlabel metal2 305368 307314 305368 307314 0 mprj/c1_o_c_data_page
rlabel metal2 305816 305634 305816 305634 0 mprj/c1_o_c_instr_long
rlabel metal2 306264 304794 306264 304794 0 mprj/c1_o_c_instr_page
rlabel metal4 310856 305133 310856 305133 0 mprj/c1_o_icache_flush
rlabel metal2 312536 305970 312536 305970 0 mprj/c1_o_instr_long_addr\[0\]
rlabel metal2 318360 306026 318360 306026 0 mprj/c1_o_instr_long_addr\[1\]
rlabel metal4 324184 305267 324184 305267 0 mprj/c1_o_instr_long_addr\[2\]
rlabel metal2 329560 304122 329560 304122 0 mprj/c1_o_instr_long_addr\[3\]
rlabel metal2 334936 307482 334936 307482 0 mprj/c1_o_instr_long_addr\[4\]
rlabel metal2 340312 304010 340312 304010 0 mprj/c1_o_instr_long_addr\[5\]
rlabel metal2 345688 307202 345688 307202 0 mprj/c1_o_instr_long_addr\[6\]
rlabel metal2 371448 305172 371448 305172 0 mprj/c1_o_instr_long_addr\[7\]
rlabel metal2 312984 304906 312984 304906 0 mprj/c1_o_mem_addr\[0\]
rlabel metal2 385896 299670 385896 299670 0 mprj/c1_o_mem_addr\[10\]
rlabel metal2 369880 304010 369880 304010 0 mprj/c1_o_mem_addr\[11\]
rlabel metal4 374360 301945 374360 301945 0 mprj/c1_o_mem_addr\[12\]
rlabel metal2 378840 307650 378840 307650 0 mprj/c1_o_mem_addr\[13\]
rlabel metal2 383320 307706 383320 307706 0 mprj/c1_o_mem_addr\[14\]
rlabel metal3 391328 304808 391328 304808 0 mprj/c1_o_mem_addr\[15\]
rlabel metal2 318808 304010 318808 304010 0 mprj/c1_o_mem_addr\[1\]
rlabel metal4 324632 304547 324632 304547 0 mprj/c1_o_mem_addr\[2\]
rlabel metal2 330008 307370 330008 307370 0 mprj/c1_o_mem_addr\[3\]
rlabel metal4 336504 305357 336504 305357 0 mprj/c1_o_mem_addr\[4\]
rlabel metal2 340830 308056 340830 308056 0 mprj/c1_o_mem_addr\[5\]
rlabel metal2 346136 304066 346136 304066 0 mprj/c1_o_mem_addr\[6\]
rlabel metal2 351512 306306 351512 306306 0 mprj/c1_o_mem_addr\[7\]
rlabel metal2 376936 299894 376936 299894 0 mprj/c1_o_mem_addr\[8\]
rlabel metal4 381416 303349 381416 303349 0 mprj/c1_o_mem_addr\[9\]
rlabel metal2 313880 304234 313880 304234 0 mprj/c1_o_mem_addr_high\[0\]
rlabel metal3 331800 305368 331800 305368 0 mprj/c1_o_mem_addr_high\[1\]
rlabel metal2 325528 306362 325528 306362 0 mprj/c1_o_mem_addr_high\[2\]
rlabel metal2 330904 306194 330904 306194 0 mprj/c1_o_mem_addr_high\[3\]
rlabel metal2 336280 306698 336280 306698 0 mprj/c1_o_mem_addr_high\[4\]
rlabel metal4 354424 303520 354424 303520 0 mprj/c1_o_mem_addr_high\[5\]
rlabel metal2 347032 306810 347032 306810 0 mprj/c1_o_mem_addr_high\[6\]
rlabel metal4 352408 304907 352408 304907 0 mprj/c1_o_mem_addr_high\[7\]
rlabel metal2 313432 306810 313432 306810 0 mprj/c1_o_mem_data\[0\]
rlabel metal4 371112 303352 371112 303352 0 mprj/c1_o_mem_data\[10\]
rlabel metal2 370328 306810 370328 306810 0 mprj/c1_o_mem_data\[11\]
rlabel metal2 374808 307202 374808 307202 0 mprj/c1_o_mem_data\[12\]
rlabel metal2 379288 304794 379288 304794 0 mprj/c1_o_mem_data\[13\]
rlabel metal2 383768 304906 383768 304906 0 mprj/c1_o_mem_data\[14\]
rlabel metal2 388248 304178 388248 304178 0 mprj/c1_o_mem_data\[15\]
rlabel metal2 319256 305690 319256 305690 0 mprj/c1_o_mem_data\[1\]
rlabel metal2 325080 306474 325080 306474 0 mprj/c1_o_mem_data\[2\]
rlabel metal4 330456 304907 330456 304907 0 mprj/c1_o_mem_data\[3\]
rlabel metal2 335832 304794 335832 304794 0 mprj/c1_o_mem_data\[4\]
rlabel metal3 355320 305088 355320 305088 0 mprj/c1_o_mem_data\[5\]
rlabel metal2 346584 306474 346584 306474 0 mprj/c1_o_mem_data\[6\]
rlabel metal2 351960 306138 351960 306138 0 mprj/c1_o_mem_data\[7\]
rlabel metal2 377384 299838 377384 299838 0 mprj/c1_o_mem_data\[8\]
rlabel metal2 381864 300118 381864 300118 0 mprj/c1_o_mem_data\[9\]
rlabel metal2 307160 306586 307160 306586 0 mprj/c1_o_mem_long
rlabel metal2 307608 306698 307608 306698 0 mprj/c1_o_mem_req
rlabel metal2 334824 301966 334824 301966 0 mprj/c1_o_mem_sel\[0\]
rlabel metal3 321832 305256 321832 305256 0 mprj/c1_o_mem_sel\[1\]
rlabel metal2 308056 306754 308056 306754 0 mprj/c1_o_mem_we
rlabel metal2 308504 306866 308504 306866 0 mprj/c1_o_req_active
rlabel metal2 335272 300566 335272 300566 0 mprj/c1_o_req_addr\[0\]
rlabel metal2 386792 302134 386792 302134 0 mprj/c1_o_req_addr\[10\]
rlabel metal2 370776 306530 370776 306530 0 mprj/c1_o_req_addr\[11\]
rlabel metal2 375256 306418 375256 306418 0 mprj/c1_o_req_addr\[12\]
rlabel metal2 379736 304962 379736 304962 0 mprj/c1_o_req_addr\[13\]
rlabel metal2 384216 306250 384216 306250 0 mprj/c1_o_req_addr\[14\]
rlabel metal2 402360 303576 402360 303576 0 mprj/c1_o_req_addr\[15\]
rlabel metal2 320600 305018 320600 305018 0 mprj/c1_o_req_addr\[1\]
rlabel metal2 335048 304640 335048 304640 0 mprj/c1_o_req_addr\[2\]
rlabel metal3 332808 305144 332808 305144 0 mprj/c1_o_req_addr\[3\]
rlabel metal2 336728 306418 336728 306418 0 mprj/c1_o_req_addr\[4\]
rlabel metal3 344960 305144 344960 305144 0 mprj/c1_o_req_addr\[5\]
rlabel metal2 347480 304738 347480 304738 0 mprj/c1_o_req_addr\[6\]
rlabel metal2 352856 304850 352856 304850 0 mprj/c1_o_req_addr\[7\]
rlabel metal2 377832 300454 377832 300454 0 mprj/c1_o_req_addr\[8\]
rlabel metal2 382312 299894 382312 299894 0 mprj/c1_o_req_addr\[9\]
rlabel metal2 308952 306362 308952 306362 0 mprj/c1_o_req_ppl_submit
rlabel metal2 309400 304682 309400 304682 0 mprj/c1_rst
rlabel metal4 331016 304248 331016 304248 0 mprj/c1_sr_bus_addr\[0\]
rlabel metal4 383096 303576 383096 303576 0 mprj/c1_sr_bus_addr\[10\]
rlabel metal2 371042 308056 371042 308056 0 mprj/c1_sr_bus_addr\[11\]
rlabel metal3 376656 304024 376656 304024 0 mprj/c1_sr_bus_addr\[12\]
rlabel metal2 380184 306306 380184 306306 0 mprj/c1_sr_bus_addr\[13\]
rlabel metal2 384664 305018 384664 305018 0 mprj/c1_sr_bus_addr\[14\]
rlabel metal2 389144 306586 389144 306586 0 mprj/c1_sr_bus_addr\[15\]
rlabel metal3 321832 302456 321832 302456 0 mprj/c1_sr_bus_addr\[1\]
rlabel metal2 326424 306306 326424 306306 0 mprj/c1_sr_bus_addr\[2\]
rlabel metal2 331800 306810 331800 306810 0 mprj/c1_sr_bus_addr\[3\]
rlabel metal2 337176 304962 337176 304962 0 mprj/c1_sr_bus_addr\[4\]
rlabel metal4 342552 304997 342552 304997 0 mprj/c1_sr_bus_addr\[5\]
rlabel metal2 347928 306642 347928 306642 0 mprj/c1_sr_bus_addr\[6\]
rlabel metal2 353304 305018 353304 305018 0 mprj/c1_sr_bus_addr\[7\]
rlabel metal2 378280 300566 378280 300566 0 mprj/c1_sr_bus_addr\[8\]
rlabel metal2 382760 300342 382760 300342 0 mprj/c1_sr_bus_addr\[9\]
rlabel metal2 336168 299894 336168 299894 0 mprj/c1_sr_bus_data_o\[0\]
rlabel metal4 378840 305312 378840 305312 0 mprj/c1_sr_bus_data_o\[10\]
rlabel metal2 371672 306642 371672 306642 0 mprj/c1_sr_bus_data_o\[11\]
rlabel metal2 376152 304850 376152 304850 0 mprj/c1_sr_bus_data_o\[12\]
rlabel metal3 382312 304024 382312 304024 0 mprj/c1_sr_bus_data_o\[13\]
rlabel metal2 405608 303422 405608 303422 0 mprj/c1_sr_bus_data_o\[14\]
rlabel metal4 399784 301453 399784 301453 0 mprj/c1_sr_bus_data_o\[15\]
rlabel metal2 321496 305074 321496 305074 0 mprj/c1_sr_bus_data_o\[1\]
rlabel metal2 326872 304850 326872 304850 0 mprj/c1_sr_bus_data_o\[2\]
rlabel metal2 332318 308056 332318 308056 0 mprj/c1_sr_bus_data_o\[3\]
rlabel metal2 337624 304906 337624 304906 0 mprj/c1_sr_bus_data_o\[4\]
rlabel metal4 343000 304817 343000 304817 0 mprj/c1_sr_bus_data_o\[5\]
rlabel metal2 348376 304570 348376 304570 0 mprj/c1_sr_bus_data_o\[6\]
rlabel metal3 353752 305424 353752 305424 0 mprj/c1_sr_bus_data_o\[7\]
rlabel metal2 378728 300230 378728 300230 0 mprj/c1_sr_bus_data_o\[8\]
rlabel metal2 383208 299838 383208 299838 0 mprj/c1_sr_bus_data_o\[9\]
rlabel metal2 309848 304962 309848 304962 0 mprj/c1_sr_bus_we
rlabel metal2 27944 387002 27944 387002 0 mprj/dcache_clk
rlabel metal2 36008 393722 36008 393722 0 mprj/dcache_mem_ack
rlabel metal2 80360 392042 80360 392042 0 mprj/dcache_mem_addr\[0\]
rlabel metal2 316344 384566 316344 384566 0 mprj/dcache_mem_addr\[10\]
rlabel metal3 331576 386344 331576 386344 0 mprj/dcache_mem_addr\[11\]
rlabel metal2 337848 386358 337848 386358 0 mprj/dcache_mem_addr\[12\]
rlabel metal2 348600 386582 348600 386582 0 mprj/dcache_mem_addr\[13\]
rlabel metal2 359352 386302 359352 386302 0 mprj/dcache_mem_addr\[14\]
rlabel metal2 370104 385742 370104 385742 0 mprj/dcache_mem_addr\[15\]
rlabel metal2 380856 386414 380856 386414 0 mprj/dcache_mem_addr\[16\]
rlabel metal2 384440 384734 384440 384734 0 mprj/dcache_mem_addr\[17\]
rlabel metal2 499688 392154 499688 392154 0 mprj/dcache_mem_addr\[18\]
rlabel metal2 391608 384678 391608 384678 0 mprj/dcache_mem_addr\[19\]
rlabel metal2 215992 386470 215992 386470 0 mprj/dcache_mem_addr\[1\]
rlabel metal2 515816 391202 515816 391202 0 mprj/dcache_mem_addr\[20\]
rlabel metal2 398776 386358 398776 386358 0 mprj/dcache_mem_addr\[21\]
rlabel metal2 402360 385518 402360 385518 0 mprj/dcache_mem_addr\[22\]
rlabel metal2 405944 384566 405944 384566 0 mprj/dcache_mem_addr\[23\]
rlabel metal2 144872 393106 144872 393106 0 mprj/dcache_mem_addr\[2\]
rlabel metal2 169064 392826 169064 392826 0 mprj/dcache_mem_addr\[3\]
rlabel metal2 193256 392882 193256 392882 0 mprj/dcache_mem_addr\[4\]
rlabel metal2 217448 391258 217448 391258 0 mprj/dcache_mem_addr\[5\]
rlabel metal2 241640 392826 241640 392826 0 mprj/dcache_mem_addr\[6\]
rlabel metal2 265832 390306 265832 390306 0 mprj/dcache_mem_addr\[7\]
rlabel metal2 290024 393666 290024 393666 0 mprj/dcache_mem_addr\[8\]
rlabel metal2 305592 386246 305592 386246 0 mprj/dcache_mem_addr\[9\]
rlabel metal2 40040 391146 40040 391146 0 mprj/dcache_mem_cache_enable
rlabel metal2 44072 391202 44072 391202 0 mprj/dcache_mem_exception
rlabel metal2 84392 391314 84392 391314 0 mprj/dcache_mem_i_data\[0\]
rlabel metal2 318136 387086 318136 387086 0 mprj/dcache_mem_i_data\[10\]
rlabel metal2 328888 384678 328888 384678 0 mprj/dcache_mem_i_data\[11\]
rlabel metal3 342104 386008 342104 386008 0 mprj/dcache_mem_i_data\[12\]
rlabel metal3 351120 386344 351120 386344 0 mprj/dcache_mem_i_data\[13\]
rlabel metal2 361144 383334 361144 383334 0 mprj/dcache_mem_i_data\[14\]
rlabel metal2 371896 385686 371896 385686 0 mprj/dcache_mem_i_data\[15\]
rlabel metal2 116648 392098 116648 392098 0 mprj/dcache_mem_i_data\[1\]
rlabel metal2 148904 391426 148904 391426 0 mprj/dcache_mem_i_data\[2\]
rlabel metal2 242872 384902 242872 384902 0 mprj/dcache_mem_i_data\[3\]
rlabel metal2 197288 391986 197288 391986 0 mprj/dcache_mem_i_data\[4\]
rlabel metal2 264376 386358 264376 386358 0 mprj/dcache_mem_i_data\[5\]
rlabel metal2 265496 389816 265496 389816 0 mprj/dcache_mem_i_data\[6\]
rlabel metal2 285880 383782 285880 383782 0 mprj/dcache_mem_i_data\[7\]
rlabel metal3 295344 386344 295344 386344 0 mprj/dcache_mem_i_data\[8\]
rlabel metal2 307384 383726 307384 383726 0 mprj/dcache_mem_i_data\[9\]
rlabel metal2 88424 391370 88424 391370 0 mprj/dcache_mem_o_data\[0\]
rlabel metal2 319928 383726 319928 383726 0 mprj/dcache_mem_o_data\[10\]
rlabel metal2 330680 383782 330680 383782 0 mprj/dcache_mem_o_data\[11\]
rlabel metal2 341432 384566 341432 384566 0 mprj/dcache_mem_o_data\[12\]
rlabel metal2 352184 383306 352184 383306 0 mprj/dcache_mem_o_data\[13\]
rlabel metal3 365456 386232 365456 386232 0 mprj/dcache_mem_o_data\[14\]
rlabel metal2 373688 382998 373688 382998 0 mprj/dcache_mem_o_data\[15\]
rlabel metal2 120680 392154 120680 392154 0 mprj/dcache_mem_o_data\[1\]
rlabel metal2 233912 386582 233912 386582 0 mprj/dcache_mem_o_data\[2\]
rlabel metal2 177128 392210 177128 392210 0 mprj/dcache_mem_o_data\[3\]
rlabel metal2 255416 384622 255416 384622 0 mprj/dcache_mem_o_data\[4\]
rlabel metal2 266168 386414 266168 386414 0 mprj/dcache_mem_o_data\[5\]
rlabel metal2 249704 393666 249704 393666 0 mprj/dcache_mem_o_data\[6\]
rlabel metal2 287672 387086 287672 387086 0 mprj/dcache_mem_o_data\[7\]
rlabel metal2 298242 381864 298242 381864 0 mprj/dcache_mem_o_data\[8\]
rlabel metal2 309176 383782 309176 383782 0 mprj/dcache_mem_o_data\[9\]
rlabel metal2 185528 382998 185528 382998 0 mprj/dcache_mem_req
rlabel metal2 92456 389634 92456 389634 0 mprj/dcache_mem_sel\[0\]
rlabel metal2 124712 389690 124712 389690 0 mprj/dcache_mem_sel\[1\]
rlabel metal2 52136 393834 52136 393834 0 mprj/dcache_mem_we
rlabel metal2 189112 385406 189112 385406 0 mprj/dcache_rst
rlabel metal2 70504 389984 70504 389984 0 mprj/dcache_wb_4_burst
rlabel metal2 164584 391552 164584 391552 0 mprj/dcache_wb_ack
rlabel metal2 96488 394058 96488 394058 0 mprj/dcache_wb_adr\[0\]
rlabel metal2 350504 392826 350504 392826 0 mprj/dcache_wb_adr\[10\]
rlabel metal2 332472 385462 332472 385462 0 mprj/dcache_wb_adr\[11\]
rlabel metal2 398888 391482 398888 391482 0 mprj/dcache_wb_adr\[12\]
rlabel metal2 353976 383894 353976 383894 0 mprj/dcache_wb_adr\[13\]
rlabel metal2 447272 389634 447272 389634 0 mprj/dcache_wb_adr\[14\]
rlabel metal2 375480 382942 375480 382942 0 mprj/dcache_wb_adr\[15\]
rlabel metal2 382648 383950 382648 383950 0 mprj/dcache_wb_adr\[16\]
rlabel metal2 495656 390474 495656 390474 0 mprj/dcache_wb_adr\[17\]
rlabel metal2 389816 383838 389816 383838 0 mprj/dcache_wb_adr\[18\]
rlabel metal2 393400 387198 393400 387198 0 mprj/dcache_wb_adr\[19\]
rlabel metal2 186424 392168 186424 392168 0 mprj/dcache_wb_adr\[1\]
rlabel metal2 396984 387142 396984 387142 0 mprj/dcache_wb_adr\[20\]
rlabel metal2 400568 383782 400568 383782 0 mprj/dcache_wb_adr\[21\]
rlabel metal2 404152 387086 404152 387086 0 mprj/dcache_wb_adr\[22\]
rlabel metal2 407736 386638 407736 386638 0 mprj/dcache_wb_adr\[23\]
rlabel metal2 235704 388094 235704 388094 0 mprj/dcache_wb_adr\[2\]
rlabel metal3 184800 387184 184800 387184 0 mprj/dcache_wb_adr\[3\]
rlabel metal2 257208 383726 257208 383726 0 mprj/dcache_wb_adr\[4\]
rlabel metal2 238616 390880 238616 390880 0 mprj/dcache_wb_adr\[5\]
rlabel metal2 253736 392098 253736 392098 0 mprj/dcache_wb_adr\[6\]
rlabel metal2 289464 383838 289464 383838 0 mprj/dcache_wb_adr\[7\]
rlabel metal3 301168 388024 301168 388024 0 mprj/dcache_wb_adr\[8\]
rlabel metal2 310968 387310 310968 387310 0 mprj/dcache_wb_adr\[9\]
rlabel metal2 194488 383726 194488 383726 0 mprj/dcache_wb_cyc
rlabel metal2 68264 390362 68264 390362 0 mprj/dcache_wb_err
rlabel metal2 100520 393778 100520 393778 0 mprj/dcache_wb_i_dat\[0\]
rlabel metal2 334488 390040 334488 390040 0 mprj/dcache_wb_i_dat\[10\]
rlabel metal2 334264 387142 334264 387142 0 mprj/dcache_wb_i_dat\[11\]
rlabel metal2 355320 389144 355320 389144 0 mprj/dcache_wb_i_dat\[12\]
rlabel metal3 357672 386344 357672 386344 0 mprj/dcache_wb_i_dat\[13\]
rlabel metal2 446824 388416 446824 388416 0 mprj/dcache_wb_i_dat\[14\]
rlabel metal3 378000 386120 378000 386120 0 mprj/dcache_wb_i_dat\[15\]
rlabel metal2 136136 388808 136136 388808 0 mprj/dcache_wb_i_dat\[1\]
rlabel metal2 237496 387366 237496 387366 0 mprj/dcache_wb_i_dat\[2\]
rlabel metal2 185192 393722 185192 393722 0 mprj/dcache_wb_i_dat\[3\]
rlabel metal2 210056 388584 210056 388584 0 mprj/dcache_wb_i_dat\[4\]
rlabel metal2 233576 393778 233576 393778 0 mprj/dcache_wb_i_dat\[5\]
rlabel metal2 257768 391986 257768 391986 0 mprj/dcache_wb_i_dat\[6\]
rlabel metal2 281960 391146 281960 391146 0 mprj/dcache_wb_i_dat\[7\]
rlabel metal2 306152 392882 306152 392882 0 mprj/dcache_wb_i_dat\[8\]
rlabel metal2 312760 387142 312760 387142 0 mprj/dcache_wb_i_dat\[9\]
rlabel metal2 212408 383894 212408 383894 0 mprj/dcache_wb_o_dat\[0\]
rlabel metal2 358568 393834 358568 393834 0 mprj/dcache_wb_o_dat\[10\]
rlabel metal2 336056 383894 336056 383894 0 mprj/dcache_wb_o_dat\[11\]
rlabel metal2 401464 388528 401464 388528 0 mprj/dcache_wb_o_dat\[12\]
rlabel metal2 357560 383782 357560 383782 0 mprj/dcache_wb_o_dat\[13\]
rlabel metal2 368312 384062 368312 384062 0 mprj/dcache_wb_o_dat\[14\]
rlabel metal3 380240 386120 380240 386120 0 mprj/dcache_wb_o_dat\[15\]
rlabel metal2 136808 393890 136808 393890 0 mprj/dcache_wb_o_dat\[1\]
rlabel metal2 165032 393330 165032 393330 0 mprj/dcache_wb_o_dat\[2\]
rlabel metal2 189224 393666 189224 393666 0 mprj/dcache_wb_o_dat\[3\]
rlabel metal2 213416 390418 213416 390418 0 mprj/dcache_wb_o_dat\[4\]
rlabel metal2 237608 393834 237608 393834 0 mprj/dcache_wb_o_dat\[5\]
rlabel metal2 261800 392154 261800 392154 0 mprj/dcache_wb_o_dat\[6\]
rlabel metal2 285992 390754 285992 390754 0 mprj/dcache_wb_o_dat\[7\]
rlabel metal3 306992 389704 306992 389704 0 mprj/dcache_wb_o_dat\[8\]
rlabel metal2 334376 393778 334376 393778 0 mprj/dcache_wb_o_dat\[9\]
rlabel metal2 214200 383950 214200 383950 0 mprj/dcache_wb_sel\[0\]
rlabel metal2 140840 393834 140840 393834 0 mprj/dcache_wb_sel\[1\]
rlabel metal2 72296 393666 72296 393666 0 mprj/dcache_wb_stb
rlabel metal2 76328 390418 76328 390418 0 mprj/dcache_wb_we
rlabel metal2 170968 77462 170968 77462 0 mprj/ic0_clk
rlabel metal4 170520 202104 170520 202104 0 mprj/ic0_mem_ack
rlabel metal4 172200 202944 172200 202944 0 mprj/ic0_mem_addr\[0\]
rlabel metal4 169064 285600 169064 285600 0 mprj/ic0_mem_addr\[10\]
rlabel metal4 170856 294112 170856 294112 0 mprj/ic0_mem_addr\[11\]
rlabel metal4 172536 302624 172536 302624 0 mprj/ic0_mem_addr\[12\]
rlabel metal3 169400 289016 169400 289016 0 mprj/ic0_mem_addr\[13\]
rlabel metal4 169288 319648 169288 319648 0 mprj/ic0_mem_addr\[14\]
rlabel metal4 172648 328160 172648 328160 0 mprj/ic0_mem_addr\[15\]
rlabel metal4 172312 207984 172312 207984 0 mprj/ic0_mem_addr\[1\]
rlabel metal3 173600 327320 173600 327320 0 mprj/ic0_mem_addr\[2\]
rlabel metal4 167272 226016 167272 226016 0 mprj/ic0_mem_addr\[3\]
rlabel metal4 170520 326592 170520 326592 0 mprj/ic0_mem_addr\[4\]
rlabel metal4 169848 332976 169848 332976 0 mprj/ic0_mem_addr\[5\]
rlabel metal3 152894 164584 152894 164584 0 mprj/ic0_mem_addr\[6\]
rlabel metal3 152950 178920 152950 178920 0 mprj/ic0_mem_addr\[7\]
rlabel metal3 153006 193256 153006 193256 0 mprj/ic0_mem_addr\[8\]
rlabel metal3 161966 207592 161966 207592 0 mprj/ic0_mem_addr\[9\]
rlabel metal4 170968 239400 170968 239400 0 mprj/ic0_mem_cache_flush
rlabel metal4 169960 318416 169960 318416 0 mprj/ic0_mem_data\[0\]
rlabel metal4 169176 287728 169176 287728 0 mprj/ic0_mem_data\[10\]
rlabel metal4 171304 351036 171304 351036 0 mprj/ic0_mem_data\[11\]
rlabel metal4 169848 354480 169848 354480 0 mprj/ic0_mem_data\[12\]
rlabel metal3 173656 357560 173656 357560 0 mprj/ic0_mem_data\[13\]
rlabel metal3 168952 355096 168952 355096 0 mprj/ic0_mem_data\[14\]
rlabel metal3 167384 334376 167384 334376 0 mprj/ic0_mem_data\[15\]
rlabel metal4 170856 362880 170856 362880 0 mprj/ic0_mem_data\[16\]
rlabel metal3 153902 311528 153902 311528 0 mprj/ic0_mem_data\[17\]
rlabel metal3 152558 315112 152558 315112 0 mprj/ic0_mem_data\[18\]
rlabel metal3 153398 318696 153398 318696 0 mprj/ic0_mem_data\[19\]
rlabel metal4 169848 321776 169848 321776 0 mprj/ic0_mem_data\[1\]
rlabel metal3 152670 322280 152670 322280 0 mprj/ic0_mem_data\[20\]
rlabel metal3 152782 325864 152782 325864 0 mprj/ic0_mem_data\[21\]
rlabel metal3 152502 329448 152502 329448 0 mprj/ic0_mem_data\[22\]
rlabel metal4 169848 368592 169848 368592 0 mprj/ic0_mem_data\[23\]
rlabel metal3 155190 336616 155190 336616 0 mprj/ic0_mem_data\[24\]
rlabel metal3 153566 340200 153566 340200 0 mprj/ic0_mem_data\[25\]
rlabel metal4 168840 357952 168840 357952 0 mprj/ic0_mem_data\[26\]
rlabel metal3 151830 347368 151830 347368 0 mprj/ic0_mem_data\[27\]
rlabel metal3 152222 350952 152222 350952 0 mprj/ic0_mem_data\[28\]
rlabel metal3 152166 354536 152166 354536 0 mprj/ic0_mem_data\[29\]
rlabel metal4 169848 326872 169848 326872 0 mprj/ic0_mem_data\[2\]
rlabel metal3 151886 358120 151886 358120 0 mprj/ic0_mem_data\[30\]
rlabel metal4 165480 368592 165480 368592 0 mprj/ic0_mem_data\[31\]
rlabel metal3 153622 125160 153622 125160 0 mprj/ic0_mem_data\[3\]
rlabel metal3 153678 139496 153678 139496 0 mprj/ic0_mem_data\[4\]
rlabel metal3 165802 336504 165802 336504 0 mprj/ic0_mem_data\[5\]
rlabel metal3 153790 168168 153790 168168 0 mprj/ic0_mem_data\[6\]
rlabel metal3 150486 182504 150486 182504 0 mprj/ic0_mem_data\[7\]
rlabel metal4 172424 270704 172424 270704 0 mprj/ic0_mem_data\[8\]
rlabel metal3 161854 211176 161854 211176 0 mprj/ic0_mem_data\[9\]
rlabel metal4 170744 220416 170744 220416 0 mprj/ic0_mem_ppl_submit
rlabel metal4 169848 315672 169848 315672 0 mprj/ic0_mem_req
rlabel metal4 168840 196168 168840 196168 0 mprj/ic0_rst
rlabel metal4 167160 196224 167160 196224 0 mprj/ic0_wb_ack
rlabel metal3 151886 78568 151886 78568 0 mprj/ic0_wb_adr\[0\]
rlabel metal4 170968 345464 170968 345464 0 mprj/ic0_wb_adr\[10\]
rlabel metal3 154294 243432 154294 243432 0 mprj/ic0_wb_adr\[11\]
rlabel metal3 154238 257768 154238 257768 0 mprj/ic0_wb_adr\[12\]
rlabel metal3 165914 358680 165914 358680 0 mprj/ic0_wb_adr\[13\]
rlabel metal3 155582 286440 155582 286440 0 mprj/ic0_wb_adr\[14\]
rlabel metal4 169848 363104 169848 363104 0 mprj/ic0_wb_adr\[15\]
rlabel metal3 151438 96488 151438 96488 0 mprj/ic0_wb_adr\[1\]
rlabel metal3 155302 114408 155302 114408 0 mprj/ic0_wb_adr\[2\]
rlabel metal3 166474 331800 166474 331800 0 mprj/ic0_wb_adr\[3\]
rlabel metal3 155358 143080 155358 143080 0 mprj/ic0_wb_adr\[4\]
rlabel metal3 162022 157416 162022 157416 0 mprj/ic0_wb_adr\[5\]
rlabel metal3 155414 171752 155414 171752 0 mprj/ic0_wb_adr\[6\]
rlabel metal3 167440 329224 167440 329224 0 mprj/ic0_wb_adr\[7\]
rlabel metal3 155526 200424 155526 200424 0 mprj/ic0_wb_adr\[8\]
rlabel metal4 165704 281344 165704 281344 0 mprj/ic0_wb_adr\[9\]
rlabel metal3 152054 57064 152054 57064 0 mprj/ic0_wb_cyc
rlabel metal4 171192 311136 171192 311136 0 mprj/ic0_wb_err
rlabel metal3 155190 82152 155190 82152 0 mprj/ic0_wb_i_dat\[0\]
rlabel metal3 166152 351064 166152 351064 0 mprj/ic0_wb_i_dat\[10\]
rlabel metal3 165130 353976 165130 353976 0 mprj/ic0_wb_i_dat\[11\]
rlabel metal4 169400 330792 169400 330792 0 mprj/ic0_wb_i_dat\[12\]
rlabel metal4 166152 317520 166152 317520 0 mprj/ic0_wb_i_dat\[13\]
rlabel metal4 167496 326032 167496 326032 0 mprj/ic0_wb_i_dat\[14\]
rlabel metal3 151942 304360 151942 304360 0 mprj/ic0_wb_i_dat\[15\]
rlabel metal3 151886 100072 151886 100072 0 mprj/ic0_wb_i_dat\[1\]
rlabel metal4 168952 226632 168952 226632 0 mprj/ic0_wb_i_dat\[2\]
rlabel metal3 164066 332472 164066 332472 0 mprj/ic0_wb_i_dat\[3\]
rlabel metal4 167384 247800 167384 247800 0 mprj/ic0_wb_i_dat\[4\]
rlabel metal3 152054 161000 152054 161000 0 mprj/ic0_wb_i_dat\[5\]
rlabel metal4 165592 257936 165592 257936 0 mprj/ic0_wb_i_dat\[6\]
rlabel metal3 152110 189672 152110 189672 0 mprj/ic0_wb_i_dat\[7\]
rlabel metal4 170632 274960 170632 274960 0 mprj/ic0_wb_i_dat\[8\]
rlabel metal3 152166 218344 152166 218344 0 mprj/ic0_wb_i_dat\[9\]
rlabel metal3 151830 85736 151830 85736 0 mprj/ic0_wb_sel\[0\]
rlabel metal4 162456 215376 162456 215376 0 mprj/ic0_wb_sel\[1\]
rlabel metal4 162008 292600 162008 292600 0 mprj/ic0_wb_stb
rlabel metal4 165480 194152 165480 194152 0 mprj/ic0_wb_we
rlabel metal2 220696 78302 220696 78302 0 mprj/ic1_clk
rlabel metal3 436520 45304 436520 45304 0 mprj/ic1_mem_ack
rlabel metal3 441098 71400 441098 71400 0 mprj/ic1_mem_addr\[0\]
rlabel metal4 426440 285600 426440 285600 0 mprj/ic1_mem_addr\[10\]
rlabel metal4 427896 294112 427896 294112 0 mprj/ic1_mem_addr\[11\]
rlabel metal3 423598 354648 423598 354648 0 mprj/ic1_mem_addr\[12\]
rlabel metal4 431256 311136 431256 311136 0 mprj/ic1_mem_addr\[13\]
rlabel metal3 439530 279272 439530 279272 0 mprj/ic1_mem_addr\[14\]
rlabel metal3 441266 293608 441266 293608 0 mprj/ic1_mem_addr\[15\]
rlabel metal4 425992 206864 425992 206864 0 mprj/ic1_mem_addr\[1\]
rlabel metal4 427672 217504 427672 217504 0 mprj/ic1_mem_addr\[2\]
rlabel metal3 440314 121576 440314 121576 0 mprj/ic1_mem_addr\[3\]
rlabel metal3 424326 333144 424326 333144 0 mprj/ic1_mem_addr\[4\]
rlabel metal4 431032 243040 431032 243040 0 mprj/ic1_mem_addr\[5\]
rlabel metal3 438578 164584 438578 164584 0 mprj/ic1_mem_addr\[6\]
rlabel metal4 424312 260064 424312 260064 0 mprj/ic1_mem_addr\[7\]
rlabel metal4 427784 268576 427784 268576 0 mprj/ic1_mem_addr\[8\]
rlabel metal4 426328 277088 426328 277088 0 mprj/ic1_mem_addr\[9\]
rlabel metal4 430920 182280 430920 182280 0 mprj/ic1_mem_cache_flush
rlabel metal3 442274 74984 442274 74984 0 mprj/ic1_mem_data\[0\]
rlabel metal3 426454 349944 426454 349944 0 mprj/ic1_mem_data\[10\]
rlabel metal4 429240 296240 429240 296240 0 mprj/ic1_mem_data\[11\]
rlabel metal3 425278 355320 425278 355320 0 mprj/ic1_mem_data\[12\]
rlabel metal3 416822 358008 416822 358008 0 mprj/ic1_mem_data\[13\]
rlabel metal3 416878 360696 416878 360696 0 mprj/ic1_mem_data\[14\]
rlabel metal3 440762 297192 440762 297192 0 mprj/ic1_mem_data\[15\]
rlabel metal3 432026 307944 432026 307944 0 mprj/ic1_mem_data\[16\]
rlabel metal3 431578 311528 431578 311528 0 mprj/ic1_mem_data\[17\]
rlabel metal3 437080 334376 437080 334376 0 mprj/ic1_mem_data\[18\]
rlabel metal4 429464 343784 429464 343784 0 mprj/ic1_mem_data\[19\]
rlabel metal3 431690 92904 431690 92904 0 mprj/ic1_mem_data\[1\]
rlabel metal3 442554 322280 442554 322280 0 mprj/ic1_mem_data\[20\]
rlabel metal3 416150 368760 416150 368760 0 mprj/ic1_mem_data\[21\]
rlabel metal4 428008 354872 428008 354872 0 mprj/ic1_mem_data\[22\]
rlabel metal4 425992 355992 425992 355992 0 mprj/ic1_mem_data\[23\]
rlabel metal4 421064 365568 421064 365568 0 mprj/ic1_mem_data\[24\]
rlabel metal3 415926 371448 415926 371448 0 mprj/ic1_mem_data\[25\]
rlabel metal3 429520 353640 429520 353640 0 mprj/ic1_mem_data\[26\]
rlabel metal3 438522 347368 438522 347368 0 mprj/ic1_mem_data\[27\]
rlabel metal3 415758 373464 415758 373464 0 mprj/ic1_mem_data\[28\]
rlabel metal4 422632 365568 422632 365568 0 mprj/ic1_mem_data\[29\]
rlabel metal3 416654 328440 416654 328440 0 mprj/ic1_mem_data\[2\]
rlabel metal4 420952 366464 420952 366464 0 mprj/ic1_mem_data\[30\]
rlabel metal3 413784 375354 413784 375354 0 mprj/ic1_mem_data\[31\]
rlabel metal3 439362 125160 439362 125160 0 mprj/ic1_mem_data\[3\]
rlabel metal3 416710 333816 416710 333816 0 mprj/ic1_mem_data\[4\]
rlabel metal3 423430 336504 423430 336504 0 mprj/ic1_mem_data\[5\]
rlabel metal4 426216 253680 426216 253680 0 mprj/ic1_mem_data\[6\]
rlabel metal3 415310 341880 415310 341880 0 mprj/ic1_mem_data\[7\]
rlabel metal4 424424 270704 424424 270704 0 mprj/ic1_mem_data\[8\]
rlabel metal3 441154 211176 441154 211176 0 mprj/ic1_mem_data\[9\]
rlabel metal4 420952 199472 420952 199472 0 mprj/ic1_mem_ppl_submit
rlabel metal3 442666 49896 442666 49896 0 mprj/ic1_mem_req
rlabel metal5 428400 75510 428400 75510 0 mprj/ic1_rst
rlabel metal4 420840 201376 420840 201376 0 mprj/ic1_wb_ack
rlabel metal3 442778 78568 442778 78568 0 mprj/ic1_wb_adr\[0\]
rlabel metal3 416094 350616 416094 350616 0 mprj/ic1_wb_adr\[10\]
rlabel metal4 429352 294392 429352 294392 0 mprj/ic1_wb_adr\[11\]
rlabel metal4 421624 306880 421624 306880 0 mprj/ic1_wb_adr\[12\]
rlabel metal3 428246 358680 428246 358680 0 mprj/ic1_wb_adr\[13\]
rlabel metal4 420728 323904 420728 323904 0 mprj/ic1_wb_adr\[14\]
rlabel metal4 420840 347984 420840 347984 0 mprj/ic1_wb_adr\[15\]
rlabel metal4 421064 211120 421064 211120 0 mprj/ic1_wb_adr\[1\]
rlabel metal4 424536 311976 424536 311976 0 mprj/ic1_wb_adr\[2\]
rlabel metal4 421288 230272 421288 230272 0 mprj/ic1_wb_adr\[3\]
rlabel metal4 421400 238784 421400 238784 0 mprj/ic1_wb_adr\[4\]
rlabel metal4 421512 255528 421512 255528 0 mprj/ic1_wb_adr\[5\]
rlabel metal3 442778 171752 442778 171752 0 mprj/ic1_wb_adr\[6\]
rlabel metal3 442834 186088 442834 186088 0 mprj/ic1_wb_adr\[7\]
rlabel metal4 431144 261968 431144 261968 0 mprj/ic1_wb_adr\[8\]
rlabel metal3 438634 214760 438634 214760 0 mprj/ic1_wb_adr\[9\]
rlabel metal4 426104 202440 426104 202440 0 mprj/ic1_wb_cyc
rlabel metal4 429464 311136 429464 311136 0 mprj/ic1_wb_err
rlabel metal4 421176 190456 421176 190456 0 mprj/ic1_wb_i_dat\[0\]
rlabel metal4 420952 344064 420952 344064 0 mprj/ic1_wb_i_dat\[10\]
rlabel metal3 414862 353976 414862 353976 0 mprj/ic1_wb_i_dat\[11\]
rlabel metal3 415870 356664 415870 356664 0 mprj/ic1_wb_i_dat\[12\]
rlabel metal4 424648 288792 424648 288792 0 mprj/ic1_wb_i_dat\[13\]
rlabel metal4 422520 346080 422520 346080 0 mprj/ic1_wb_i_dat\[14\]
rlabel metal3 430122 304360 430122 304360 0 mprj/ic1_wb_i_dat\[15\]
rlabel metal4 422856 215712 422856 215712 0 mprj/ic1_wb_i_dat\[1\]
rlabel metal4 422744 224952 422744 224952 0 mprj/ic1_wb_i_dat\[2\]
rlabel metal4 422968 232400 422968 232400 0 mprj/ic1_wb_i_dat\[3\]
rlabel metal3 442946 146664 442946 146664 0 mprj/ic1_wb_i_dat\[4\]
rlabel metal4 423080 249424 423080 249424 0 mprj/ic1_wb_i_dat\[5\]
rlabel metal4 423192 257936 423192 257936 0 mprj/ic1_wb_i_dat\[6\]
rlabel metal4 423304 266448 423304 266448 0 mprj/ic1_wb_i_dat\[7\]
rlabel metal3 415814 345912 415814 345912 0 mprj/ic1_wb_i_dat\[8\]
rlabel metal3 442890 218344 442890 218344 0 mprj/ic1_wb_i_dat\[9\]
rlabel metal3 415310 323736 415310 323736 0 mprj/ic1_wb_sel\[0\]
rlabel metal4 422632 215376 422632 215376 0 mprj/ic1_wb_sel\[1\]
rlabel metal3 442666 64232 442666 64232 0 mprj/ic1_wb_stb
rlabel metal4 422520 199360 422520 199360 0 mprj/ic1_wb_we
rlabel metal2 172312 187334 172312 187334 0 mprj/inner_clock
rlabel metal2 172984 77462 172984 77462 0 mprj/inner_disable
rlabel metal3 223776 93352 223776 93352 0 mprj/inner_embed_mode
rlabel metal2 273112 306530 273112 306530 0 mprj/inner_ext_irq
rlabel metal3 226128 100184 226128 100184 0 mprj/inner_reset
rlabel metal3 225400 94920 225400 94920 0 mprj/inner_wb_4_burst
rlabel metal2 274008 306642 274008 306642 0 mprj/inner_wb_8_burst
rlabel metal2 177016 79534 177016 79534 0 mprj/inner_wb_ack
rlabel metal2 180376 79590 180376 79590 0 mprj/inner_wb_adr\[0\]
rlabel metal2 201880 79646 201880 79646 0 mprj/inner_wb_adr\[10\]
rlabel metal3 248136 100408 248136 100408 0 mprj/inner_wb_adr\[11\]
rlabel metal3 249816 98840 249816 98840 0 mprj/inner_wb_adr\[12\]
rlabel metal3 251496 93576 251496 93576 0 mprj/inner_wb_adr\[13\]
rlabel metal2 209944 86478 209944 86478 0 mprj/inner_wb_adr\[14\]
rlabel metal2 211960 80374 211960 80374 0 mprj/inner_wb_adr\[15\]
rlabel metal4 213976 82817 213976 82817 0 mprj/inner_wb_adr\[16\]
rlabel metal2 214774 75880 214774 75880 0 mprj/inner_wb_adr\[17\]
rlabel metal2 215320 80430 215320 80430 0 mprj/inner_wb_adr\[18\]
rlabel metal2 215992 80486 215992 80486 0 mprj/inner_wb_adr\[19\]
rlabel metal3 230776 101864 230776 101864 0 mprj/inner_wb_adr\[1\]
rlabel metal2 216664 79758 216664 79758 0 mprj/inner_wb_adr\[20\]
rlabel metal2 217336 78022 217336 78022 0 mprj/inner_wb_adr\[21\]
rlabel metal2 218008 79702 218008 79702 0 mprj/inner_wb_adr\[22\]
rlabel metal2 218680 88662 218680 88662 0 mprj/inner_wb_adr\[23\]
rlabel metal2 185752 87150 185752 87150 0 mprj/inner_wb_adr\[2\]
rlabel metal2 187768 81214 187768 81214 0 mprj/inner_wb_adr\[3\]
rlabel metal2 189658 75880 189658 75880 0 mprj/inner_wb_adr\[4\]
rlabel metal2 191800 81270 191800 81270 0 mprj/inner_wb_adr\[5\]
rlabel metal3 285208 305256 285208 305256 0 mprj/inner_wb_adr\[6\]
rlabel metal3 285040 305368 285040 305368 0 mprj/inner_wb_adr\[7\]
rlabel metal2 288344 194810 288344 194810 0 mprj/inner_wb_adr\[8\]
rlabel metal2 289688 204778 289688 204778 0 mprj/inner_wb_adr\[9\]
rlabel metal3 227752 98504 227752 98504 0 mprj/inner_wb_cyc
rlabel metal3 226856 101640 226856 101640 0 mprj/inner_wb_err
rlabel metal3 229096 101752 229096 101752 0 mprj/inner_wb_i_dat\[0\]
rlabel metal3 291088 305256 291088 305256 0 mprj/inner_wb_i_dat\[10\]
rlabel metal2 204750 75880 204750 75880 0 mprj/inner_wb_i_dat\[11\]
rlabel metal2 294168 306642 294168 306642 0 mprj/inner_wb_i_dat\[12\]
rlabel metal3 212688 80472 212688 80472 0 mprj/inner_wb_i_dat\[13\]
rlabel metal2 210616 82110 210616 82110 0 mprj/inner_wb_i_dat\[14\]
rlabel metal2 212632 81382 212632 81382 0 mprj/inner_wb_i_dat\[15\]
rlabel metal2 278936 201586 278936 201586 0 mprj/inner_wb_i_dat\[1\]
rlabel metal2 186424 82894 186424 82894 0 mprj/inner_wb_i_dat\[2\]
rlabel metal2 188440 87262 188440 87262 0 mprj/inner_wb_i_dat\[3\]
rlabel metal3 191576 80584 191576 80584 0 mprj/inner_wb_i_dat\[4\]
rlabel metal3 285264 305480 285264 305480 0 mprj/inner_wb_i_dat\[5\]
rlabel metal2 194488 77070 194488 77070 0 mprj/inner_wb_i_dat\[6\]
rlabel metal2 196504 77462 196504 77462 0 mprj/inner_wb_i_dat\[7\]
rlabel metal2 288792 199066 288792 199066 0 mprj/inner_wb_i_dat\[8\]
rlabel metal2 290136 203378 290136 203378 0 mprj/inner_wb_i_dat\[9\]
rlabel metal3 227360 93464 227360 93464 0 mprj/inner_wb_o_dat\[0\]
rlabel metal2 203224 83118 203224 83118 0 mprj/inner_wb_o_dat\[10\]
rlabel metal2 205240 83174 205240 83174 0 mprj/inner_wb_o_dat\[11\]
rlabel metal2 207256 83230 207256 83230 0 mprj/inner_wb_o_dat\[12\]
rlabel metal2 209272 84798 209272 84798 0 mprj/inner_wb_o_dat\[13\]
rlabel metal2 211288 85582 211288 85582 0 mprj/inner_wb_o_dat\[14\]
rlabel metal2 213304 78806 213304 78806 0 mprj/inner_wb_o_dat\[15\]
rlabel metal2 279384 199906 279384 199906 0 mprj/inner_wb_o_dat\[1\]
rlabel metal2 281176 306194 281176 306194 0 mprj/inner_wb_o_dat\[2\]
rlabel metal2 282520 306474 282520 306474 0 mprj/inner_wb_o_dat\[3\]
rlabel metal3 282632 305144 282632 305144 0 mprj/inner_wb_o_dat\[4\]
rlabel metal3 194432 80584 194432 80584 0 mprj/inner_wb_o_dat\[5\]
rlabel metal3 285768 305144 285768 305144 0 mprj/inner_wb_o_dat\[6\]
rlabel metal2 237720 83496 237720 83496 0 mprj/inner_wb_o_dat\[7\]
rlabel metal2 238616 85512 238616 85512 0 mprj/inner_wb_o_dat\[8\]
rlabel metal2 290584 200074 290584 200074 0 mprj/inner_wb_o_dat\[9\]
rlabel metal3 230216 91672 230216 91672 0 mprj/inner_wb_sel\[0\]
rlabel metal3 186200 80584 186200 80584 0 mprj/inner_wb_sel\[1\]
rlabel metal2 234360 90160 234360 90160 0 mprj/inner_wb_stb
rlabel metal3 227976 91560 227976 91560 0 mprj/inner_wb_we
rlabel metal3 267414 22344 267414 22344 0 mprj/iram_addr\[0\]
rlabel metal4 265944 24248 265944 24248 0 mprj/iram_addr\[1\]
rlabel metal3 267470 30408 267470 30408 0 mprj/iram_addr\[2\]
rlabel metal3 266070 34440 266070 34440 0 mprj/iram_addr\[3\]
rlabel metal4 270088 37352 270088 37352 0 mprj/iram_addr\[4\]
rlabel metal3 265944 42098 265944 42098 0 mprj/iram_addr\[5\]
rlabel metal3 268002 14280 268002 14280 0 mprj/iram_clk
rlabel metal3 267470 23688 267470 23688 0 mprj/iram_i_data\[0\]
rlabel metal3 265944 57526 265944 57526 0 mprj/iram_i_data\[10\]
rlabel metal3 265944 60326 265944 60326 0 mprj/iram_i_data\[11\]
rlabel metal3 265944 63014 265944 63014 0 mprj/iram_i_data\[12\]
rlabel metal3 268030 65352 268030 65352 0 mprj/iram_i_data\[13\]
rlabel metal3 265944 68278 265944 68278 0 mprj/iram_i_data\[14\]
rlabel metal4 268968 72296 268968 72296 0 mprj/iram_i_data\[15\]
rlabel metal3 268030 27720 268030 27720 0 mprj/iram_i_data\[1\]
rlabel metal4 265944 30072 265944 30072 0 mprj/iram_i_data\[2\]
rlabel metal3 265944 35658 265944 35658 0 mprj/iram_i_data\[3\]
rlabel metal4 268856 38808 268856 38808 0 mprj/iram_i_data\[4\]
rlabel metal3 265944 43498 265944 43498 0 mprj/iram_i_data\[5\]
rlabel metal3 265944 46298 265944 46298 0 mprj/iram_i_data\[6\]
rlabel metal3 265944 48986 265944 48986 0 mprj/iram_i_data\[7\]
rlabel metal3 268016 51912 268016 51912 0 mprj/iram_i_data\[8\]
rlabel metal3 265944 54838 265944 54838 0 mprj/iram_i_data\[9\]
rlabel metal3 266518 25032 266518 25032 0 mprj/iram_o_data\[0\]
rlabel metal3 265944 58982 265944 58982 0 mprj/iram_o_data\[10\]
rlabel metal3 265944 61726 265944 61726 0 mprj/iram_o_data\[11\]
rlabel metal4 265944 65016 265944 65016 0 mprj/iram_o_data\[12\]
rlabel metal3 269458 69160 269458 69160 0 mprj/iram_o_data\[13\]
rlabel metal4 265944 71008 265944 71008 0 mprj/iram_o_data\[14\]
rlabel metal3 267414 72072 267414 72072 0 mprj/iram_o_data\[15\]
rlabel metal3 267414 29064 267414 29064 0 mprj/iram_o_data\[1\]
rlabel metal3 269458 29960 269458 29960 0 mprj/iram_o_data\[2\]
rlabel metal4 265944 36120 265944 36120 0 mprj/iram_o_data\[3\]
rlabel metal3 265944 40810 265944 40810 0 mprj/iram_o_data\[4\]
rlabel metal3 265944 44898 265944 44898 0 mprj/iram_o_data\[5\]
rlabel metal3 265944 47698 265944 47698 0 mprj/iram_o_data\[6\]
rlabel metal3 265944 50442 265944 50442 0 mprj/iram_o_data\[7\]
rlabel metal3 265944 53382 265944 53382 0 mprj/iram_o_data\[8\]
rlabel metal3 265944 56294 265944 56294 0 mprj/iram_o_data\[9\]
rlabel metal3 268030 21000 268030 21000 0 mprj/iram_we
rlabel via4 210168 13397 210168 13397 0 user_clock2
rlabel metal4 209496 13217 209496 13217 0 user_irq[0]
rlabel metal4 169624 44925 169624 44925 0 user_irq[1]
rlabel metal4 209944 13307 209944 13307 0 user_irq[2]
rlabel metal3 185472 12264 185472 12264 0 wb_clk_i
rlabel metal3 185752 12488 185752 12488 0 wb_rst_i
rlabel metal2 15400 1470 15400 1470 0 wbs_ack_o
rlabel metal2 23016 2366 23016 2366 0 wbs_adr_i[0]
rlabel metal3 191576 13496 191576 13496 0 wbs_adr_i[10]
rlabel metal2 93464 2534 93464 2534 0 wbs_adr_i[11]
rlabel metal2 99064 1638 99064 1638 0 wbs_adr_i[12]
rlabel metal2 104664 7070 104664 7070 0 wbs_adr_i[13]
rlabel metal2 110600 1694 110600 1694 0 wbs_adr_i[14]
rlabel metal2 116312 3374 116312 3374 0 wbs_adr_i[15]
rlabel metal2 122024 3430 122024 3430 0 wbs_adr_i[16]
rlabel metal2 127624 3486 127624 3486 0 wbs_adr_i[17]
rlabel metal2 133224 7574 133224 7574 0 wbs_adr_i[18]
rlabel metal2 139160 1806 139160 1806 0 wbs_adr_i[19]
rlabel metal2 30632 3150 30632 3150 0 wbs_adr_i[1]
rlabel metal2 144648 7630 144648 7630 0 wbs_adr_i[20]
rlabel metal2 150584 1862 150584 1862 0 wbs_adr_i[21]
rlabel metal2 156184 2590 156184 2590 0 wbs_adr_i[22]
rlabel metal2 162008 1414 162008 1414 0 wbs_adr_i[23]
rlabel metal2 167496 7406 167496 7406 0 wbs_adr_i[24]
rlabel metal2 173432 4382 173432 4382 0 wbs_adr_i[25]
rlabel metal2 179144 3934 179144 3934 0 wbs_adr_i[26]
rlabel metal3 195440 8232 195440 8232 0 wbs_adr_i[27]
rlabel metal2 206808 13482 206808 13482 0 wbs_adr_i[28]
rlabel metal2 196280 4410 196280 4410 0 wbs_adr_i[29]
rlabel metal2 38360 280 38360 280 0 wbs_adr_i[2]
rlabel metal3 205072 10024 205072 10024 0 wbs_adr_i[30]
rlabel metal2 208824 14714 208824 14714 0 wbs_adr_i[31]
rlabel metal2 45976 336 45976 336 0 wbs_adr_i[3]
rlabel metal2 53256 6958 53256 6958 0 wbs_adr_i[4]
rlabel metal2 59304 392 59304 392 0 wbs_adr_i[5]
rlabel metal3 192024 448 192024 448 0 wbs_adr_i[6]
rlabel metal2 70504 3262 70504 3262 0 wbs_adr_i[7]
rlabel metal2 76328 462 76328 462 0 wbs_adr_i[8]
rlabel metal2 194040 11858 194040 11858 0 wbs_adr_i[9]
rlabel metal4 186200 10767 186200 10767 0 wbs_cyc_i
rlabel metal2 24920 4830 24920 4830 0 wbs_dat_i[0]
rlabel metal2 194936 12754 194936 12754 0 wbs_dat_i[10]
rlabel metal2 95368 1582 95368 1582 0 wbs_dat_i[11]
rlabel metal2 101080 518 101080 518 0 wbs_dat_i[12]
rlabel metal2 106568 7518 106568 7518 0 wbs_dat_i[13]
rlabel metal2 112504 5054 112504 5054 0 wbs_dat_i[14]
rlabel metal2 117992 7798 117992 7798 0 wbs_dat_i[15]
rlabel metal2 123928 1750 123928 1750 0 wbs_dat_i[16]
rlabel metal2 129640 5894 129640 5894 0 wbs_dat_i[17]
rlabel metal2 135352 5950 135352 5950 0 wbs_dat_i[18]
rlabel metal2 141064 5838 141064 5838 0 wbs_dat_i[19]
rlabel metal2 188216 13482 188216 13482 0 wbs_dat_i[1]
rlabel metal2 146776 4270 146776 4270 0 wbs_dat_i[20]
rlabel metal2 152488 5110 152488 5110 0 wbs_dat_i[21]
rlabel metal2 158200 6006 158200 6006 0 wbs_dat_i[22]
rlabel metal2 163912 3542 163912 3542 0 wbs_dat_i[23]
rlabel metal2 169624 5222 169624 5222 0 wbs_dat_i[24]
rlabel metal2 175336 6062 175336 6062 0 wbs_dat_i[25]
rlabel metal3 193368 5768 193368 5768 0 wbs_dat_i[26]
rlabel metal3 196560 4984 196560 4984 0 wbs_dat_i[27]
rlabel metal2 192472 2310 192472 2310 0 wbs_dat_i[28]
rlabel metal2 198184 2310 198184 2310 0 wbs_dat_i[29]
rlabel metal3 188664 12264 188664 12264 0 wbs_dat_i[2]
rlabel metal2 208376 12250 208376 12250 0 wbs_dat_i[30]
rlabel metal2 209272 4200 209272 4200 0 wbs_dat_i[31]
rlabel metal2 47768 5726 47768 5726 0 wbs_dat_i[3]
rlabel metal2 55384 2142 55384 2142 0 wbs_dat_i[4]
rlabel metal2 191576 12698 191576 12698 0 wbs_dat_i[5]
rlabel metal2 192248 11018 192248 11018 0 wbs_dat_i[6]
rlabel metal2 72520 3990 72520 3990 0 wbs_dat_i[7]
rlabel metal2 78232 5782 78232 5782 0 wbs_dat_i[8]
rlabel metal3 193312 12488 193312 12488 0 wbs_dat_i[9]
rlabel metal2 26824 1918 26824 1918 0 wbs_dat_o[0]
rlabel metal2 91560 4158 91560 4158 0 wbs_dat_o[10]
rlabel metal2 97272 4998 97272 4998 0 wbs_dat_o[11]
rlabel metal2 196504 8554 196504 8554 0 wbs_dat_o[12]
rlabel metal2 108696 4214 108696 4214 0 wbs_dat_o[13]
rlabel metal2 114296 8246 114296 8246 0 wbs_dat_o[14]
rlabel metal2 120120 3318 120120 3318 0 wbs_dat_o[15]
rlabel metal2 125832 630 125832 630 0 wbs_dat_o[16]
rlabel metal2 131544 4326 131544 4326 0 wbs_dat_o[17]
rlabel metal2 137032 8190 137032 8190 0 wbs_dat_o[18]
rlabel metal2 142856 7854 142856 7854 0 wbs_dat_o[19]
rlabel metal2 116760 9688 116760 9688 0 wbs_dat_o[1]
rlabel metal2 148456 8134 148456 8134 0 wbs_dat_o[20]
rlabel metal2 154168 6846 154168 6846 0 wbs_dat_o[21]
rlabel metal2 160104 5166 160104 5166 0 wbs_dat_o[22]
rlabel metal2 165592 6230 165592 6230 0 wbs_dat_o[23]
rlabel metal2 171528 5614 171528 5614 0 wbs_dat_o[24]
rlabel metal2 177240 4774 177240 4774 0 wbs_dat_o[25]
rlabel metal3 194432 4872 194432 4872 0 wbs_dat_o[26]
rlabel metal2 206584 12642 206584 12642 0 wbs_dat_o[27]
rlabel metal2 194152 6622 194152 6622 0 wbs_dat_o[28]
rlabel metal3 204008 9912 204008 9912 0 wbs_dat_o[29]
rlabel metal2 189336 15162 189336 15162 0 wbs_dat_o[2]
rlabel metal2 208600 14658 208600 14658 0 wbs_dat_o[30]
rlabel metal3 210280 4424 210280 4424 0 wbs_dat_o[31]
rlabel metal2 49672 5838 49672 5838 0 wbs_dat_o[3]
rlabel metal3 190232 12152 190232 12152 0 wbs_dat_o[4]
rlabel metal1 186200 12936 186200 12936 0 wbs_dat_o[5]
rlabel metal2 68712 2254 68712 2254 0 wbs_dat_o[6]
rlabel metal2 74200 6622 74200 6622 0 wbs_dat_o[7]
rlabel metal3 193144 12152 193144 12152 0 wbs_dat_o[8]
rlabel metal2 92344 10752 92344 10752 0 wbs_dat_o[9]
rlabel metal2 28728 2366 28728 2366 0 wbs_sel_i[0]
rlabel metal2 188664 14322 188664 14322 0 wbs_sel_i[1]
rlabel metal2 43960 2422 43960 2422 0 wbs_sel_i[2]
rlabel metal2 51576 3598 51576 3598 0 wbs_sel_i[3]
rlabel metal2 186648 10122 186648 10122 0 wbs_stb_i
rlabel metal2 21112 3990 21112 3990 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
