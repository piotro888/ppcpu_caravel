magic
tech sky130B
magscale 1 2
timestamp 1662742412
<< nwell >>
rect 1066 149317 149170 149883
rect 1066 148229 149170 148795
rect 1066 147141 149170 147707
rect 1066 146053 149170 146619
rect 1066 144965 149170 145531
rect 1066 143877 149170 144443
rect 1066 142789 149170 143355
rect 1066 141701 149170 142267
rect 1066 140613 149170 141179
rect 1066 139525 149170 140091
rect 1066 138437 149170 139003
rect 1066 137349 149170 137915
rect 1066 136261 149170 136827
rect 1066 135173 149170 135739
rect 1066 134085 149170 134651
rect 1066 132997 149170 133563
rect 1066 131909 149170 132475
rect 1066 130821 149170 131387
rect 1066 129733 149170 130299
rect 1066 128645 149170 129211
rect 1066 127557 149170 128123
rect 1066 126469 149170 127035
rect 1066 125381 149170 125947
rect 1066 124293 149170 124859
rect 1066 123205 149170 123771
rect 1066 122117 149170 122683
rect 1066 121029 149170 121595
rect 1066 119941 149170 120507
rect 1066 118853 149170 119419
rect 1066 117765 149170 118331
rect 1066 116677 149170 117243
rect 1066 115589 149170 116155
rect 1066 114501 149170 115067
rect 1066 113413 149170 113979
rect 1066 112325 149170 112891
rect 1066 111237 149170 111803
rect 1066 110149 149170 110715
rect 1066 109061 149170 109627
rect 1066 107973 149170 108539
rect 1066 106885 149170 107451
rect 1066 105797 149170 106363
rect 1066 104709 149170 105275
rect 1066 103621 149170 104187
rect 1066 102533 149170 103099
rect 1066 101445 149170 102011
rect 1066 100357 149170 100923
rect 1066 99269 149170 99835
rect 1066 98181 149170 98747
rect 1066 97093 149170 97659
rect 1066 96005 149170 96571
rect 1066 94917 149170 95483
rect 1066 93829 149170 94395
rect 1066 92741 149170 93307
rect 1066 91653 149170 92219
rect 1066 90565 149170 91131
rect 1066 89477 149170 90043
rect 1066 88389 149170 88955
rect 1066 87301 149170 87867
rect 1066 86213 149170 86779
rect 1066 85125 149170 85691
rect 1066 84037 149170 84603
rect 1066 82949 149170 83515
rect 1066 81861 149170 82427
rect 1066 80773 149170 81339
rect 1066 79685 149170 80251
rect 1066 78597 149170 79163
rect 1066 77509 149170 78075
rect 1066 76421 149170 76987
rect 1066 75333 149170 75899
rect 1066 74245 149170 74811
rect 1066 73157 149170 73723
rect 1066 72069 149170 72635
rect 1066 70981 149170 71547
rect 1066 69893 149170 70459
rect 1066 68805 149170 69371
rect 1066 67717 149170 68283
rect 1066 66629 149170 67195
rect 1066 65541 149170 66107
rect 1066 64453 149170 65019
rect 1066 63365 149170 63931
rect 1066 62277 149170 62843
rect 1066 61189 149170 61755
rect 1066 60101 149170 60667
rect 1066 59013 149170 59579
rect 1066 57925 149170 58491
rect 1066 56837 149170 57403
rect 1066 55749 149170 56315
rect 1066 54661 149170 55227
rect 1066 53573 149170 54139
rect 1066 52485 149170 53051
rect 1066 51397 149170 51963
rect 1066 50309 149170 50875
rect 1066 49221 149170 49787
rect 1066 48133 149170 48699
rect 1066 47045 149170 47611
rect 1066 45957 149170 46523
rect 1066 44869 149170 45435
rect 1066 43781 149170 44347
rect 1066 42693 149170 43259
rect 1066 41605 149170 42171
rect 1066 40517 149170 41083
rect 1066 39429 149170 39995
rect 1066 38341 149170 38907
rect 1066 37253 149170 37819
rect 1066 36165 149170 36731
rect 1066 35077 149170 35643
rect 1066 33989 149170 34555
rect 1066 32901 149170 33467
rect 1066 31813 149170 32379
rect 1066 30725 149170 31291
rect 1066 29637 149170 30203
rect 1066 28549 149170 29115
rect 1066 27461 149170 28027
rect 1066 26373 149170 26939
rect 1066 25285 149170 25851
rect 1066 24197 149170 24763
rect 1066 23109 149170 23675
rect 1066 22021 149170 22587
rect 1066 20933 149170 21499
rect 1066 19845 149170 20411
rect 1066 18757 149170 19323
rect 1066 17669 149170 18235
rect 1066 16581 149170 17147
rect 1066 15493 149170 16059
rect 1066 14405 149170 14971
rect 1066 13317 149170 13883
rect 1066 12229 149170 12795
rect 1066 11141 149170 11707
rect 1066 10053 149170 10619
rect 1066 8965 149170 9531
rect 1066 7877 149170 8443
rect 1066 6789 149170 7355
rect 1066 5701 149170 6267
rect 1066 4613 149170 5179
rect 1066 3525 149170 4091
rect 1066 2437 149170 3003
<< obsli1 >>
rect 1104 2159 149132 150161
<< obsm1 >>
rect 1104 1640 149132 150408
<< metal2 >>
rect 5262 151637 5318 152437
rect 6274 151637 6330 152437
rect 7286 151637 7342 152437
rect 8298 151637 8354 152437
rect 9310 151637 9366 152437
rect 10322 151637 10378 152437
rect 11334 151637 11390 152437
rect 12346 151637 12402 152437
rect 13358 151637 13414 152437
rect 14370 151637 14426 152437
rect 15382 151637 15438 152437
rect 16394 151637 16450 152437
rect 17406 151637 17462 152437
rect 18418 151637 18474 152437
rect 19430 151637 19486 152437
rect 20442 151637 20498 152437
rect 21454 151637 21510 152437
rect 22466 151637 22522 152437
rect 23478 151637 23534 152437
rect 24490 151637 24546 152437
rect 25502 151637 25558 152437
rect 26514 151637 26570 152437
rect 27526 151637 27582 152437
rect 28538 151637 28594 152437
rect 29550 151637 29606 152437
rect 30562 151637 30618 152437
rect 31574 151637 31630 152437
rect 32586 151637 32642 152437
rect 33598 151637 33654 152437
rect 34610 151637 34666 152437
rect 35622 151637 35678 152437
rect 36634 151637 36690 152437
rect 37646 151637 37702 152437
rect 38658 151637 38714 152437
rect 39670 151637 39726 152437
rect 40682 151637 40738 152437
rect 41694 151637 41750 152437
rect 42706 151637 42762 152437
rect 43718 151637 43774 152437
rect 44730 151637 44786 152437
rect 45742 151637 45798 152437
rect 46754 151637 46810 152437
rect 47766 151637 47822 152437
rect 48778 151637 48834 152437
rect 49790 151637 49846 152437
rect 50802 151637 50858 152437
rect 51814 151637 51870 152437
rect 52826 151637 52882 152437
rect 53838 151637 53894 152437
rect 54850 151637 54906 152437
rect 55862 151637 55918 152437
rect 56874 151637 56930 152437
rect 57886 151637 57942 152437
rect 58898 151637 58954 152437
rect 59910 151637 59966 152437
rect 60922 151637 60978 152437
rect 61934 151637 61990 152437
rect 62946 151637 63002 152437
rect 63958 151637 64014 152437
rect 64970 151637 65026 152437
rect 65982 151637 66038 152437
rect 66994 151637 67050 152437
rect 68006 151637 68062 152437
rect 69018 151637 69074 152437
rect 70030 151637 70086 152437
rect 71042 151637 71098 152437
rect 72054 151637 72110 152437
rect 73066 151637 73122 152437
rect 74078 151637 74134 152437
rect 75090 151637 75146 152437
rect 76102 151637 76158 152437
rect 77114 151637 77170 152437
rect 78126 151637 78182 152437
rect 79138 151637 79194 152437
rect 80150 151637 80206 152437
rect 81162 151637 81218 152437
rect 82174 151637 82230 152437
rect 83186 151637 83242 152437
rect 84198 151637 84254 152437
rect 85210 151637 85266 152437
rect 86222 151637 86278 152437
rect 87234 151637 87290 152437
rect 88246 151637 88302 152437
rect 89258 151637 89314 152437
rect 90270 151637 90326 152437
rect 91282 151637 91338 152437
rect 92294 151637 92350 152437
rect 93306 151637 93362 152437
rect 94318 151637 94374 152437
rect 95330 151637 95386 152437
rect 96342 151637 96398 152437
rect 97354 151637 97410 152437
rect 98366 151637 98422 152437
rect 99378 151637 99434 152437
rect 100390 151637 100446 152437
rect 101402 151637 101458 152437
rect 102414 151637 102470 152437
rect 103426 151637 103482 152437
rect 104438 151637 104494 152437
rect 105450 151637 105506 152437
rect 106462 151637 106518 152437
rect 107474 151637 107530 152437
rect 108486 151637 108542 152437
rect 109498 151637 109554 152437
rect 110510 151637 110566 152437
rect 111522 151637 111578 152437
rect 112534 151637 112590 152437
rect 113546 151637 113602 152437
rect 114558 151637 114614 152437
rect 115570 151637 115626 152437
rect 116582 151637 116638 152437
rect 117594 151637 117650 152437
rect 118606 151637 118662 152437
rect 119618 151637 119674 152437
rect 120630 151637 120686 152437
rect 121642 151637 121698 152437
rect 122654 151637 122710 152437
rect 123666 151637 123722 152437
rect 124678 151637 124734 152437
rect 125690 151637 125746 152437
rect 126702 151637 126758 152437
rect 127714 151637 127770 152437
rect 128726 151637 128782 152437
rect 129738 151637 129794 152437
rect 130750 151637 130806 152437
rect 131762 151637 131818 152437
rect 132774 151637 132830 152437
rect 133786 151637 133842 152437
rect 134798 151637 134854 152437
rect 135810 151637 135866 152437
rect 136822 151637 136878 152437
rect 137834 151637 137890 152437
rect 138846 151637 138902 152437
rect 139858 151637 139914 152437
rect 140870 151637 140926 152437
rect 141882 151637 141938 152437
rect 142894 151637 142950 152437
rect 143906 151637 143962 152437
rect 144918 151637 144974 152437
rect 3238 0 3294 800
rect 4250 0 4306 800
rect 5262 0 5318 800
rect 6274 0 6330 800
rect 7286 0 7342 800
rect 8298 0 8354 800
rect 9310 0 9366 800
rect 10322 0 10378 800
rect 11334 0 11390 800
rect 12346 0 12402 800
rect 13358 0 13414 800
rect 14370 0 14426 800
rect 15382 0 15438 800
rect 16394 0 16450 800
rect 17406 0 17462 800
rect 18418 0 18474 800
rect 19430 0 19486 800
rect 20442 0 20498 800
rect 21454 0 21510 800
rect 22466 0 22522 800
rect 23478 0 23534 800
rect 24490 0 24546 800
rect 25502 0 25558 800
rect 26514 0 26570 800
rect 27526 0 27582 800
rect 28538 0 28594 800
rect 29550 0 29606 800
rect 30562 0 30618 800
rect 31574 0 31630 800
rect 32586 0 32642 800
rect 33598 0 33654 800
rect 34610 0 34666 800
rect 35622 0 35678 800
rect 36634 0 36690 800
rect 37646 0 37702 800
rect 38658 0 38714 800
rect 39670 0 39726 800
rect 40682 0 40738 800
rect 41694 0 41750 800
rect 42706 0 42762 800
rect 43718 0 43774 800
rect 44730 0 44786 800
rect 45742 0 45798 800
rect 46754 0 46810 800
rect 47766 0 47822 800
rect 48778 0 48834 800
rect 49790 0 49846 800
rect 50802 0 50858 800
rect 51814 0 51870 800
rect 52826 0 52882 800
rect 53838 0 53894 800
rect 54850 0 54906 800
rect 55862 0 55918 800
rect 56874 0 56930 800
rect 57886 0 57942 800
rect 58898 0 58954 800
rect 59910 0 59966 800
rect 60922 0 60978 800
rect 61934 0 61990 800
rect 62946 0 63002 800
rect 63958 0 64014 800
rect 64970 0 65026 800
rect 65982 0 66038 800
rect 66994 0 67050 800
rect 68006 0 68062 800
rect 69018 0 69074 800
rect 70030 0 70086 800
rect 71042 0 71098 800
rect 72054 0 72110 800
rect 73066 0 73122 800
rect 74078 0 74134 800
rect 75090 0 75146 800
rect 76102 0 76158 800
rect 77114 0 77170 800
rect 78126 0 78182 800
rect 79138 0 79194 800
rect 80150 0 80206 800
rect 81162 0 81218 800
rect 82174 0 82230 800
rect 83186 0 83242 800
rect 84198 0 84254 800
rect 85210 0 85266 800
rect 86222 0 86278 800
rect 87234 0 87290 800
rect 88246 0 88302 800
rect 89258 0 89314 800
rect 90270 0 90326 800
rect 91282 0 91338 800
rect 92294 0 92350 800
rect 93306 0 93362 800
rect 94318 0 94374 800
rect 95330 0 95386 800
rect 96342 0 96398 800
rect 97354 0 97410 800
rect 98366 0 98422 800
rect 99378 0 99434 800
rect 100390 0 100446 800
rect 101402 0 101458 800
rect 102414 0 102470 800
rect 103426 0 103482 800
rect 104438 0 104494 800
rect 105450 0 105506 800
rect 106462 0 106518 800
rect 107474 0 107530 800
rect 108486 0 108542 800
rect 109498 0 109554 800
rect 110510 0 110566 800
rect 111522 0 111578 800
rect 112534 0 112590 800
rect 113546 0 113602 800
rect 114558 0 114614 800
rect 115570 0 115626 800
rect 116582 0 116638 800
rect 117594 0 117650 800
rect 118606 0 118662 800
rect 119618 0 119674 800
rect 120630 0 120686 800
rect 121642 0 121698 800
rect 122654 0 122710 800
rect 123666 0 123722 800
rect 124678 0 124734 800
rect 125690 0 125746 800
rect 126702 0 126758 800
rect 127714 0 127770 800
rect 128726 0 128782 800
rect 129738 0 129794 800
rect 130750 0 130806 800
rect 131762 0 131818 800
rect 132774 0 132830 800
rect 133786 0 133842 800
rect 134798 0 134854 800
rect 135810 0 135866 800
rect 136822 0 136878 800
rect 137834 0 137890 800
rect 138846 0 138902 800
rect 139858 0 139914 800
rect 140870 0 140926 800
rect 141882 0 141938 800
rect 142894 0 142950 800
rect 143906 0 143962 800
rect 144918 0 144974 800
rect 145930 0 145986 800
rect 146942 0 146998 800
<< obsm2 >>
rect 2228 151581 5206 151722
rect 5374 151581 6218 151722
rect 6386 151581 7230 151722
rect 7398 151581 8242 151722
rect 8410 151581 9254 151722
rect 9422 151581 10266 151722
rect 10434 151581 11278 151722
rect 11446 151581 12290 151722
rect 12458 151581 13302 151722
rect 13470 151581 14314 151722
rect 14482 151581 15326 151722
rect 15494 151581 16338 151722
rect 16506 151581 17350 151722
rect 17518 151581 18362 151722
rect 18530 151581 19374 151722
rect 19542 151581 20386 151722
rect 20554 151581 21398 151722
rect 21566 151581 22410 151722
rect 22578 151581 23422 151722
rect 23590 151581 24434 151722
rect 24602 151581 25446 151722
rect 25614 151581 26458 151722
rect 26626 151581 27470 151722
rect 27638 151581 28482 151722
rect 28650 151581 29494 151722
rect 29662 151581 30506 151722
rect 30674 151581 31518 151722
rect 31686 151581 32530 151722
rect 32698 151581 33542 151722
rect 33710 151581 34554 151722
rect 34722 151581 35566 151722
rect 35734 151581 36578 151722
rect 36746 151581 37590 151722
rect 37758 151581 38602 151722
rect 38770 151581 39614 151722
rect 39782 151581 40626 151722
rect 40794 151581 41638 151722
rect 41806 151581 42650 151722
rect 42818 151581 43662 151722
rect 43830 151581 44674 151722
rect 44842 151581 45686 151722
rect 45854 151581 46698 151722
rect 46866 151581 47710 151722
rect 47878 151581 48722 151722
rect 48890 151581 49734 151722
rect 49902 151581 50746 151722
rect 50914 151581 51758 151722
rect 51926 151581 52770 151722
rect 52938 151581 53782 151722
rect 53950 151581 54794 151722
rect 54962 151581 55806 151722
rect 55974 151581 56818 151722
rect 56986 151581 57830 151722
rect 57998 151581 58842 151722
rect 59010 151581 59854 151722
rect 60022 151581 60866 151722
rect 61034 151581 61878 151722
rect 62046 151581 62890 151722
rect 63058 151581 63902 151722
rect 64070 151581 64914 151722
rect 65082 151581 65926 151722
rect 66094 151581 66938 151722
rect 67106 151581 67950 151722
rect 68118 151581 68962 151722
rect 69130 151581 69974 151722
rect 70142 151581 70986 151722
rect 71154 151581 71998 151722
rect 72166 151581 73010 151722
rect 73178 151581 74022 151722
rect 74190 151581 75034 151722
rect 75202 151581 76046 151722
rect 76214 151581 77058 151722
rect 77226 151581 78070 151722
rect 78238 151581 79082 151722
rect 79250 151581 80094 151722
rect 80262 151581 81106 151722
rect 81274 151581 82118 151722
rect 82286 151581 83130 151722
rect 83298 151581 84142 151722
rect 84310 151581 85154 151722
rect 85322 151581 86166 151722
rect 86334 151581 87178 151722
rect 87346 151581 88190 151722
rect 88358 151581 89202 151722
rect 89370 151581 90214 151722
rect 90382 151581 91226 151722
rect 91394 151581 92238 151722
rect 92406 151581 93250 151722
rect 93418 151581 94262 151722
rect 94430 151581 95274 151722
rect 95442 151581 96286 151722
rect 96454 151581 97298 151722
rect 97466 151581 98310 151722
rect 98478 151581 99322 151722
rect 99490 151581 100334 151722
rect 100502 151581 101346 151722
rect 101514 151581 102358 151722
rect 102526 151581 103370 151722
rect 103538 151581 104382 151722
rect 104550 151581 105394 151722
rect 105562 151581 106406 151722
rect 106574 151581 107418 151722
rect 107586 151581 108430 151722
rect 108598 151581 109442 151722
rect 109610 151581 110454 151722
rect 110622 151581 111466 151722
rect 111634 151581 112478 151722
rect 112646 151581 113490 151722
rect 113658 151581 114502 151722
rect 114670 151581 115514 151722
rect 115682 151581 116526 151722
rect 116694 151581 117538 151722
rect 117706 151581 118550 151722
rect 118718 151581 119562 151722
rect 119730 151581 120574 151722
rect 120742 151581 121586 151722
rect 121754 151581 122598 151722
rect 122766 151581 123610 151722
rect 123778 151581 124622 151722
rect 124790 151581 125634 151722
rect 125802 151581 126646 151722
rect 126814 151581 127658 151722
rect 127826 151581 128670 151722
rect 128838 151581 129682 151722
rect 129850 151581 130694 151722
rect 130862 151581 131706 151722
rect 131874 151581 132718 151722
rect 132886 151581 133730 151722
rect 133898 151581 134742 151722
rect 134910 151581 135754 151722
rect 135922 151581 136766 151722
rect 136934 151581 137778 151722
rect 137946 151581 138790 151722
rect 138958 151581 139802 151722
rect 139970 151581 140814 151722
rect 140982 151581 141826 151722
rect 141994 151581 142838 151722
rect 143006 151581 143850 151722
rect 144018 151581 144862 151722
rect 145030 151581 148470 151722
rect 2228 856 148470 151581
rect 2228 734 3182 856
rect 3350 734 4194 856
rect 4362 734 5206 856
rect 5374 734 6218 856
rect 6386 734 7230 856
rect 7398 734 8242 856
rect 8410 734 9254 856
rect 9422 734 10266 856
rect 10434 734 11278 856
rect 11446 734 12290 856
rect 12458 734 13302 856
rect 13470 734 14314 856
rect 14482 734 15326 856
rect 15494 734 16338 856
rect 16506 734 17350 856
rect 17518 734 18362 856
rect 18530 734 19374 856
rect 19542 734 20386 856
rect 20554 734 21398 856
rect 21566 734 22410 856
rect 22578 734 23422 856
rect 23590 734 24434 856
rect 24602 734 25446 856
rect 25614 734 26458 856
rect 26626 734 27470 856
rect 27638 734 28482 856
rect 28650 734 29494 856
rect 29662 734 30506 856
rect 30674 734 31518 856
rect 31686 734 32530 856
rect 32698 734 33542 856
rect 33710 734 34554 856
rect 34722 734 35566 856
rect 35734 734 36578 856
rect 36746 734 37590 856
rect 37758 734 38602 856
rect 38770 734 39614 856
rect 39782 734 40626 856
rect 40794 734 41638 856
rect 41806 734 42650 856
rect 42818 734 43662 856
rect 43830 734 44674 856
rect 44842 734 45686 856
rect 45854 734 46698 856
rect 46866 734 47710 856
rect 47878 734 48722 856
rect 48890 734 49734 856
rect 49902 734 50746 856
rect 50914 734 51758 856
rect 51926 734 52770 856
rect 52938 734 53782 856
rect 53950 734 54794 856
rect 54962 734 55806 856
rect 55974 734 56818 856
rect 56986 734 57830 856
rect 57998 734 58842 856
rect 59010 734 59854 856
rect 60022 734 60866 856
rect 61034 734 61878 856
rect 62046 734 62890 856
rect 63058 734 63902 856
rect 64070 734 64914 856
rect 65082 734 65926 856
rect 66094 734 66938 856
rect 67106 734 67950 856
rect 68118 734 68962 856
rect 69130 734 69974 856
rect 70142 734 70986 856
rect 71154 734 71998 856
rect 72166 734 73010 856
rect 73178 734 74022 856
rect 74190 734 75034 856
rect 75202 734 76046 856
rect 76214 734 77058 856
rect 77226 734 78070 856
rect 78238 734 79082 856
rect 79250 734 80094 856
rect 80262 734 81106 856
rect 81274 734 82118 856
rect 82286 734 83130 856
rect 83298 734 84142 856
rect 84310 734 85154 856
rect 85322 734 86166 856
rect 86334 734 87178 856
rect 87346 734 88190 856
rect 88358 734 89202 856
rect 89370 734 90214 856
rect 90382 734 91226 856
rect 91394 734 92238 856
rect 92406 734 93250 856
rect 93418 734 94262 856
rect 94430 734 95274 856
rect 95442 734 96286 856
rect 96454 734 97298 856
rect 97466 734 98310 856
rect 98478 734 99322 856
rect 99490 734 100334 856
rect 100502 734 101346 856
rect 101514 734 102358 856
rect 102526 734 103370 856
rect 103538 734 104382 856
rect 104550 734 105394 856
rect 105562 734 106406 856
rect 106574 734 107418 856
rect 107586 734 108430 856
rect 108598 734 109442 856
rect 109610 734 110454 856
rect 110622 734 111466 856
rect 111634 734 112478 856
rect 112646 734 113490 856
rect 113658 734 114502 856
rect 114670 734 115514 856
rect 115682 734 116526 856
rect 116694 734 117538 856
rect 117706 734 118550 856
rect 118718 734 119562 856
rect 119730 734 120574 856
rect 120742 734 121586 856
rect 121754 734 122598 856
rect 122766 734 123610 856
rect 123778 734 124622 856
rect 124790 734 125634 856
rect 125802 734 126646 856
rect 126814 734 127658 856
rect 127826 734 128670 856
rect 128838 734 129682 856
rect 129850 734 130694 856
rect 130862 734 131706 856
rect 131874 734 132718 856
rect 132886 734 133730 856
rect 133898 734 134742 856
rect 134910 734 135754 856
rect 135922 734 136766 856
rect 136934 734 137778 856
rect 137946 734 138790 856
rect 138958 734 139802 856
rect 139970 734 140814 856
rect 140982 734 141826 856
rect 141994 734 142838 856
rect 143006 734 143850 856
rect 144018 734 144862 856
rect 145030 734 145874 856
rect 146042 734 146886 856
rect 147054 734 148470 856
<< metal3 >>
rect 149493 114248 150293 114368
rect 149493 38088 150293 38208
<< obsm3 >>
rect 4210 114448 149493 150381
rect 4210 114168 149413 114448
rect 4210 38288 149493 114168
rect 4210 38008 149413 38288
rect 4210 2143 149493 38008
<< metal4 >>
rect 4208 2128 4528 150192
rect 19568 2128 19888 150192
rect 34928 2128 35248 150192
rect 50288 2128 50608 150192
rect 65648 2128 65968 150192
rect 81008 2128 81328 150192
rect 96368 2128 96688 150192
rect 111728 2128 112048 150192
rect 127088 2128 127408 150192
rect 142448 2128 142768 150192
<< obsm4 >>
rect 12203 150272 141621 150381
rect 12203 2347 19488 150272
rect 19968 2347 34848 150272
rect 35328 2347 50208 150272
rect 50688 2347 65568 150272
rect 66048 2347 80928 150272
rect 81408 2347 96288 150272
rect 96768 2347 111648 150272
rect 112128 2347 127008 150272
rect 127488 2347 141621 150272
<< labels >>
rlabel metal2 s 3238 0 3294 800 6 i_addr[0]
port 1 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 i_addr[1]
port 2 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 i_addr[2]
port 3 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 i_addr[3]
port 4 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 i_addr[4]
port 5 nsew signal input
rlabel metal3 s 149493 38088 150293 38208 6 i_clk
port 6 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 i_data[0]
port 7 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 i_data[100]
port 8 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 i_data[101]
port 9 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 i_data[102]
port 10 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 i_data[103]
port 11 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 i_data[104]
port 12 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 i_data[105]
port 13 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 i_data[106]
port 14 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 i_data[107]
port 15 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 i_data[108]
port 16 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 i_data[109]
port 17 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 i_data[10]
port 18 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 i_data[110]
port 19 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 i_data[111]
port 20 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 i_data[112]
port 21 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 i_data[113]
port 22 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 i_data[114]
port 23 nsew signal input
rlabel metal2 s 124678 0 124734 800 6 i_data[115]
port 24 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 i_data[116]
port 25 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 i_data[117]
port 26 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 i_data[118]
port 27 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 i_data[119]
port 28 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 i_data[11]
port 29 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 i_data[120]
port 30 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 i_data[121]
port 31 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 i_data[122]
port 32 nsew signal input
rlabel metal2 s 132774 0 132830 800 6 i_data[123]
port 33 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 i_data[124]
port 34 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 i_data[125]
port 35 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 i_data[126]
port 36 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 i_data[127]
port 37 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 i_data[128]
port 38 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 i_data[129]
port 39 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 i_data[12]
port 40 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 i_data[130]
port 41 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 i_data[131]
port 42 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 i_data[132]
port 43 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 i_data[133]
port 44 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 i_data[134]
port 45 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 i_data[135]
port 46 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 i_data[136]
port 47 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 i_data[137]
port 48 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 i_data[13]
port 49 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 i_data[14]
port 50 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 i_data[15]
port 51 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 i_data[16]
port 52 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 i_data[17]
port 53 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 i_data[18]
port 54 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 i_data[19]
port 55 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 i_data[1]
port 56 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 i_data[20]
port 57 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 i_data[21]
port 58 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 i_data[22]
port 59 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 i_data[23]
port 60 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 i_data[24]
port 61 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 i_data[25]
port 62 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 i_data[26]
port 63 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 i_data[27]
port 64 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 i_data[28]
port 65 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 i_data[29]
port 66 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 i_data[2]
port 67 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 i_data[30]
port 68 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 i_data[31]
port 69 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 i_data[32]
port 70 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 i_data[33]
port 71 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 i_data[34]
port 72 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 i_data[35]
port 73 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 i_data[36]
port 74 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 i_data[37]
port 75 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 i_data[38]
port 76 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 i_data[39]
port 77 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 i_data[3]
port 78 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 i_data[40]
port 79 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 i_data[41]
port 80 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 i_data[42]
port 81 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 i_data[43]
port 82 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 i_data[44]
port 83 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 i_data[45]
port 84 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 i_data[46]
port 85 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 i_data[47]
port 86 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 i_data[48]
port 87 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 i_data[49]
port 88 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 i_data[4]
port 89 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 i_data[50]
port 90 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 i_data[51]
port 91 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 i_data[52]
port 92 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 i_data[53]
port 93 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 i_data[54]
port 94 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 i_data[55]
port 95 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 i_data[56]
port 96 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 i_data[57]
port 97 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 i_data[58]
port 98 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 i_data[59]
port 99 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 i_data[5]
port 100 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 i_data[60]
port 101 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 i_data[61]
port 102 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 i_data[62]
port 103 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 i_data[63]
port 104 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 i_data[64]
port 105 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 i_data[65]
port 106 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 i_data[66]
port 107 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 i_data[67]
port 108 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 i_data[68]
port 109 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 i_data[69]
port 110 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 i_data[6]
port 111 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 i_data[70]
port 112 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 i_data[71]
port 113 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 i_data[72]
port 114 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 i_data[73]
port 115 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 i_data[74]
port 116 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 i_data[75]
port 117 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 i_data[76]
port 118 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 i_data[77]
port 119 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 i_data[78]
port 120 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 i_data[79]
port 121 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 i_data[7]
port 122 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 i_data[80]
port 123 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 i_data[81]
port 124 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 i_data[82]
port 125 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 i_data[83]
port 126 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 i_data[84]
port 127 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 i_data[85]
port 128 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 i_data[86]
port 129 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 i_data[87]
port 130 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 i_data[88]
port 131 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 i_data[89]
port 132 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 i_data[8]
port 133 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 i_data[90]
port 134 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 i_data[91]
port 135 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 i_data[92]
port 136 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 i_data[93]
port 137 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 i_data[94]
port 138 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 i_data[95]
port 139 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 i_data[96]
port 140 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 i_data[97]
port 141 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 i_data[98]
port 142 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 i_data[99]
port 143 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 i_data[9]
port 144 nsew signal input
rlabel metal3 s 149493 114248 150293 114368 6 i_rst
port 145 nsew signal input
rlabel metal2 s 144918 151637 144974 152437 6 i_we
port 146 nsew signal input
rlabel metal2 s 5262 151637 5318 152437 6 o_data[0]
port 147 nsew signal output
rlabel metal2 s 106462 151637 106518 152437 6 o_data[100]
port 148 nsew signal output
rlabel metal2 s 107474 151637 107530 152437 6 o_data[101]
port 149 nsew signal output
rlabel metal2 s 108486 151637 108542 152437 6 o_data[102]
port 150 nsew signal output
rlabel metal2 s 109498 151637 109554 152437 6 o_data[103]
port 151 nsew signal output
rlabel metal2 s 110510 151637 110566 152437 6 o_data[104]
port 152 nsew signal output
rlabel metal2 s 111522 151637 111578 152437 6 o_data[105]
port 153 nsew signal output
rlabel metal2 s 112534 151637 112590 152437 6 o_data[106]
port 154 nsew signal output
rlabel metal2 s 113546 151637 113602 152437 6 o_data[107]
port 155 nsew signal output
rlabel metal2 s 114558 151637 114614 152437 6 o_data[108]
port 156 nsew signal output
rlabel metal2 s 115570 151637 115626 152437 6 o_data[109]
port 157 nsew signal output
rlabel metal2 s 15382 151637 15438 152437 6 o_data[10]
port 158 nsew signal output
rlabel metal2 s 116582 151637 116638 152437 6 o_data[110]
port 159 nsew signal output
rlabel metal2 s 117594 151637 117650 152437 6 o_data[111]
port 160 nsew signal output
rlabel metal2 s 118606 151637 118662 152437 6 o_data[112]
port 161 nsew signal output
rlabel metal2 s 119618 151637 119674 152437 6 o_data[113]
port 162 nsew signal output
rlabel metal2 s 120630 151637 120686 152437 6 o_data[114]
port 163 nsew signal output
rlabel metal2 s 121642 151637 121698 152437 6 o_data[115]
port 164 nsew signal output
rlabel metal2 s 122654 151637 122710 152437 6 o_data[116]
port 165 nsew signal output
rlabel metal2 s 123666 151637 123722 152437 6 o_data[117]
port 166 nsew signal output
rlabel metal2 s 124678 151637 124734 152437 6 o_data[118]
port 167 nsew signal output
rlabel metal2 s 125690 151637 125746 152437 6 o_data[119]
port 168 nsew signal output
rlabel metal2 s 16394 151637 16450 152437 6 o_data[11]
port 169 nsew signal output
rlabel metal2 s 126702 151637 126758 152437 6 o_data[120]
port 170 nsew signal output
rlabel metal2 s 127714 151637 127770 152437 6 o_data[121]
port 171 nsew signal output
rlabel metal2 s 128726 151637 128782 152437 6 o_data[122]
port 172 nsew signal output
rlabel metal2 s 129738 151637 129794 152437 6 o_data[123]
port 173 nsew signal output
rlabel metal2 s 130750 151637 130806 152437 6 o_data[124]
port 174 nsew signal output
rlabel metal2 s 131762 151637 131818 152437 6 o_data[125]
port 175 nsew signal output
rlabel metal2 s 132774 151637 132830 152437 6 o_data[126]
port 176 nsew signal output
rlabel metal2 s 133786 151637 133842 152437 6 o_data[127]
port 177 nsew signal output
rlabel metal2 s 134798 151637 134854 152437 6 o_data[128]
port 178 nsew signal output
rlabel metal2 s 135810 151637 135866 152437 6 o_data[129]
port 179 nsew signal output
rlabel metal2 s 17406 151637 17462 152437 6 o_data[12]
port 180 nsew signal output
rlabel metal2 s 136822 151637 136878 152437 6 o_data[130]
port 181 nsew signal output
rlabel metal2 s 137834 151637 137890 152437 6 o_data[131]
port 182 nsew signal output
rlabel metal2 s 138846 151637 138902 152437 6 o_data[132]
port 183 nsew signal output
rlabel metal2 s 139858 151637 139914 152437 6 o_data[133]
port 184 nsew signal output
rlabel metal2 s 140870 151637 140926 152437 6 o_data[134]
port 185 nsew signal output
rlabel metal2 s 141882 151637 141938 152437 6 o_data[135]
port 186 nsew signal output
rlabel metal2 s 142894 151637 142950 152437 6 o_data[136]
port 187 nsew signal output
rlabel metal2 s 143906 151637 143962 152437 6 o_data[137]
port 188 nsew signal output
rlabel metal2 s 18418 151637 18474 152437 6 o_data[13]
port 189 nsew signal output
rlabel metal2 s 19430 151637 19486 152437 6 o_data[14]
port 190 nsew signal output
rlabel metal2 s 20442 151637 20498 152437 6 o_data[15]
port 191 nsew signal output
rlabel metal2 s 21454 151637 21510 152437 6 o_data[16]
port 192 nsew signal output
rlabel metal2 s 22466 151637 22522 152437 6 o_data[17]
port 193 nsew signal output
rlabel metal2 s 23478 151637 23534 152437 6 o_data[18]
port 194 nsew signal output
rlabel metal2 s 24490 151637 24546 152437 6 o_data[19]
port 195 nsew signal output
rlabel metal2 s 6274 151637 6330 152437 6 o_data[1]
port 196 nsew signal output
rlabel metal2 s 25502 151637 25558 152437 6 o_data[20]
port 197 nsew signal output
rlabel metal2 s 26514 151637 26570 152437 6 o_data[21]
port 198 nsew signal output
rlabel metal2 s 27526 151637 27582 152437 6 o_data[22]
port 199 nsew signal output
rlabel metal2 s 28538 151637 28594 152437 6 o_data[23]
port 200 nsew signal output
rlabel metal2 s 29550 151637 29606 152437 6 o_data[24]
port 201 nsew signal output
rlabel metal2 s 30562 151637 30618 152437 6 o_data[25]
port 202 nsew signal output
rlabel metal2 s 31574 151637 31630 152437 6 o_data[26]
port 203 nsew signal output
rlabel metal2 s 32586 151637 32642 152437 6 o_data[27]
port 204 nsew signal output
rlabel metal2 s 33598 151637 33654 152437 6 o_data[28]
port 205 nsew signal output
rlabel metal2 s 34610 151637 34666 152437 6 o_data[29]
port 206 nsew signal output
rlabel metal2 s 7286 151637 7342 152437 6 o_data[2]
port 207 nsew signal output
rlabel metal2 s 35622 151637 35678 152437 6 o_data[30]
port 208 nsew signal output
rlabel metal2 s 36634 151637 36690 152437 6 o_data[31]
port 209 nsew signal output
rlabel metal2 s 37646 151637 37702 152437 6 o_data[32]
port 210 nsew signal output
rlabel metal2 s 38658 151637 38714 152437 6 o_data[33]
port 211 nsew signal output
rlabel metal2 s 39670 151637 39726 152437 6 o_data[34]
port 212 nsew signal output
rlabel metal2 s 40682 151637 40738 152437 6 o_data[35]
port 213 nsew signal output
rlabel metal2 s 41694 151637 41750 152437 6 o_data[36]
port 214 nsew signal output
rlabel metal2 s 42706 151637 42762 152437 6 o_data[37]
port 215 nsew signal output
rlabel metal2 s 43718 151637 43774 152437 6 o_data[38]
port 216 nsew signal output
rlabel metal2 s 44730 151637 44786 152437 6 o_data[39]
port 217 nsew signal output
rlabel metal2 s 8298 151637 8354 152437 6 o_data[3]
port 218 nsew signal output
rlabel metal2 s 45742 151637 45798 152437 6 o_data[40]
port 219 nsew signal output
rlabel metal2 s 46754 151637 46810 152437 6 o_data[41]
port 220 nsew signal output
rlabel metal2 s 47766 151637 47822 152437 6 o_data[42]
port 221 nsew signal output
rlabel metal2 s 48778 151637 48834 152437 6 o_data[43]
port 222 nsew signal output
rlabel metal2 s 49790 151637 49846 152437 6 o_data[44]
port 223 nsew signal output
rlabel metal2 s 50802 151637 50858 152437 6 o_data[45]
port 224 nsew signal output
rlabel metal2 s 51814 151637 51870 152437 6 o_data[46]
port 225 nsew signal output
rlabel metal2 s 52826 151637 52882 152437 6 o_data[47]
port 226 nsew signal output
rlabel metal2 s 53838 151637 53894 152437 6 o_data[48]
port 227 nsew signal output
rlabel metal2 s 54850 151637 54906 152437 6 o_data[49]
port 228 nsew signal output
rlabel metal2 s 9310 151637 9366 152437 6 o_data[4]
port 229 nsew signal output
rlabel metal2 s 55862 151637 55918 152437 6 o_data[50]
port 230 nsew signal output
rlabel metal2 s 56874 151637 56930 152437 6 o_data[51]
port 231 nsew signal output
rlabel metal2 s 57886 151637 57942 152437 6 o_data[52]
port 232 nsew signal output
rlabel metal2 s 58898 151637 58954 152437 6 o_data[53]
port 233 nsew signal output
rlabel metal2 s 59910 151637 59966 152437 6 o_data[54]
port 234 nsew signal output
rlabel metal2 s 60922 151637 60978 152437 6 o_data[55]
port 235 nsew signal output
rlabel metal2 s 61934 151637 61990 152437 6 o_data[56]
port 236 nsew signal output
rlabel metal2 s 62946 151637 63002 152437 6 o_data[57]
port 237 nsew signal output
rlabel metal2 s 63958 151637 64014 152437 6 o_data[58]
port 238 nsew signal output
rlabel metal2 s 64970 151637 65026 152437 6 o_data[59]
port 239 nsew signal output
rlabel metal2 s 10322 151637 10378 152437 6 o_data[5]
port 240 nsew signal output
rlabel metal2 s 65982 151637 66038 152437 6 o_data[60]
port 241 nsew signal output
rlabel metal2 s 66994 151637 67050 152437 6 o_data[61]
port 242 nsew signal output
rlabel metal2 s 68006 151637 68062 152437 6 o_data[62]
port 243 nsew signal output
rlabel metal2 s 69018 151637 69074 152437 6 o_data[63]
port 244 nsew signal output
rlabel metal2 s 70030 151637 70086 152437 6 o_data[64]
port 245 nsew signal output
rlabel metal2 s 71042 151637 71098 152437 6 o_data[65]
port 246 nsew signal output
rlabel metal2 s 72054 151637 72110 152437 6 o_data[66]
port 247 nsew signal output
rlabel metal2 s 73066 151637 73122 152437 6 o_data[67]
port 248 nsew signal output
rlabel metal2 s 74078 151637 74134 152437 6 o_data[68]
port 249 nsew signal output
rlabel metal2 s 75090 151637 75146 152437 6 o_data[69]
port 250 nsew signal output
rlabel metal2 s 11334 151637 11390 152437 6 o_data[6]
port 251 nsew signal output
rlabel metal2 s 76102 151637 76158 152437 6 o_data[70]
port 252 nsew signal output
rlabel metal2 s 77114 151637 77170 152437 6 o_data[71]
port 253 nsew signal output
rlabel metal2 s 78126 151637 78182 152437 6 o_data[72]
port 254 nsew signal output
rlabel metal2 s 79138 151637 79194 152437 6 o_data[73]
port 255 nsew signal output
rlabel metal2 s 80150 151637 80206 152437 6 o_data[74]
port 256 nsew signal output
rlabel metal2 s 81162 151637 81218 152437 6 o_data[75]
port 257 nsew signal output
rlabel metal2 s 82174 151637 82230 152437 6 o_data[76]
port 258 nsew signal output
rlabel metal2 s 83186 151637 83242 152437 6 o_data[77]
port 259 nsew signal output
rlabel metal2 s 84198 151637 84254 152437 6 o_data[78]
port 260 nsew signal output
rlabel metal2 s 85210 151637 85266 152437 6 o_data[79]
port 261 nsew signal output
rlabel metal2 s 12346 151637 12402 152437 6 o_data[7]
port 262 nsew signal output
rlabel metal2 s 86222 151637 86278 152437 6 o_data[80]
port 263 nsew signal output
rlabel metal2 s 87234 151637 87290 152437 6 o_data[81]
port 264 nsew signal output
rlabel metal2 s 88246 151637 88302 152437 6 o_data[82]
port 265 nsew signal output
rlabel metal2 s 89258 151637 89314 152437 6 o_data[83]
port 266 nsew signal output
rlabel metal2 s 90270 151637 90326 152437 6 o_data[84]
port 267 nsew signal output
rlabel metal2 s 91282 151637 91338 152437 6 o_data[85]
port 268 nsew signal output
rlabel metal2 s 92294 151637 92350 152437 6 o_data[86]
port 269 nsew signal output
rlabel metal2 s 93306 151637 93362 152437 6 o_data[87]
port 270 nsew signal output
rlabel metal2 s 94318 151637 94374 152437 6 o_data[88]
port 271 nsew signal output
rlabel metal2 s 95330 151637 95386 152437 6 o_data[89]
port 272 nsew signal output
rlabel metal2 s 13358 151637 13414 152437 6 o_data[8]
port 273 nsew signal output
rlabel metal2 s 96342 151637 96398 152437 6 o_data[90]
port 274 nsew signal output
rlabel metal2 s 97354 151637 97410 152437 6 o_data[91]
port 275 nsew signal output
rlabel metal2 s 98366 151637 98422 152437 6 o_data[92]
port 276 nsew signal output
rlabel metal2 s 99378 151637 99434 152437 6 o_data[93]
port 277 nsew signal output
rlabel metal2 s 100390 151637 100446 152437 6 o_data[94]
port 278 nsew signal output
rlabel metal2 s 101402 151637 101458 152437 6 o_data[95]
port 279 nsew signal output
rlabel metal2 s 102414 151637 102470 152437 6 o_data[96]
port 280 nsew signal output
rlabel metal2 s 103426 151637 103482 152437 6 o_data[97]
port 281 nsew signal output
rlabel metal2 s 104438 151637 104494 152437 6 o_data[98]
port 282 nsew signal output
rlabel metal2 s 105450 151637 105506 152437 6 o_data[99]
port 283 nsew signal output
rlabel metal2 s 14370 151637 14426 152437 6 o_data[9]
port 284 nsew signal output
rlabel metal4 s 4208 2128 4528 150192 6 vccd1
port 285 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 150192 6 vccd1
port 285 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 150192 6 vccd1
port 285 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 150192 6 vccd1
port 285 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 150192 6 vccd1
port 285 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 150192 6 vssd1
port 286 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 150192 6 vssd1
port 286 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 150192 6 vssd1
port 286 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 150192 6 vssd1
port 286 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 150192 6 vssd1
port 286 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 150293 152437
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 57125620
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/icache_ram/runs/22_09_09_18_43/results/signoff/icache_ram.magic.gds
string GDS_START 288304
<< end >>

