magic
tech gf180mcuD
magscale 1 10
timestamp 1699806575
<< nwell >>
rect 1258 66233 158678 66726
rect 1258 66208 30248 66233
rect 1258 65479 14749 65504
rect 1258 64665 158678 65479
rect 1258 64640 14637 64665
rect 1258 63911 19005 63936
rect 1258 63097 158678 63911
rect 1258 63072 10381 63097
rect 1258 62343 14301 62368
rect 1258 61529 158678 62343
rect 1258 61504 24829 61529
rect 1258 60775 10381 60800
rect 1258 59961 158678 60775
rect 1258 59936 9821 59961
rect 1258 59207 13629 59232
rect 1258 58393 158678 59207
rect 1258 58368 25432 58393
rect 1258 57639 10381 57664
rect 1258 56825 158678 57639
rect 1258 56800 9597 56825
rect 1258 56071 29981 56096
rect 1258 55257 158678 56071
rect 1258 55232 10493 55257
rect 1258 54503 18669 54528
rect 1258 53689 158678 54503
rect 1258 53664 7021 53689
rect 1258 52935 6909 52960
rect 1258 52121 158678 52935
rect 1258 52096 7805 52121
rect 1258 51367 13181 51392
rect 1258 50553 158678 51367
rect 1258 50528 6461 50553
rect 1258 49799 18669 49824
rect 1258 48985 158678 49799
rect 1258 48960 8365 48985
rect 1258 48231 6349 48256
rect 1258 47417 158678 48231
rect 1258 47392 9261 47417
rect 1258 46663 19677 46688
rect 1258 45849 158678 46663
rect 1258 45824 2989 45849
rect 1258 45095 10381 45120
rect 1258 44281 158678 45095
rect 1258 44256 9485 44281
rect 1258 43527 3549 43552
rect 1258 42713 158678 43527
rect 1258 42688 2989 42713
rect 1258 41959 22029 41984
rect 1258 41145 158678 41959
rect 1258 41120 14301 41145
rect 1258 40391 3213 40416
rect 1258 39577 158678 40391
rect 1258 39552 2989 39577
rect 1258 38823 14120 38848
rect 1258 38009 158678 38823
rect 1258 37984 2989 38009
rect 1258 37255 19565 37280
rect 1258 36441 158678 37255
rect 1258 36416 8701 36441
rect 1258 35687 4669 35712
rect 1258 34873 158678 35687
rect 1258 34848 2989 34873
rect 1258 34119 4445 34144
rect 1258 33305 158678 34119
rect 1258 33280 6461 33305
rect 1258 32551 20573 32576
rect 1258 31737 158678 32551
rect 1258 31712 32669 31737
rect 1258 30983 4109 31008
rect 1258 30169 158678 30983
rect 1258 30144 7581 30169
rect 1258 29415 5901 29440
rect 1258 28601 158678 29415
rect 1258 28576 8141 28601
rect 1258 27847 12733 27872
rect 1258 27033 158678 27847
rect 1258 27008 26509 27033
rect 1258 26279 13965 26304
rect 1258 25465 158678 26279
rect 1258 25440 8589 25465
rect 1258 24711 11277 24736
rect 1258 23897 158678 24711
rect 1258 23872 6797 23897
rect 1258 23143 19341 23168
rect 1258 22329 158678 23143
rect 1258 22304 10381 22329
rect 1258 21575 6909 21600
rect 1258 20761 158678 21575
rect 1258 20736 18333 20761
rect 1258 20007 6909 20032
rect 1258 19193 158678 20007
rect 1258 19168 14301 19193
rect 1258 18439 27853 18464
rect 1258 17625 158678 18439
rect 1258 17600 8813 17625
rect 1258 16871 7736 16896
rect 1258 16057 158678 16871
rect 1258 16032 14301 16057
rect 1258 15303 18669 15328
rect 1258 14489 158678 15303
rect 1258 14464 25725 14489
rect 1258 13735 21736 13760
rect 1258 12921 158678 13735
rect 1258 12896 9821 12921
rect 1258 12167 10381 12192
rect 1258 11353 158678 12167
rect 1258 11328 34349 11353
rect 1258 10599 20685 10624
rect 1258 9785 158678 10599
rect 1258 9760 10829 9785
rect 1258 9031 11277 9056
rect 1258 8217 158678 9031
rect 1258 8192 15981 8217
rect 1258 7463 36365 7488
rect 1258 6649 158678 7463
rect 1258 6624 14301 6649
rect 1258 5895 19789 5920
rect 1258 5081 158678 5895
rect 1258 5056 17213 5081
rect 1258 4327 14189 4352
rect 1258 3513 158678 4327
rect 1258 3488 33005 3513
<< pwell >>
rect 1258 65504 158678 66208
rect 1258 63936 158678 64640
rect 1258 62368 158678 63072
rect 1258 60800 158678 61504
rect 1258 59232 158678 59936
rect 1258 57664 158678 58368
rect 1258 56096 158678 56800
rect 1258 54528 158678 55232
rect 1258 52960 158678 53664
rect 1258 51392 158678 52096
rect 1258 49824 158678 50528
rect 1258 48256 158678 48960
rect 1258 46688 158678 47392
rect 1258 45120 158678 45824
rect 1258 43552 158678 44256
rect 1258 41984 158678 42688
rect 1258 40416 158678 41120
rect 1258 38848 158678 39552
rect 1258 37280 158678 37984
rect 1258 35712 158678 36416
rect 1258 34144 158678 34848
rect 1258 32576 158678 33280
rect 1258 31008 158678 31712
rect 1258 29440 158678 30144
rect 1258 27872 158678 28576
rect 1258 26304 158678 27008
rect 1258 24736 158678 25440
rect 1258 23168 158678 23872
rect 1258 21600 158678 22304
rect 1258 20032 158678 20736
rect 1258 18464 158678 19168
rect 1258 16896 158678 17600
rect 1258 15328 158678 16032
rect 1258 13760 158678 14464
rect 1258 12192 158678 12896
rect 1258 10624 158678 11328
rect 1258 9056 158678 9760
rect 1258 7488 158678 8192
rect 1258 5920 158678 6624
rect 1258 4352 158678 5056
rect 1258 3050 158678 3488
<< obsm1 >>
rect 1344 3076 158592 66834
<< obsm2 >>
rect 1932 578 158564 67966
<< metal3 >>
rect 159200 65408 160000 65520
rect 159200 63840 160000 63952
rect 159200 62272 160000 62384
rect 159200 60704 160000 60816
rect 159200 59136 160000 59248
rect 159200 57568 160000 57680
rect 159200 56000 160000 56112
rect 159200 54432 160000 54544
rect 159200 52864 160000 52976
rect 159200 51296 160000 51408
rect 159200 49728 160000 49840
rect 159200 48160 160000 48272
rect 159200 46592 160000 46704
rect 159200 45024 160000 45136
rect 159200 43456 160000 43568
rect 159200 41888 160000 42000
rect 159200 40320 160000 40432
rect 159200 38752 160000 38864
rect 159200 37184 160000 37296
rect 159200 35616 160000 35728
rect 159200 34048 160000 34160
rect 159200 32480 160000 32592
rect 159200 30912 160000 31024
rect 159200 29344 160000 29456
rect 159200 27776 160000 27888
rect 159200 26208 160000 26320
rect 159200 24640 160000 24752
rect 159200 23072 160000 23184
rect 159200 21504 160000 21616
rect 159200 19936 160000 20048
rect 159200 18368 160000 18480
rect 159200 16800 160000 16912
rect 159200 15232 160000 15344
rect 159200 13664 160000 13776
rect 159200 12096 160000 12208
rect 159200 10528 160000 10640
rect 159200 8960 160000 9072
rect 159200 7392 160000 7504
rect 159200 5824 160000 5936
rect 159200 4256 160000 4368
<< obsm3 >>
rect 1922 65580 159200 67956
rect 1922 65348 159140 65580
rect 1922 64012 159200 65348
rect 1922 63780 159140 64012
rect 1922 62444 159200 63780
rect 1922 62212 159140 62444
rect 1922 60876 159200 62212
rect 1922 60644 159140 60876
rect 1922 59308 159200 60644
rect 1922 59076 159140 59308
rect 1922 57740 159200 59076
rect 1922 57508 159140 57740
rect 1922 56172 159200 57508
rect 1922 55940 159140 56172
rect 1922 54604 159200 55940
rect 1922 54372 159140 54604
rect 1922 53036 159200 54372
rect 1922 52804 159140 53036
rect 1922 51468 159200 52804
rect 1922 51236 159140 51468
rect 1922 49900 159200 51236
rect 1922 49668 159140 49900
rect 1922 48332 159200 49668
rect 1922 48100 159140 48332
rect 1922 46764 159200 48100
rect 1922 46532 159140 46764
rect 1922 45196 159200 46532
rect 1922 44964 159140 45196
rect 1922 43628 159200 44964
rect 1922 43396 159140 43628
rect 1922 42060 159200 43396
rect 1922 41828 159140 42060
rect 1922 40492 159200 41828
rect 1922 40260 159140 40492
rect 1922 38924 159200 40260
rect 1922 38692 159140 38924
rect 1922 37356 159200 38692
rect 1922 37124 159140 37356
rect 1922 35788 159200 37124
rect 1922 35556 159140 35788
rect 1922 34220 159200 35556
rect 1922 33988 159140 34220
rect 1922 32652 159200 33988
rect 1922 32420 159140 32652
rect 1922 31084 159200 32420
rect 1922 30852 159140 31084
rect 1922 29516 159200 30852
rect 1922 29284 159140 29516
rect 1922 27948 159200 29284
rect 1922 27716 159140 27948
rect 1922 26380 159200 27716
rect 1922 26148 159140 26380
rect 1922 24812 159200 26148
rect 1922 24580 159140 24812
rect 1922 23244 159200 24580
rect 1922 23012 159140 23244
rect 1922 21676 159200 23012
rect 1922 21444 159140 21676
rect 1922 20108 159200 21444
rect 1922 19876 159140 20108
rect 1922 18540 159200 19876
rect 1922 18308 159140 18540
rect 1922 16972 159200 18308
rect 1922 16740 159140 16972
rect 1922 15404 159200 16740
rect 1922 15172 159140 15404
rect 1922 13836 159200 15172
rect 1922 13604 159140 13836
rect 1922 12268 159200 13604
rect 1922 12036 159140 12268
rect 1922 10700 159200 12036
rect 1922 10468 159140 10700
rect 1922 9132 159200 10468
rect 1922 8900 159140 9132
rect 1922 7564 159200 8900
rect 1922 7332 159140 7564
rect 1922 5996 159200 7332
rect 1922 5764 159140 5996
rect 1922 4428 159200 5764
rect 1922 4196 159140 4428
rect 1922 588 159200 4196
<< metal4 >>
rect 4448 3076 4768 66700
rect 19808 3076 20128 66700
rect 35168 3076 35488 66700
rect 50528 3076 50848 66700
rect 65888 3076 66208 66700
rect 81248 3076 81568 66700
rect 96608 3076 96928 66700
rect 111968 3076 112288 66700
rect 127328 3076 127648 66700
rect 142688 3076 143008 66700
rect 158048 3076 158368 66700
<< obsm4 >>
rect 9660 66760 155764 67518
rect 9660 3016 19748 66760
rect 20188 3016 35108 66760
rect 35548 3016 50468 66760
rect 50908 3016 65828 66760
rect 66268 3016 81188 66760
rect 81628 3016 96548 66760
rect 96988 3016 111908 66760
rect 112348 3016 127268 66760
rect 127708 3016 142628 66760
rect 143068 3016 155764 66760
rect 9660 690 155764 3016
<< labels >>
rlabel metal3 s 159200 7392 160000 7504 6 i_addr[0]
port 1 nsew signal input
rlabel metal3 s 159200 12096 160000 12208 6 i_addr[1]
port 2 nsew signal input
rlabel metal3 s 159200 16800 160000 16912 6 i_addr[2]
port 3 nsew signal input
rlabel metal3 s 159200 21504 160000 21616 6 i_addr[3]
port 4 nsew signal input
rlabel metal3 s 159200 26208 160000 26320 6 i_addr[4]
port 5 nsew signal input
rlabel metal3 s 159200 30912 160000 31024 6 i_addr[5]
port 6 nsew signal input
rlabel metal3 s 159200 4256 160000 4368 6 i_clk
port 7 nsew signal input
rlabel metal3 s 159200 8960 160000 9072 6 i_data[0]
port 8 nsew signal input
rlabel metal3 s 159200 48160 160000 48272 6 i_data[10]
port 9 nsew signal input
rlabel metal3 s 159200 51296 160000 51408 6 i_data[11]
port 10 nsew signal input
rlabel metal3 s 159200 54432 160000 54544 6 i_data[12]
port 11 nsew signal input
rlabel metal3 s 159200 57568 160000 57680 6 i_data[13]
port 12 nsew signal input
rlabel metal3 s 159200 60704 160000 60816 6 i_data[14]
port 13 nsew signal input
rlabel metal3 s 159200 63840 160000 63952 6 i_data[15]
port 14 nsew signal input
rlabel metal3 s 159200 13664 160000 13776 6 i_data[1]
port 15 nsew signal input
rlabel metal3 s 159200 18368 160000 18480 6 i_data[2]
port 16 nsew signal input
rlabel metal3 s 159200 23072 160000 23184 6 i_data[3]
port 17 nsew signal input
rlabel metal3 s 159200 27776 160000 27888 6 i_data[4]
port 18 nsew signal input
rlabel metal3 s 159200 32480 160000 32592 6 i_data[5]
port 19 nsew signal input
rlabel metal3 s 159200 35616 160000 35728 6 i_data[6]
port 20 nsew signal input
rlabel metal3 s 159200 38752 160000 38864 6 i_data[7]
port 21 nsew signal input
rlabel metal3 s 159200 41888 160000 42000 6 i_data[8]
port 22 nsew signal input
rlabel metal3 s 159200 45024 160000 45136 6 i_data[9]
port 23 nsew signal input
rlabel metal3 s 159200 5824 160000 5936 6 i_we
port 24 nsew signal input
rlabel metal3 s 159200 10528 160000 10640 6 o_data[0]
port 25 nsew signal output
rlabel metal3 s 159200 49728 160000 49840 6 o_data[10]
port 26 nsew signal output
rlabel metal3 s 159200 52864 160000 52976 6 o_data[11]
port 27 nsew signal output
rlabel metal3 s 159200 56000 160000 56112 6 o_data[12]
port 28 nsew signal output
rlabel metal3 s 159200 59136 160000 59248 6 o_data[13]
port 29 nsew signal output
rlabel metal3 s 159200 62272 160000 62384 6 o_data[14]
port 30 nsew signal output
rlabel metal3 s 159200 65408 160000 65520 6 o_data[15]
port 31 nsew signal output
rlabel metal3 s 159200 15232 160000 15344 6 o_data[1]
port 32 nsew signal output
rlabel metal3 s 159200 19936 160000 20048 6 o_data[2]
port 33 nsew signal output
rlabel metal3 s 159200 24640 160000 24752 6 o_data[3]
port 34 nsew signal output
rlabel metal3 s 159200 29344 160000 29456 6 o_data[4]
port 35 nsew signal output
rlabel metal3 s 159200 34048 160000 34160 6 o_data[5]
port 36 nsew signal output
rlabel metal3 s 159200 37184 160000 37296 6 o_data[6]
port 37 nsew signal output
rlabel metal3 s 159200 40320 160000 40432 6 o_data[7]
port 38 nsew signal output
rlabel metal3 s 159200 43456 160000 43568 6 o_data[8]
port 39 nsew signal output
rlabel metal3 s 159200 46592 160000 46704 6 o_data[9]
port 40 nsew signal output
rlabel metal4 s 4448 3076 4768 66700 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 66700 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 66700 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 66700 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 66700 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 66700 6 vccd1
port 41 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 66700 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 66700 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 66700 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 66700 6 vssd1
port 42 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 66700 6 vssd1
port 42 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 160000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9276466
string GDS_FILE /home/piotro/caravel_user_project/openlane/int_ram/runs/23_11_12_17_26/results/signoff/int_ram.magic.gds
string GDS_START 223822
<< end >>

